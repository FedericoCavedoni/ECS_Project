library IEEE;
  use IEEE.std_logic_1164.all;
  use IEEE.numeric_std.all;

entity ddfs_lut_65536_16bit is
  port (
    address  : in  std_logic_vector(15 downto 0);
    ddfs_out : out std_logic_vector(15 downto 0)
  );
end entity;

architecture rtl of ddfs_lut_65536_16bit is

  type LUT_t is array (natural range 0 to 65535) of integer;
  constant LUT: LUT_t := (
    0 => 0,
    1 => 3,
    2 => 6,
    3 => 9,
    4 => 13,
    5 => 16,
    6 => 19,
    7 => 22,
    8 => 25,
    9 => 28,
    10 => 31,
    11 => 35,
    12 => 38,
    13 => 41,
    14 => 44,
    15 => 47,
    16 => 50,
    17 => 53,
    18 => 57,
    19 => 60,
    20 => 63,
    21 => 66,
    22 => 69,
    23 => 72,
    24 => 75,
    25 => 79,
    26 => 82,
    27 => 85,
    28 => 88,
    29 => 91,
    30 => 94,
    31 => 97,
    32 => 101,
    33 => 104,
    34 => 107,
    35 => 110,
    36 => 113,
    37 => 116,
    38 => 119,
    39 => 123,
    40 => 126,
    41 => 129,
    42 => 132,
    43 => 135,
    44 => 138,
    45 => 141,
    46 => 145,
    47 => 148,
    48 => 151,
    49 => 154,
    50 => 157,
    51 => 160,
    52 => 163,
    53 => 166,
    54 => 170,
    55 => 173,
    56 => 176,
    57 => 179,
    58 => 182,
    59 => 185,
    60 => 188,
    61 => 192,
    62 => 195,
    63 => 198,
    64 => 201,
    65 => 204,
    66 => 207,
    67 => 210,
    68 => 214,
    69 => 217,
    70 => 220,
    71 => 223,
    72 => 226,
    73 => 229,
    74 => 232,
    75 => 236,
    76 => 239,
    77 => 242,
    78 => 245,
    79 => 248,
    80 => 251,
    81 => 254,
    82 => 258,
    83 => 261,
    84 => 264,
    85 => 267,
    86 => 270,
    87 => 273,
    88 => 276,
    89 => 280,
    90 => 283,
    91 => 286,
    92 => 289,
    93 => 292,
    94 => 295,
    95 => 298,
    96 => 302,
    97 => 305,
    98 => 308,
    99 => 311,
    100 => 314,
    101 => 317,
    102 => 320,
    103 => 324,
    104 => 327,
    105 => 330,
    106 => 333,
    107 => 336,
    108 => 339,
    109 => 342,
    110 => 346,
    111 => 349,
    112 => 352,
    113 => 355,
    114 => 358,
    115 => 361,
    116 => 364,
    117 => 368,
    118 => 371,
    119 => 374,
    120 => 377,
    121 => 380,
    122 => 383,
    123 => 386,
    124 => 390,
    125 => 393,
    126 => 396,
    127 => 399,
    128 => 402,
    129 => 405,
    130 => 408,
    131 => 412,
    132 => 415,
    133 => 418,
    134 => 421,
    135 => 424,
    136 => 427,
    137 => 430,
    138 => 434,
    139 => 437,
    140 => 440,
    141 => 443,
    142 => 446,
    143 => 449,
    144 => 452,
    145 => 456,
    146 => 459,
    147 => 462,
    148 => 465,
    149 => 468,
    150 => 471,
    151 => 474,
    152 => 477,
    153 => 481,
    154 => 484,
    155 => 487,
    156 => 490,
    157 => 493,
    158 => 496,
    159 => 499,
    160 => 503,
    161 => 506,
    162 => 509,
    163 => 512,
    164 => 515,
    165 => 518,
    166 => 521,
    167 => 525,
    168 => 528,
    169 => 531,
    170 => 534,
    171 => 537,
    172 => 540,
    173 => 543,
    174 => 547,
    175 => 550,
    176 => 553,
    177 => 556,
    178 => 559,
    179 => 562,
    180 => 565,
    181 => 569,
    182 => 572,
    183 => 575,
    184 => 578,
    185 => 581,
    186 => 584,
    187 => 587,
    188 => 591,
    189 => 594,
    190 => 597,
    191 => 600,
    192 => 603,
    193 => 606,
    194 => 609,
    195 => 613,
    196 => 616,
    197 => 619,
    198 => 622,
    199 => 625,
    200 => 628,
    201 => 631,
    202 => 635,
    203 => 638,
    204 => 641,
    205 => 644,
    206 => 647,
    207 => 650,
    208 => 653,
    209 => 657,
    210 => 660,
    211 => 663,
    212 => 666,
    213 => 669,
    214 => 672,
    215 => 675,
    216 => 679,
    217 => 682,
    218 => 685,
    219 => 688,
    220 => 691,
    221 => 694,
    222 => 697,
    223 => 701,
    224 => 704,
    225 => 707,
    226 => 710,
    227 => 713,
    228 => 716,
    229 => 719,
    230 => 722,
    231 => 726,
    232 => 729,
    233 => 732,
    234 => 735,
    235 => 738,
    236 => 741,
    237 => 744,
    238 => 748,
    239 => 751,
    240 => 754,
    241 => 757,
    242 => 760,
    243 => 763,
    244 => 766,
    245 => 770,
    246 => 773,
    247 => 776,
    248 => 779,
    249 => 782,
    250 => 785,
    251 => 788,
    252 => 792,
    253 => 795,
    254 => 798,
    255 => 801,
    256 => 804,
    257 => 807,
    258 => 810,
    259 => 814,
    260 => 817,
    261 => 820,
    262 => 823,
    263 => 826,
    264 => 829,
    265 => 832,
    266 => 836,
    267 => 839,
    268 => 842,
    269 => 845,
    270 => 848,
    271 => 851,
    272 => 854,
    273 => 858,
    274 => 861,
    275 => 864,
    276 => 867,
    277 => 870,
    278 => 873,
    279 => 876,
    280 => 880,
    281 => 883,
    282 => 886,
    283 => 889,
    284 => 892,
    285 => 895,
    286 => 898,
    287 => 901,
    288 => 905,
    289 => 908,
    290 => 911,
    291 => 914,
    292 => 917,
    293 => 920,
    294 => 923,
    295 => 927,
    296 => 930,
    297 => 933,
    298 => 936,
    299 => 939,
    300 => 942,
    301 => 945,
    302 => 949,
    303 => 952,
    304 => 955,
    305 => 958,
    306 => 961,
    307 => 964,
    308 => 967,
    309 => 971,
    310 => 974,
    311 => 977,
    312 => 980,
    313 => 983,
    314 => 986,
    315 => 989,
    316 => 993,
    317 => 996,
    318 => 999,
    319 => 1002,
    320 => 1005,
    321 => 1008,
    322 => 1011,
    323 => 1015,
    324 => 1018,
    325 => 1021,
    326 => 1024,
    327 => 1027,
    328 => 1030,
    329 => 1033,
    330 => 1037,
    331 => 1040,
    332 => 1043,
    333 => 1046,
    334 => 1049,
    335 => 1052,
    336 => 1055,
    337 => 1059,
    338 => 1062,
    339 => 1065,
    340 => 1068,
    341 => 1071,
    342 => 1074,
    343 => 1077,
    344 => 1080,
    345 => 1084,
    346 => 1087,
    347 => 1090,
    348 => 1093,
    349 => 1096,
    350 => 1099,
    351 => 1102,
    352 => 1106,
    353 => 1109,
    354 => 1112,
    355 => 1115,
    356 => 1118,
    357 => 1121,
    358 => 1124,
    359 => 1128,
    360 => 1131,
    361 => 1134,
    362 => 1137,
    363 => 1140,
    364 => 1143,
    365 => 1146,
    366 => 1150,
    367 => 1153,
    368 => 1156,
    369 => 1159,
    370 => 1162,
    371 => 1165,
    372 => 1168,
    373 => 1172,
    374 => 1175,
    375 => 1178,
    376 => 1181,
    377 => 1184,
    378 => 1187,
    379 => 1190,
    380 => 1194,
    381 => 1197,
    382 => 1200,
    383 => 1203,
    384 => 1206,
    385 => 1209,
    386 => 1212,
    387 => 1215,
    388 => 1219,
    389 => 1222,
    390 => 1225,
    391 => 1228,
    392 => 1231,
    393 => 1234,
    394 => 1237,
    395 => 1241,
    396 => 1244,
    397 => 1247,
    398 => 1250,
    399 => 1253,
    400 => 1256,
    401 => 1259,
    402 => 1263,
    403 => 1266,
    404 => 1269,
    405 => 1272,
    406 => 1275,
    407 => 1278,
    408 => 1281,
    409 => 1285,
    410 => 1288,
    411 => 1291,
    412 => 1294,
    413 => 1297,
    414 => 1300,
    415 => 1303,
    416 => 1307,
    417 => 1310,
    418 => 1313,
    419 => 1316,
    420 => 1319,
    421 => 1322,
    422 => 1325,
    423 => 1328,
    424 => 1332,
    425 => 1335,
    426 => 1338,
    427 => 1341,
    428 => 1344,
    429 => 1347,
    430 => 1350,
    431 => 1354,
    432 => 1357,
    433 => 1360,
    434 => 1363,
    435 => 1366,
    436 => 1369,
    437 => 1372,
    438 => 1376,
    439 => 1379,
    440 => 1382,
    441 => 1385,
    442 => 1388,
    443 => 1391,
    444 => 1394,
    445 => 1398,
    446 => 1401,
    447 => 1404,
    448 => 1407,
    449 => 1410,
    450 => 1413,
    451 => 1416,
    452 => 1420,
    453 => 1423,
    454 => 1426,
    455 => 1429,
    456 => 1432,
    457 => 1435,
    458 => 1438,
    459 => 1441,
    460 => 1445,
    461 => 1448,
    462 => 1451,
    463 => 1454,
    464 => 1457,
    465 => 1460,
    466 => 1463,
    467 => 1467,
    468 => 1470,
    469 => 1473,
    470 => 1476,
    471 => 1479,
    472 => 1482,
    473 => 1485,
    474 => 1489,
    475 => 1492,
    476 => 1495,
    477 => 1498,
    478 => 1501,
    479 => 1504,
    480 => 1507,
    481 => 1511,
    482 => 1514,
    483 => 1517,
    484 => 1520,
    485 => 1523,
    486 => 1526,
    487 => 1529,
    488 => 1532,
    489 => 1536,
    490 => 1539,
    491 => 1542,
    492 => 1545,
    493 => 1548,
    494 => 1551,
    495 => 1554,
    496 => 1558,
    497 => 1561,
    498 => 1564,
    499 => 1567,
    500 => 1570,
    501 => 1573,
    502 => 1576,
    503 => 1580,
    504 => 1583,
    505 => 1586,
    506 => 1589,
    507 => 1592,
    508 => 1595,
    509 => 1598,
    510 => 1602,
    511 => 1605,
    512 => 1608,
    513 => 1611,
    514 => 1614,
    515 => 1617,
    516 => 1620,
    517 => 1623,
    518 => 1627,
    519 => 1630,
    520 => 1633,
    521 => 1636,
    522 => 1639,
    523 => 1642,
    524 => 1645,
    525 => 1649,
    526 => 1652,
    527 => 1655,
    528 => 1658,
    529 => 1661,
    530 => 1664,
    531 => 1667,
    532 => 1671,
    533 => 1674,
    534 => 1677,
    535 => 1680,
    536 => 1683,
    537 => 1686,
    538 => 1689,
    539 => 1693,
    540 => 1696,
    541 => 1699,
    542 => 1702,
    543 => 1705,
    544 => 1708,
    545 => 1711,
    546 => 1714,
    547 => 1718,
    548 => 1721,
    549 => 1724,
    550 => 1727,
    551 => 1730,
    552 => 1733,
    553 => 1736,
    554 => 1740,
    555 => 1743,
    556 => 1746,
    557 => 1749,
    558 => 1752,
    559 => 1755,
    560 => 1758,
    561 => 1762,
    562 => 1765,
    563 => 1768,
    564 => 1771,
    565 => 1774,
    566 => 1777,
    567 => 1780,
    568 => 1783,
    569 => 1787,
    570 => 1790,
    571 => 1793,
    572 => 1796,
    573 => 1799,
    574 => 1802,
    575 => 1805,
    576 => 1809,
    577 => 1812,
    578 => 1815,
    579 => 1818,
    580 => 1821,
    581 => 1824,
    582 => 1827,
    583 => 1831,
    584 => 1834,
    585 => 1837,
    586 => 1840,
    587 => 1843,
    588 => 1846,
    589 => 1849,
    590 => 1852,
    591 => 1856,
    592 => 1859,
    593 => 1862,
    594 => 1865,
    595 => 1868,
    596 => 1871,
    597 => 1874,
    598 => 1878,
    599 => 1881,
    600 => 1884,
    601 => 1887,
    602 => 1890,
    603 => 1893,
    604 => 1896,
    605 => 1900,
    606 => 1903,
    607 => 1906,
    608 => 1909,
    609 => 1912,
    610 => 1915,
    611 => 1918,
    612 => 1921,
    613 => 1925,
    614 => 1928,
    615 => 1931,
    616 => 1934,
    617 => 1937,
    618 => 1940,
    619 => 1943,
    620 => 1947,
    621 => 1950,
    622 => 1953,
    623 => 1956,
    624 => 1959,
    625 => 1962,
    626 => 1965,
    627 => 1969,
    628 => 1972,
    629 => 1975,
    630 => 1978,
    631 => 1981,
    632 => 1984,
    633 => 1987,
    634 => 1990,
    635 => 1994,
    636 => 1997,
    637 => 2000,
    638 => 2003,
    639 => 2006,
    640 => 2009,
    641 => 2012,
    642 => 2016,
    643 => 2019,
    644 => 2022,
    645 => 2025,
    646 => 2028,
    647 => 2031,
    648 => 2034,
    649 => 2038,
    650 => 2041,
    651 => 2044,
    652 => 2047,
    653 => 2050,
    654 => 2053,
    655 => 2056,
    656 => 2059,
    657 => 2063,
    658 => 2066,
    659 => 2069,
    660 => 2072,
    661 => 2075,
    662 => 2078,
    663 => 2081,
    664 => 2085,
    665 => 2088,
    666 => 2091,
    667 => 2094,
    668 => 2097,
    669 => 2100,
    670 => 2103,
    671 => 2106,
    672 => 2110,
    673 => 2113,
    674 => 2116,
    675 => 2119,
    676 => 2122,
    677 => 2125,
    678 => 2128,
    679 => 2132,
    680 => 2135,
    681 => 2138,
    682 => 2141,
    683 => 2144,
    684 => 2147,
    685 => 2150,
    686 => 2154,
    687 => 2157,
    688 => 2160,
    689 => 2163,
    690 => 2166,
    691 => 2169,
    692 => 2172,
    693 => 2175,
    694 => 2179,
    695 => 2182,
    696 => 2185,
    697 => 2188,
    698 => 2191,
    699 => 2194,
    700 => 2197,
    701 => 2201,
    702 => 2204,
    703 => 2207,
    704 => 2210,
    705 => 2213,
    706 => 2216,
    707 => 2219,
    708 => 2222,
    709 => 2226,
    710 => 2229,
    711 => 2232,
    712 => 2235,
    713 => 2238,
    714 => 2241,
    715 => 2244,
    716 => 2248,
    717 => 2251,
    718 => 2254,
    719 => 2257,
    720 => 2260,
    721 => 2263,
    722 => 2266,
    723 => 2269,
    724 => 2273,
    725 => 2276,
    726 => 2279,
    727 => 2282,
    728 => 2285,
    729 => 2288,
    730 => 2291,
    731 => 2295,
    732 => 2298,
    733 => 2301,
    734 => 2304,
    735 => 2307,
    736 => 2310,
    737 => 2313,
    738 => 2316,
    739 => 2320,
    740 => 2323,
    741 => 2326,
    742 => 2329,
    743 => 2332,
    744 => 2335,
    745 => 2338,
    746 => 2342,
    747 => 2345,
    748 => 2348,
    749 => 2351,
    750 => 2354,
    751 => 2357,
    752 => 2360,
    753 => 2363,
    754 => 2367,
    755 => 2370,
    756 => 2373,
    757 => 2376,
    758 => 2379,
    759 => 2382,
    760 => 2385,
    761 => 2389,
    762 => 2392,
    763 => 2395,
    764 => 2398,
    765 => 2401,
    766 => 2404,
    767 => 2407,
    768 => 2410,
    769 => 2414,
    770 => 2417,
    771 => 2420,
    772 => 2423,
    773 => 2426,
    774 => 2429,
    775 => 2432,
    776 => 2436,
    777 => 2439,
    778 => 2442,
    779 => 2445,
    780 => 2448,
    781 => 2451,
    782 => 2454,
    783 => 2457,
    784 => 2461,
    785 => 2464,
    786 => 2467,
    787 => 2470,
    788 => 2473,
    789 => 2476,
    790 => 2479,
    791 => 2483,
    792 => 2486,
    793 => 2489,
    794 => 2492,
    795 => 2495,
    796 => 2498,
    797 => 2501,
    798 => 2504,
    799 => 2508,
    800 => 2511,
    801 => 2514,
    802 => 2517,
    803 => 2520,
    804 => 2523,
    805 => 2526,
    806 => 2530,
    807 => 2533,
    808 => 2536,
    809 => 2539,
    810 => 2542,
    811 => 2545,
    812 => 2548,
    813 => 2551,
    814 => 2555,
    815 => 2558,
    816 => 2561,
    817 => 2564,
    818 => 2567,
    819 => 2570,
    820 => 2573,
    821 => 2577,
    822 => 2580,
    823 => 2583,
    824 => 2586,
    825 => 2589,
    826 => 2592,
    827 => 2595,
    828 => 2598,
    829 => 2602,
    830 => 2605,
    831 => 2608,
    832 => 2611,
    833 => 2614,
    834 => 2617,
    835 => 2620,
    836 => 2623,
    837 => 2627,
    838 => 2630,
    839 => 2633,
    840 => 2636,
    841 => 2639,
    842 => 2642,
    843 => 2645,
    844 => 2649,
    845 => 2652,
    846 => 2655,
    847 => 2658,
    848 => 2661,
    849 => 2664,
    850 => 2667,
    851 => 2670,
    852 => 2674,
    853 => 2677,
    854 => 2680,
    855 => 2683,
    856 => 2686,
    857 => 2689,
    858 => 2692,
    859 => 2695,
    860 => 2699,
    861 => 2702,
    862 => 2705,
    863 => 2708,
    864 => 2711,
    865 => 2714,
    866 => 2717,
    867 => 2721,
    868 => 2724,
    869 => 2727,
    870 => 2730,
    871 => 2733,
    872 => 2736,
    873 => 2739,
    874 => 2742,
    875 => 2746,
    876 => 2749,
    877 => 2752,
    878 => 2755,
    879 => 2758,
    880 => 2761,
    881 => 2764,
    882 => 2767,
    883 => 2771,
    884 => 2774,
    885 => 2777,
    886 => 2780,
    887 => 2783,
    888 => 2786,
    889 => 2789,
    890 => 2793,
    891 => 2796,
    892 => 2799,
    893 => 2802,
    894 => 2805,
    895 => 2808,
    896 => 2811,
    897 => 2814,
    898 => 2818,
    899 => 2821,
    900 => 2824,
    901 => 2827,
    902 => 2830,
    903 => 2833,
    904 => 2836,
    905 => 2839,
    906 => 2843,
    907 => 2846,
    908 => 2849,
    909 => 2852,
    910 => 2855,
    911 => 2858,
    912 => 2861,
    913 => 2865,
    914 => 2868,
    915 => 2871,
    916 => 2874,
    917 => 2877,
    918 => 2880,
    919 => 2883,
    920 => 2886,
    921 => 2890,
    922 => 2893,
    923 => 2896,
    924 => 2899,
    925 => 2902,
    926 => 2905,
    927 => 2908,
    928 => 2911,
    929 => 2915,
    930 => 2918,
    931 => 2921,
    932 => 2924,
    933 => 2927,
    934 => 2930,
    935 => 2933,
    936 => 2936,
    937 => 2940,
    938 => 2943,
    939 => 2946,
    940 => 2949,
    941 => 2952,
    942 => 2955,
    943 => 2958,
    944 => 2962,
    945 => 2965,
    946 => 2968,
    947 => 2971,
    948 => 2974,
    949 => 2977,
    950 => 2980,
    951 => 2983,
    952 => 2987,
    953 => 2990,
    954 => 2993,
    955 => 2996,
    956 => 2999,
    957 => 3002,
    958 => 3005,
    959 => 3008,
    960 => 3012,
    961 => 3015,
    962 => 3018,
    963 => 3021,
    964 => 3024,
    965 => 3027,
    966 => 3030,
    967 => 3033,
    968 => 3037,
    969 => 3040,
    970 => 3043,
    971 => 3046,
    972 => 3049,
    973 => 3052,
    974 => 3055,
    975 => 3059,
    976 => 3062,
    977 => 3065,
    978 => 3068,
    979 => 3071,
    980 => 3074,
    981 => 3077,
    982 => 3080,
    983 => 3084,
    984 => 3087,
    985 => 3090,
    986 => 3093,
    987 => 3096,
    988 => 3099,
    989 => 3102,
    990 => 3105,
    991 => 3109,
    992 => 3112,
    993 => 3115,
    994 => 3118,
    995 => 3121,
    996 => 3124,
    997 => 3127,
    998 => 3130,
    999 => 3134,
    1000 => 3137,
    1001 => 3140,
    1002 => 3143,
    1003 => 3146,
    1004 => 3149,
    1005 => 3152,
    1006 => 3155,
    1007 => 3159,
    1008 => 3162,
    1009 => 3165,
    1010 => 3168,
    1011 => 3171,
    1012 => 3174,
    1013 => 3177,
    1014 => 3180,
    1015 => 3184,
    1016 => 3187,
    1017 => 3190,
    1018 => 3193,
    1019 => 3196,
    1020 => 3199,
    1021 => 3202,
    1022 => 3205,
    1023 => 3209,
    1024 => 3212,
    1025 => 3215,
    1026 => 3218,
    1027 => 3221,
    1028 => 3224,
    1029 => 3227,
    1030 => 3230,
    1031 => 3234,
    1032 => 3237,
    1033 => 3240,
    1034 => 3243,
    1035 => 3246,
    1036 => 3249,
    1037 => 3252,
    1038 => 3255,
    1039 => 3259,
    1040 => 3262,
    1041 => 3265,
    1042 => 3268,
    1043 => 3271,
    1044 => 3274,
    1045 => 3277,
    1046 => 3281,
    1047 => 3284,
    1048 => 3287,
    1049 => 3290,
    1050 => 3293,
    1051 => 3296,
    1052 => 3299,
    1053 => 3302,
    1054 => 3306,
    1055 => 3309,
    1056 => 3312,
    1057 => 3315,
    1058 => 3318,
    1059 => 3321,
    1060 => 3324,
    1061 => 3327,
    1062 => 3331,
    1063 => 3334,
    1064 => 3337,
    1065 => 3340,
    1066 => 3343,
    1067 => 3346,
    1068 => 3349,
    1069 => 3352,
    1070 => 3356,
    1071 => 3359,
    1072 => 3362,
    1073 => 3365,
    1074 => 3368,
    1075 => 3371,
    1076 => 3374,
    1077 => 3377,
    1078 => 3381,
    1079 => 3384,
    1080 => 3387,
    1081 => 3390,
    1082 => 3393,
    1083 => 3396,
    1084 => 3399,
    1085 => 3402,
    1086 => 3406,
    1087 => 3409,
    1088 => 3412,
    1089 => 3415,
    1090 => 3418,
    1091 => 3421,
    1092 => 3424,
    1093 => 3427,
    1094 => 3430,
    1095 => 3434,
    1096 => 3437,
    1097 => 3440,
    1098 => 3443,
    1099 => 3446,
    1100 => 3449,
    1101 => 3452,
    1102 => 3455,
    1103 => 3459,
    1104 => 3462,
    1105 => 3465,
    1106 => 3468,
    1107 => 3471,
    1108 => 3474,
    1109 => 3477,
    1110 => 3480,
    1111 => 3484,
    1112 => 3487,
    1113 => 3490,
    1114 => 3493,
    1115 => 3496,
    1116 => 3499,
    1117 => 3502,
    1118 => 3505,
    1119 => 3509,
    1120 => 3512,
    1121 => 3515,
    1122 => 3518,
    1123 => 3521,
    1124 => 3524,
    1125 => 3527,
    1126 => 3530,
    1127 => 3534,
    1128 => 3537,
    1129 => 3540,
    1130 => 3543,
    1131 => 3546,
    1132 => 3549,
    1133 => 3552,
    1134 => 3555,
    1135 => 3559,
    1136 => 3562,
    1137 => 3565,
    1138 => 3568,
    1139 => 3571,
    1140 => 3574,
    1141 => 3577,
    1142 => 3580,
    1143 => 3584,
    1144 => 3587,
    1145 => 3590,
    1146 => 3593,
    1147 => 3596,
    1148 => 3599,
    1149 => 3602,
    1150 => 3605,
    1151 => 3609,
    1152 => 3612,
    1153 => 3615,
    1154 => 3618,
    1155 => 3621,
    1156 => 3624,
    1157 => 3627,
    1158 => 3630,
    1159 => 3634,
    1160 => 3637,
    1161 => 3640,
    1162 => 3643,
    1163 => 3646,
    1164 => 3649,
    1165 => 3652,
    1166 => 3655,
    1167 => 3658,
    1168 => 3662,
    1169 => 3665,
    1170 => 3668,
    1171 => 3671,
    1172 => 3674,
    1173 => 3677,
    1174 => 3680,
    1175 => 3683,
    1176 => 3687,
    1177 => 3690,
    1178 => 3693,
    1179 => 3696,
    1180 => 3699,
    1181 => 3702,
    1182 => 3705,
    1183 => 3708,
    1184 => 3712,
    1185 => 3715,
    1186 => 3718,
    1187 => 3721,
    1188 => 3724,
    1189 => 3727,
    1190 => 3730,
    1191 => 3733,
    1192 => 3737,
    1193 => 3740,
    1194 => 3743,
    1195 => 3746,
    1196 => 3749,
    1197 => 3752,
    1198 => 3755,
    1199 => 3758,
    1200 => 3761,
    1201 => 3765,
    1202 => 3768,
    1203 => 3771,
    1204 => 3774,
    1205 => 3777,
    1206 => 3780,
    1207 => 3783,
    1208 => 3786,
    1209 => 3790,
    1210 => 3793,
    1211 => 3796,
    1212 => 3799,
    1213 => 3802,
    1214 => 3805,
    1215 => 3808,
    1216 => 3811,
    1217 => 3815,
    1218 => 3818,
    1219 => 3821,
    1220 => 3824,
    1221 => 3827,
    1222 => 3830,
    1223 => 3833,
    1224 => 3836,
    1225 => 3839,
    1226 => 3843,
    1227 => 3846,
    1228 => 3849,
    1229 => 3852,
    1230 => 3855,
    1231 => 3858,
    1232 => 3861,
    1233 => 3864,
    1234 => 3868,
    1235 => 3871,
    1236 => 3874,
    1237 => 3877,
    1238 => 3880,
    1239 => 3883,
    1240 => 3886,
    1241 => 3889,
    1242 => 3893,
    1243 => 3896,
    1244 => 3899,
    1245 => 3902,
    1246 => 3905,
    1247 => 3908,
    1248 => 3911,
    1249 => 3914,
    1250 => 3917,
    1251 => 3921,
    1252 => 3924,
    1253 => 3927,
    1254 => 3930,
    1255 => 3933,
    1256 => 3936,
    1257 => 3939,
    1258 => 3942,
    1259 => 3946,
    1260 => 3949,
    1261 => 3952,
    1262 => 3955,
    1263 => 3958,
    1264 => 3961,
    1265 => 3964,
    1266 => 3967,
    1267 => 3970,
    1268 => 3974,
    1269 => 3977,
    1270 => 3980,
    1271 => 3983,
    1272 => 3986,
    1273 => 3989,
    1274 => 3992,
    1275 => 3995,
    1276 => 3999,
    1277 => 4002,
    1278 => 4005,
    1279 => 4008,
    1280 => 4011,
    1281 => 4014,
    1282 => 4017,
    1283 => 4020,
    1284 => 4024,
    1285 => 4027,
    1286 => 4030,
    1287 => 4033,
    1288 => 4036,
    1289 => 4039,
    1290 => 4042,
    1291 => 4045,
    1292 => 4048,
    1293 => 4052,
    1294 => 4055,
    1295 => 4058,
    1296 => 4061,
    1297 => 4064,
    1298 => 4067,
    1299 => 4070,
    1300 => 4073,
    1301 => 4076,
    1302 => 4080,
    1303 => 4083,
    1304 => 4086,
    1305 => 4089,
    1306 => 4092,
    1307 => 4095,
    1308 => 4098,
    1309 => 4101,
    1310 => 4105,
    1311 => 4108,
    1312 => 4111,
    1313 => 4114,
    1314 => 4117,
    1315 => 4120,
    1316 => 4123,
    1317 => 4126,
    1318 => 4129,
    1319 => 4133,
    1320 => 4136,
    1321 => 4139,
    1322 => 4142,
    1323 => 4145,
    1324 => 4148,
    1325 => 4151,
    1326 => 4154,
    1327 => 4158,
    1328 => 4161,
    1329 => 4164,
    1330 => 4167,
    1331 => 4170,
    1332 => 4173,
    1333 => 4176,
    1334 => 4179,
    1335 => 4182,
    1336 => 4186,
    1337 => 4189,
    1338 => 4192,
    1339 => 4195,
    1340 => 4198,
    1341 => 4201,
    1342 => 4204,
    1343 => 4207,
    1344 => 4210,
    1345 => 4214,
    1346 => 4217,
    1347 => 4220,
    1348 => 4223,
    1349 => 4226,
    1350 => 4229,
    1351 => 4232,
    1352 => 4235,
    1353 => 4239,
    1354 => 4242,
    1355 => 4245,
    1356 => 4248,
    1357 => 4251,
    1358 => 4254,
    1359 => 4257,
    1360 => 4260,
    1361 => 4263,
    1362 => 4267,
    1363 => 4270,
    1364 => 4273,
    1365 => 4276,
    1366 => 4279,
    1367 => 4282,
    1368 => 4285,
    1369 => 4288,
    1370 => 4291,
    1371 => 4295,
    1372 => 4298,
    1373 => 4301,
    1374 => 4304,
    1375 => 4307,
    1376 => 4310,
    1377 => 4313,
    1378 => 4316,
    1379 => 4320,
    1380 => 4323,
    1381 => 4326,
    1382 => 4329,
    1383 => 4332,
    1384 => 4335,
    1385 => 4338,
    1386 => 4341,
    1387 => 4344,
    1388 => 4348,
    1389 => 4351,
    1390 => 4354,
    1391 => 4357,
    1392 => 4360,
    1393 => 4363,
    1394 => 4366,
    1395 => 4369,
    1396 => 4372,
    1397 => 4376,
    1398 => 4379,
    1399 => 4382,
    1400 => 4385,
    1401 => 4388,
    1402 => 4391,
    1403 => 4394,
    1404 => 4397,
    1405 => 4400,
    1406 => 4404,
    1407 => 4407,
    1408 => 4410,
    1409 => 4413,
    1410 => 4416,
    1411 => 4419,
    1412 => 4422,
    1413 => 4425,
    1414 => 4428,
    1415 => 4432,
    1416 => 4435,
    1417 => 4438,
    1418 => 4441,
    1419 => 4444,
    1420 => 4447,
    1421 => 4450,
    1422 => 4453,
    1423 => 4456,
    1424 => 4460,
    1425 => 4463,
    1426 => 4466,
    1427 => 4469,
    1428 => 4472,
    1429 => 4475,
    1430 => 4478,
    1431 => 4481,
    1432 => 4485,
    1433 => 4488,
    1434 => 4491,
    1435 => 4494,
    1436 => 4497,
    1437 => 4500,
    1438 => 4503,
    1439 => 4506,
    1440 => 4509,
    1441 => 4513,
    1442 => 4516,
    1443 => 4519,
    1444 => 4522,
    1445 => 4525,
    1446 => 4528,
    1447 => 4531,
    1448 => 4534,
    1449 => 4537,
    1450 => 4541,
    1451 => 4544,
    1452 => 4547,
    1453 => 4550,
    1454 => 4553,
    1455 => 4556,
    1456 => 4559,
    1457 => 4562,
    1458 => 4565,
    1459 => 4569,
    1460 => 4572,
    1461 => 4575,
    1462 => 4578,
    1463 => 4581,
    1464 => 4584,
    1465 => 4587,
    1466 => 4590,
    1467 => 4593,
    1468 => 4597,
    1469 => 4600,
    1470 => 4603,
    1471 => 4606,
    1472 => 4609,
    1473 => 4612,
    1474 => 4615,
    1475 => 4618,
    1476 => 4621,
    1477 => 4624,
    1478 => 4628,
    1479 => 4631,
    1480 => 4634,
    1481 => 4637,
    1482 => 4640,
    1483 => 4643,
    1484 => 4646,
    1485 => 4649,
    1486 => 4652,
    1487 => 4656,
    1488 => 4659,
    1489 => 4662,
    1490 => 4665,
    1491 => 4668,
    1492 => 4671,
    1493 => 4674,
    1494 => 4677,
    1495 => 4680,
    1496 => 4684,
    1497 => 4687,
    1498 => 4690,
    1499 => 4693,
    1500 => 4696,
    1501 => 4699,
    1502 => 4702,
    1503 => 4705,
    1504 => 4708,
    1505 => 4712,
    1506 => 4715,
    1507 => 4718,
    1508 => 4721,
    1509 => 4724,
    1510 => 4727,
    1511 => 4730,
    1512 => 4733,
    1513 => 4736,
    1514 => 4740,
    1515 => 4743,
    1516 => 4746,
    1517 => 4749,
    1518 => 4752,
    1519 => 4755,
    1520 => 4758,
    1521 => 4761,
    1522 => 4764,
    1523 => 4768,
    1524 => 4771,
    1525 => 4774,
    1526 => 4777,
    1527 => 4780,
    1528 => 4783,
    1529 => 4786,
    1530 => 4789,
    1531 => 4792,
    1532 => 4795,
    1533 => 4799,
    1534 => 4802,
    1535 => 4805,
    1536 => 4808,
    1537 => 4811,
    1538 => 4814,
    1539 => 4817,
    1540 => 4820,
    1541 => 4823,
    1542 => 4827,
    1543 => 4830,
    1544 => 4833,
    1545 => 4836,
    1546 => 4839,
    1547 => 4842,
    1548 => 4845,
    1549 => 4848,
    1550 => 4851,
    1551 => 4855,
    1552 => 4858,
    1553 => 4861,
    1554 => 4864,
    1555 => 4867,
    1556 => 4870,
    1557 => 4873,
    1558 => 4876,
    1559 => 4879,
    1560 => 4882,
    1561 => 4886,
    1562 => 4889,
    1563 => 4892,
    1564 => 4895,
    1565 => 4898,
    1566 => 4901,
    1567 => 4904,
    1568 => 4907,
    1569 => 4910,
    1570 => 4914,
    1571 => 4917,
    1572 => 4920,
    1573 => 4923,
    1574 => 4926,
    1575 => 4929,
    1576 => 4932,
    1577 => 4935,
    1578 => 4938,
    1579 => 4941,
    1580 => 4945,
    1581 => 4948,
    1582 => 4951,
    1583 => 4954,
    1584 => 4957,
    1585 => 4960,
    1586 => 4963,
    1587 => 4966,
    1588 => 4969,
    1589 => 4973,
    1590 => 4976,
    1591 => 4979,
    1592 => 4982,
    1593 => 4985,
    1594 => 4988,
    1595 => 4991,
    1596 => 4994,
    1597 => 4997,
    1598 => 5000,
    1599 => 5004,
    1600 => 5007,
    1601 => 5010,
    1602 => 5013,
    1603 => 5016,
    1604 => 5019,
    1605 => 5022,
    1606 => 5025,
    1607 => 5028,
    1608 => 5032,
    1609 => 5035,
    1610 => 5038,
    1611 => 5041,
    1612 => 5044,
    1613 => 5047,
    1614 => 5050,
    1615 => 5053,
    1616 => 5056,
    1617 => 5059,
    1618 => 5063,
    1619 => 5066,
    1620 => 5069,
    1621 => 5072,
    1622 => 5075,
    1623 => 5078,
    1624 => 5081,
    1625 => 5084,
    1626 => 5087,
    1627 => 5091,
    1628 => 5094,
    1629 => 5097,
    1630 => 5100,
    1631 => 5103,
    1632 => 5106,
    1633 => 5109,
    1634 => 5112,
    1635 => 5115,
    1636 => 5118,
    1637 => 5122,
    1638 => 5125,
    1639 => 5128,
    1640 => 5131,
    1641 => 5134,
    1642 => 5137,
    1643 => 5140,
    1644 => 5143,
    1645 => 5146,
    1646 => 5149,
    1647 => 5153,
    1648 => 5156,
    1649 => 5159,
    1650 => 5162,
    1651 => 5165,
    1652 => 5168,
    1653 => 5171,
    1654 => 5174,
    1655 => 5177,
    1656 => 5180,
    1657 => 5184,
    1658 => 5187,
    1659 => 5190,
    1660 => 5193,
    1661 => 5196,
    1662 => 5199,
    1663 => 5202,
    1664 => 5205,
    1665 => 5208,
    1666 => 5212,
    1667 => 5215,
    1668 => 5218,
    1669 => 5221,
    1670 => 5224,
    1671 => 5227,
    1672 => 5230,
    1673 => 5233,
    1674 => 5236,
    1675 => 5239,
    1676 => 5243,
    1677 => 5246,
    1678 => 5249,
    1679 => 5252,
    1680 => 5255,
    1681 => 5258,
    1682 => 5261,
    1683 => 5264,
    1684 => 5267,
    1685 => 5270,
    1686 => 5274,
    1687 => 5277,
    1688 => 5280,
    1689 => 5283,
    1690 => 5286,
    1691 => 5289,
    1692 => 5292,
    1693 => 5295,
    1694 => 5298,
    1695 => 5301,
    1696 => 5305,
    1697 => 5308,
    1698 => 5311,
    1699 => 5314,
    1700 => 5317,
    1701 => 5320,
    1702 => 5323,
    1703 => 5326,
    1704 => 5329,
    1705 => 5332,
    1706 => 5336,
    1707 => 5339,
    1708 => 5342,
    1709 => 5345,
    1710 => 5348,
    1711 => 5351,
    1712 => 5354,
    1713 => 5357,
    1714 => 5360,
    1715 => 5363,
    1716 => 5367,
    1717 => 5370,
    1718 => 5373,
    1719 => 5376,
    1720 => 5379,
    1721 => 5382,
    1722 => 5385,
    1723 => 5388,
    1724 => 5391,
    1725 => 5394,
    1726 => 5398,
    1727 => 5401,
    1728 => 5404,
    1729 => 5407,
    1730 => 5410,
    1731 => 5413,
    1732 => 5416,
    1733 => 5419,
    1734 => 5422,
    1735 => 5425,
    1736 => 5428,
    1737 => 5432,
    1738 => 5435,
    1739 => 5438,
    1740 => 5441,
    1741 => 5444,
    1742 => 5447,
    1743 => 5450,
    1744 => 5453,
    1745 => 5456,
    1746 => 5459,
    1747 => 5463,
    1748 => 5466,
    1749 => 5469,
    1750 => 5472,
    1751 => 5475,
    1752 => 5478,
    1753 => 5481,
    1754 => 5484,
    1755 => 5487,
    1756 => 5490,
    1757 => 5494,
    1758 => 5497,
    1759 => 5500,
    1760 => 5503,
    1761 => 5506,
    1762 => 5509,
    1763 => 5512,
    1764 => 5515,
    1765 => 5518,
    1766 => 5521,
    1767 => 5525,
    1768 => 5528,
    1769 => 5531,
    1770 => 5534,
    1771 => 5537,
    1772 => 5540,
    1773 => 5543,
    1774 => 5546,
    1775 => 5549,
    1776 => 5552,
    1777 => 5555,
    1778 => 5559,
    1779 => 5562,
    1780 => 5565,
    1781 => 5568,
    1782 => 5571,
    1783 => 5574,
    1784 => 5577,
    1785 => 5580,
    1786 => 5583,
    1787 => 5586,
    1788 => 5590,
    1789 => 5593,
    1790 => 5596,
    1791 => 5599,
    1792 => 5602,
    1793 => 5605,
    1794 => 5608,
    1795 => 5611,
    1796 => 5614,
    1797 => 5617,
    1798 => 5620,
    1799 => 5624,
    1800 => 5627,
    1801 => 5630,
    1802 => 5633,
    1803 => 5636,
    1804 => 5639,
    1805 => 5642,
    1806 => 5645,
    1807 => 5648,
    1808 => 5651,
    1809 => 5655,
    1810 => 5658,
    1811 => 5661,
    1812 => 5664,
    1813 => 5667,
    1814 => 5670,
    1815 => 5673,
    1816 => 5676,
    1817 => 5679,
    1818 => 5682,
    1819 => 5685,
    1820 => 5689,
    1821 => 5692,
    1822 => 5695,
    1823 => 5698,
    1824 => 5701,
    1825 => 5704,
    1826 => 5707,
    1827 => 5710,
    1828 => 5713,
    1829 => 5716,
    1830 => 5719,
    1831 => 5723,
    1832 => 5726,
    1833 => 5729,
    1834 => 5732,
    1835 => 5735,
    1836 => 5738,
    1837 => 5741,
    1838 => 5744,
    1839 => 5747,
    1840 => 5750,
    1841 => 5754,
    1842 => 5757,
    1843 => 5760,
    1844 => 5763,
    1845 => 5766,
    1846 => 5769,
    1847 => 5772,
    1848 => 5775,
    1849 => 5778,
    1850 => 5781,
    1851 => 5784,
    1852 => 5788,
    1853 => 5791,
    1854 => 5794,
    1855 => 5797,
    1856 => 5800,
    1857 => 5803,
    1858 => 5806,
    1859 => 5809,
    1860 => 5812,
    1861 => 5815,
    1862 => 5818,
    1863 => 5822,
    1864 => 5825,
    1865 => 5828,
    1866 => 5831,
    1867 => 5834,
    1868 => 5837,
    1869 => 5840,
    1870 => 5843,
    1871 => 5846,
    1872 => 5849,
    1873 => 5852,
    1874 => 5856,
    1875 => 5859,
    1876 => 5862,
    1877 => 5865,
    1878 => 5868,
    1879 => 5871,
    1880 => 5874,
    1881 => 5877,
    1882 => 5880,
    1883 => 5883,
    1884 => 5886,
    1885 => 5890,
    1886 => 5893,
    1887 => 5896,
    1888 => 5899,
    1889 => 5902,
    1890 => 5905,
    1891 => 5908,
    1892 => 5911,
    1893 => 5914,
    1894 => 5917,
    1895 => 5920,
    1896 => 5924,
    1897 => 5927,
    1898 => 5930,
    1899 => 5933,
    1900 => 5936,
    1901 => 5939,
    1902 => 5942,
    1903 => 5945,
    1904 => 5948,
    1905 => 5951,
    1906 => 5954,
    1907 => 5958,
    1908 => 5961,
    1909 => 5964,
    1910 => 5967,
    1911 => 5970,
    1912 => 5973,
    1913 => 5976,
    1914 => 5979,
    1915 => 5982,
    1916 => 5985,
    1917 => 5988,
    1918 => 5991,
    1919 => 5995,
    1920 => 5998,
    1921 => 6001,
    1922 => 6004,
    1923 => 6007,
    1924 => 6010,
    1925 => 6013,
    1926 => 6016,
    1927 => 6019,
    1928 => 6022,
    1929 => 6025,
    1930 => 6029,
    1931 => 6032,
    1932 => 6035,
    1933 => 6038,
    1934 => 6041,
    1935 => 6044,
    1936 => 6047,
    1937 => 6050,
    1938 => 6053,
    1939 => 6056,
    1940 => 6059,
    1941 => 6063,
    1942 => 6066,
    1943 => 6069,
    1944 => 6072,
    1945 => 6075,
    1946 => 6078,
    1947 => 6081,
    1948 => 6084,
    1949 => 6087,
    1950 => 6090,
    1951 => 6093,
    1952 => 6096,
    1953 => 6100,
    1954 => 6103,
    1955 => 6106,
    1956 => 6109,
    1957 => 6112,
    1958 => 6115,
    1959 => 6118,
    1960 => 6121,
    1961 => 6124,
    1962 => 6127,
    1963 => 6130,
    1964 => 6134,
    1965 => 6137,
    1966 => 6140,
    1967 => 6143,
    1968 => 6146,
    1969 => 6149,
    1970 => 6152,
    1971 => 6155,
    1972 => 6158,
    1973 => 6161,
    1974 => 6164,
    1975 => 6167,
    1976 => 6171,
    1977 => 6174,
    1978 => 6177,
    1979 => 6180,
    1980 => 6183,
    1981 => 6186,
    1982 => 6189,
    1983 => 6192,
    1984 => 6195,
    1985 => 6198,
    1986 => 6201,
    1987 => 6204,
    1988 => 6208,
    1989 => 6211,
    1990 => 6214,
    1991 => 6217,
    1992 => 6220,
    1993 => 6223,
    1994 => 6226,
    1995 => 6229,
    1996 => 6232,
    1997 => 6235,
    1998 => 6238,
    1999 => 6241,
    2000 => 6245,
    2001 => 6248,
    2002 => 6251,
    2003 => 6254,
    2004 => 6257,
    2005 => 6260,
    2006 => 6263,
    2007 => 6266,
    2008 => 6269,
    2009 => 6272,
    2010 => 6275,
    2011 => 6278,
    2012 => 6282,
    2013 => 6285,
    2014 => 6288,
    2015 => 6291,
    2016 => 6294,
    2017 => 6297,
    2018 => 6300,
    2019 => 6303,
    2020 => 6306,
    2021 => 6309,
    2022 => 6312,
    2023 => 6315,
    2024 => 6319,
    2025 => 6322,
    2026 => 6325,
    2027 => 6328,
    2028 => 6331,
    2029 => 6334,
    2030 => 6337,
    2031 => 6340,
    2032 => 6343,
    2033 => 6346,
    2034 => 6349,
    2035 => 6352,
    2036 => 6356,
    2037 => 6359,
    2038 => 6362,
    2039 => 6365,
    2040 => 6368,
    2041 => 6371,
    2042 => 6374,
    2043 => 6377,
    2044 => 6380,
    2045 => 6383,
    2046 => 6386,
    2047 => 6389,
    2048 => 6393,
    2049 => 6396,
    2050 => 6399,
    2051 => 6402,
    2052 => 6405,
    2053 => 6408,
    2054 => 6411,
    2055 => 6414,
    2056 => 6417,
    2057 => 6420,
    2058 => 6423,
    2059 => 6426,
    2060 => 6429,
    2061 => 6433,
    2062 => 6436,
    2063 => 6439,
    2064 => 6442,
    2065 => 6445,
    2066 => 6448,
    2067 => 6451,
    2068 => 6454,
    2069 => 6457,
    2070 => 6460,
    2071 => 6463,
    2072 => 6466,
    2073 => 6470,
    2074 => 6473,
    2075 => 6476,
    2076 => 6479,
    2077 => 6482,
    2078 => 6485,
    2079 => 6488,
    2080 => 6491,
    2081 => 6494,
    2082 => 6497,
    2083 => 6500,
    2084 => 6503,
    2085 => 6506,
    2086 => 6510,
    2087 => 6513,
    2088 => 6516,
    2089 => 6519,
    2090 => 6522,
    2091 => 6525,
    2092 => 6528,
    2093 => 6531,
    2094 => 6534,
    2095 => 6537,
    2096 => 6540,
    2097 => 6543,
    2098 => 6547,
    2099 => 6550,
    2100 => 6553,
    2101 => 6556,
    2102 => 6559,
    2103 => 6562,
    2104 => 6565,
    2105 => 6568,
    2106 => 6571,
    2107 => 6574,
    2108 => 6577,
    2109 => 6580,
    2110 => 6583,
    2111 => 6587,
    2112 => 6590,
    2113 => 6593,
    2114 => 6596,
    2115 => 6599,
    2116 => 6602,
    2117 => 6605,
    2118 => 6608,
    2119 => 6611,
    2120 => 6614,
    2121 => 6617,
    2122 => 6620,
    2123 => 6623,
    2124 => 6627,
    2125 => 6630,
    2126 => 6633,
    2127 => 6636,
    2128 => 6639,
    2129 => 6642,
    2130 => 6645,
    2131 => 6648,
    2132 => 6651,
    2133 => 6654,
    2134 => 6657,
    2135 => 6660,
    2136 => 6663,
    2137 => 6667,
    2138 => 6670,
    2139 => 6673,
    2140 => 6676,
    2141 => 6679,
    2142 => 6682,
    2143 => 6685,
    2144 => 6688,
    2145 => 6691,
    2146 => 6694,
    2147 => 6697,
    2148 => 6700,
    2149 => 6703,
    2150 => 6706,
    2151 => 6710,
    2152 => 6713,
    2153 => 6716,
    2154 => 6719,
    2155 => 6722,
    2156 => 6725,
    2157 => 6728,
    2158 => 6731,
    2159 => 6734,
    2160 => 6737,
    2161 => 6740,
    2162 => 6743,
    2163 => 6746,
    2164 => 6750,
    2165 => 6753,
    2166 => 6756,
    2167 => 6759,
    2168 => 6762,
    2169 => 6765,
    2170 => 6768,
    2171 => 6771,
    2172 => 6774,
    2173 => 6777,
    2174 => 6780,
    2175 => 6783,
    2176 => 6786,
    2177 => 6789,
    2178 => 6793,
    2179 => 6796,
    2180 => 6799,
    2181 => 6802,
    2182 => 6805,
    2183 => 6808,
    2184 => 6811,
    2185 => 6814,
    2186 => 6817,
    2187 => 6820,
    2188 => 6823,
    2189 => 6826,
    2190 => 6829,
    2191 => 6833,
    2192 => 6836,
    2193 => 6839,
    2194 => 6842,
    2195 => 6845,
    2196 => 6848,
    2197 => 6851,
    2198 => 6854,
    2199 => 6857,
    2200 => 6860,
    2201 => 6863,
    2202 => 6866,
    2203 => 6869,
    2204 => 6872,
    2205 => 6876,
    2206 => 6879,
    2207 => 6882,
    2208 => 6885,
    2209 => 6888,
    2210 => 6891,
    2211 => 6894,
    2212 => 6897,
    2213 => 6900,
    2214 => 6903,
    2215 => 6906,
    2216 => 6909,
    2217 => 6912,
    2218 => 6915,
    2219 => 6919,
    2220 => 6922,
    2221 => 6925,
    2222 => 6928,
    2223 => 6931,
    2224 => 6934,
    2225 => 6937,
    2226 => 6940,
    2227 => 6943,
    2228 => 6946,
    2229 => 6949,
    2230 => 6952,
    2231 => 6955,
    2232 => 6958,
    2233 => 6961,
    2234 => 6965,
    2235 => 6968,
    2236 => 6971,
    2237 => 6974,
    2238 => 6977,
    2239 => 6980,
    2240 => 6983,
    2241 => 6986,
    2242 => 6989,
    2243 => 6992,
    2244 => 6995,
    2245 => 6998,
    2246 => 7001,
    2247 => 7004,
    2248 => 7008,
    2249 => 7011,
    2250 => 7014,
    2251 => 7017,
    2252 => 7020,
    2253 => 7023,
    2254 => 7026,
    2255 => 7029,
    2256 => 7032,
    2257 => 7035,
    2258 => 7038,
    2259 => 7041,
    2260 => 7044,
    2261 => 7047,
    2262 => 7050,
    2263 => 7054,
    2264 => 7057,
    2265 => 7060,
    2266 => 7063,
    2267 => 7066,
    2268 => 7069,
    2269 => 7072,
    2270 => 7075,
    2271 => 7078,
    2272 => 7081,
    2273 => 7084,
    2274 => 7087,
    2275 => 7090,
    2276 => 7093,
    2277 => 7097,
    2278 => 7100,
    2279 => 7103,
    2280 => 7106,
    2281 => 7109,
    2282 => 7112,
    2283 => 7115,
    2284 => 7118,
    2285 => 7121,
    2286 => 7124,
    2287 => 7127,
    2288 => 7130,
    2289 => 7133,
    2290 => 7136,
    2291 => 7139,
    2292 => 7143,
    2293 => 7146,
    2294 => 7149,
    2295 => 7152,
    2296 => 7155,
    2297 => 7158,
    2298 => 7161,
    2299 => 7164,
    2300 => 7167,
    2301 => 7170,
    2302 => 7173,
    2303 => 7176,
    2304 => 7179,
    2305 => 7182,
    2306 => 7185,
    2307 => 7188,
    2308 => 7192,
    2309 => 7195,
    2310 => 7198,
    2311 => 7201,
    2312 => 7204,
    2313 => 7207,
    2314 => 7210,
    2315 => 7213,
    2316 => 7216,
    2317 => 7219,
    2318 => 7222,
    2319 => 7225,
    2320 => 7228,
    2321 => 7231,
    2322 => 7234,
    2323 => 7238,
    2324 => 7241,
    2325 => 7244,
    2326 => 7247,
    2327 => 7250,
    2328 => 7253,
    2329 => 7256,
    2330 => 7259,
    2331 => 7262,
    2332 => 7265,
    2333 => 7268,
    2334 => 7271,
    2335 => 7274,
    2336 => 7277,
    2337 => 7280,
    2338 => 7283,
    2339 => 7287,
    2340 => 7290,
    2341 => 7293,
    2342 => 7296,
    2343 => 7299,
    2344 => 7302,
    2345 => 7305,
    2346 => 7308,
    2347 => 7311,
    2348 => 7314,
    2349 => 7317,
    2350 => 7320,
    2351 => 7323,
    2352 => 7326,
    2353 => 7329,
    2354 => 7332,
    2355 => 7336,
    2356 => 7339,
    2357 => 7342,
    2358 => 7345,
    2359 => 7348,
    2360 => 7351,
    2361 => 7354,
    2362 => 7357,
    2363 => 7360,
    2364 => 7363,
    2365 => 7366,
    2366 => 7369,
    2367 => 7372,
    2368 => 7375,
    2369 => 7378,
    2370 => 7381,
    2371 => 7385,
    2372 => 7388,
    2373 => 7391,
    2374 => 7394,
    2375 => 7397,
    2376 => 7400,
    2377 => 7403,
    2378 => 7406,
    2379 => 7409,
    2380 => 7412,
    2381 => 7415,
    2382 => 7418,
    2383 => 7421,
    2384 => 7424,
    2385 => 7427,
    2386 => 7430,
    2387 => 7433,
    2388 => 7437,
    2389 => 7440,
    2390 => 7443,
    2391 => 7446,
    2392 => 7449,
    2393 => 7452,
    2394 => 7455,
    2395 => 7458,
    2396 => 7461,
    2397 => 7464,
    2398 => 7467,
    2399 => 7470,
    2400 => 7473,
    2401 => 7476,
    2402 => 7479,
    2403 => 7482,
    2404 => 7485,
    2405 => 7489,
    2406 => 7492,
    2407 => 7495,
    2408 => 7498,
    2409 => 7501,
    2410 => 7504,
    2411 => 7507,
    2412 => 7510,
    2413 => 7513,
    2414 => 7516,
    2415 => 7519,
    2416 => 7522,
    2417 => 7525,
    2418 => 7528,
    2419 => 7531,
    2420 => 7534,
    2421 => 7537,
    2422 => 7541,
    2423 => 7544,
    2424 => 7547,
    2425 => 7550,
    2426 => 7553,
    2427 => 7556,
    2428 => 7559,
    2429 => 7562,
    2430 => 7565,
    2431 => 7568,
    2432 => 7571,
    2433 => 7574,
    2434 => 7577,
    2435 => 7580,
    2436 => 7583,
    2437 => 7586,
    2438 => 7589,
    2439 => 7592,
    2440 => 7596,
    2441 => 7599,
    2442 => 7602,
    2443 => 7605,
    2444 => 7608,
    2445 => 7611,
    2446 => 7614,
    2447 => 7617,
    2448 => 7620,
    2449 => 7623,
    2450 => 7626,
    2451 => 7629,
    2452 => 7632,
    2453 => 7635,
    2454 => 7638,
    2455 => 7641,
    2456 => 7644,
    2457 => 7647,
    2458 => 7651,
    2459 => 7654,
    2460 => 7657,
    2461 => 7660,
    2462 => 7663,
    2463 => 7666,
    2464 => 7669,
    2465 => 7672,
    2466 => 7675,
    2467 => 7678,
    2468 => 7681,
    2469 => 7684,
    2470 => 7687,
    2471 => 7690,
    2472 => 7693,
    2473 => 7696,
    2474 => 7699,
    2475 => 7702,
    2476 => 7705,
    2477 => 7709,
    2478 => 7712,
    2479 => 7715,
    2480 => 7718,
    2481 => 7721,
    2482 => 7724,
    2483 => 7727,
    2484 => 7730,
    2485 => 7733,
    2486 => 7736,
    2487 => 7739,
    2488 => 7742,
    2489 => 7745,
    2490 => 7748,
    2491 => 7751,
    2492 => 7754,
    2493 => 7757,
    2494 => 7760,
    2495 => 7764,
    2496 => 7767,
    2497 => 7770,
    2498 => 7773,
    2499 => 7776,
    2500 => 7779,
    2501 => 7782,
    2502 => 7785,
    2503 => 7788,
    2504 => 7791,
    2505 => 7794,
    2506 => 7797,
    2507 => 7800,
    2508 => 7803,
    2509 => 7806,
    2510 => 7809,
    2511 => 7812,
    2512 => 7815,
    2513 => 7818,
    2514 => 7821,
    2515 => 7825,
    2516 => 7828,
    2517 => 7831,
    2518 => 7834,
    2519 => 7837,
    2520 => 7840,
    2521 => 7843,
    2522 => 7846,
    2523 => 7849,
    2524 => 7852,
    2525 => 7855,
    2526 => 7858,
    2527 => 7861,
    2528 => 7864,
    2529 => 7867,
    2530 => 7870,
    2531 => 7873,
    2532 => 7876,
    2533 => 7879,
    2534 => 7882,
    2535 => 7886,
    2536 => 7889,
    2537 => 7892,
    2538 => 7895,
    2539 => 7898,
    2540 => 7901,
    2541 => 7904,
    2542 => 7907,
    2543 => 7910,
    2544 => 7913,
    2545 => 7916,
    2546 => 7919,
    2547 => 7922,
    2548 => 7925,
    2549 => 7928,
    2550 => 7931,
    2551 => 7934,
    2552 => 7937,
    2553 => 7940,
    2554 => 7943,
    2555 => 7946,
    2556 => 7950,
    2557 => 7953,
    2558 => 7956,
    2559 => 7959,
    2560 => 7962,
    2561 => 7965,
    2562 => 7968,
    2563 => 7971,
    2564 => 7974,
    2565 => 7977,
    2566 => 7980,
    2567 => 7983,
    2568 => 7986,
    2569 => 7989,
    2570 => 7992,
    2571 => 7995,
    2572 => 7998,
    2573 => 8001,
    2574 => 8004,
    2575 => 8007,
    2576 => 8010,
    2577 => 8014,
    2578 => 8017,
    2579 => 8020,
    2580 => 8023,
    2581 => 8026,
    2582 => 8029,
    2583 => 8032,
    2584 => 8035,
    2585 => 8038,
    2586 => 8041,
    2587 => 8044,
    2588 => 8047,
    2589 => 8050,
    2590 => 8053,
    2591 => 8056,
    2592 => 8059,
    2593 => 8062,
    2594 => 8065,
    2595 => 8068,
    2596 => 8071,
    2597 => 8074,
    2598 => 8077,
    2599 => 8081,
    2600 => 8084,
    2601 => 8087,
    2602 => 8090,
    2603 => 8093,
    2604 => 8096,
    2605 => 8099,
    2606 => 8102,
    2607 => 8105,
    2608 => 8108,
    2609 => 8111,
    2610 => 8114,
    2611 => 8117,
    2612 => 8120,
    2613 => 8123,
    2614 => 8126,
    2615 => 8129,
    2616 => 8132,
    2617 => 8135,
    2618 => 8138,
    2619 => 8141,
    2620 => 8144,
    2621 => 8147,
    2622 => 8151,
    2623 => 8154,
    2624 => 8157,
    2625 => 8160,
    2626 => 8163,
    2627 => 8166,
    2628 => 8169,
    2629 => 8172,
    2630 => 8175,
    2631 => 8178,
    2632 => 8181,
    2633 => 8184,
    2634 => 8187,
    2635 => 8190,
    2636 => 8193,
    2637 => 8196,
    2638 => 8199,
    2639 => 8202,
    2640 => 8205,
    2641 => 8208,
    2642 => 8211,
    2643 => 8214,
    2644 => 8217,
    2645 => 8220,
    2646 => 8224,
    2647 => 8227,
    2648 => 8230,
    2649 => 8233,
    2650 => 8236,
    2651 => 8239,
    2652 => 8242,
    2653 => 8245,
    2654 => 8248,
    2655 => 8251,
    2656 => 8254,
    2657 => 8257,
    2658 => 8260,
    2659 => 8263,
    2660 => 8266,
    2661 => 8269,
    2662 => 8272,
    2663 => 8275,
    2664 => 8278,
    2665 => 8281,
    2666 => 8284,
    2667 => 8287,
    2668 => 8290,
    2669 => 8293,
    2670 => 8296,
    2671 => 8300,
    2672 => 8303,
    2673 => 8306,
    2674 => 8309,
    2675 => 8312,
    2676 => 8315,
    2677 => 8318,
    2678 => 8321,
    2679 => 8324,
    2680 => 8327,
    2681 => 8330,
    2682 => 8333,
    2683 => 8336,
    2684 => 8339,
    2685 => 8342,
    2686 => 8345,
    2687 => 8348,
    2688 => 8351,
    2689 => 8354,
    2690 => 8357,
    2691 => 8360,
    2692 => 8363,
    2693 => 8366,
    2694 => 8369,
    2695 => 8372,
    2696 => 8375,
    2697 => 8379,
    2698 => 8382,
    2699 => 8385,
    2700 => 8388,
    2701 => 8391,
    2702 => 8394,
    2703 => 8397,
    2704 => 8400,
    2705 => 8403,
    2706 => 8406,
    2707 => 8409,
    2708 => 8412,
    2709 => 8415,
    2710 => 8418,
    2711 => 8421,
    2712 => 8424,
    2713 => 8427,
    2714 => 8430,
    2715 => 8433,
    2716 => 8436,
    2717 => 8439,
    2718 => 8442,
    2719 => 8445,
    2720 => 8448,
    2721 => 8451,
    2722 => 8454,
    2723 => 8457,
    2724 => 8460,
    2725 => 8464,
    2726 => 8467,
    2727 => 8470,
    2728 => 8473,
    2729 => 8476,
    2730 => 8479,
    2731 => 8482,
    2732 => 8485,
    2733 => 8488,
    2734 => 8491,
    2735 => 8494,
    2736 => 8497,
    2737 => 8500,
    2738 => 8503,
    2739 => 8506,
    2740 => 8509,
    2741 => 8512,
    2742 => 8515,
    2743 => 8518,
    2744 => 8521,
    2745 => 8524,
    2746 => 8527,
    2747 => 8530,
    2748 => 8533,
    2749 => 8536,
    2750 => 8539,
    2751 => 8542,
    2752 => 8545,
    2753 => 8548,
    2754 => 8552,
    2755 => 8555,
    2756 => 8558,
    2757 => 8561,
    2758 => 8564,
    2759 => 8567,
    2760 => 8570,
    2761 => 8573,
    2762 => 8576,
    2763 => 8579,
    2764 => 8582,
    2765 => 8585,
    2766 => 8588,
    2767 => 8591,
    2768 => 8594,
    2769 => 8597,
    2770 => 8600,
    2771 => 8603,
    2772 => 8606,
    2773 => 8609,
    2774 => 8612,
    2775 => 8615,
    2776 => 8618,
    2777 => 8621,
    2778 => 8624,
    2779 => 8627,
    2780 => 8630,
    2781 => 8633,
    2782 => 8636,
    2783 => 8639,
    2784 => 8642,
    2785 => 8645,
    2786 => 8649,
    2787 => 8652,
    2788 => 8655,
    2789 => 8658,
    2790 => 8661,
    2791 => 8664,
    2792 => 8667,
    2793 => 8670,
    2794 => 8673,
    2795 => 8676,
    2796 => 8679,
    2797 => 8682,
    2798 => 8685,
    2799 => 8688,
    2800 => 8691,
    2801 => 8694,
    2802 => 8697,
    2803 => 8700,
    2804 => 8703,
    2805 => 8706,
    2806 => 8709,
    2807 => 8712,
    2808 => 8715,
    2809 => 8718,
    2810 => 8721,
    2811 => 8724,
    2812 => 8727,
    2813 => 8730,
    2814 => 8733,
    2815 => 8736,
    2816 => 8739,
    2817 => 8742,
    2818 => 8745,
    2819 => 8748,
    2820 => 8751,
    2821 => 8755,
    2822 => 8758,
    2823 => 8761,
    2824 => 8764,
    2825 => 8767,
    2826 => 8770,
    2827 => 8773,
    2828 => 8776,
    2829 => 8779,
    2830 => 8782,
    2831 => 8785,
    2832 => 8788,
    2833 => 8791,
    2834 => 8794,
    2835 => 8797,
    2836 => 8800,
    2837 => 8803,
    2838 => 8806,
    2839 => 8809,
    2840 => 8812,
    2841 => 8815,
    2842 => 8818,
    2843 => 8821,
    2844 => 8824,
    2845 => 8827,
    2846 => 8830,
    2847 => 8833,
    2848 => 8836,
    2849 => 8839,
    2850 => 8842,
    2851 => 8845,
    2852 => 8848,
    2853 => 8851,
    2854 => 8854,
    2855 => 8857,
    2856 => 8860,
    2857 => 8863,
    2858 => 8866,
    2859 => 8869,
    2860 => 8873,
    2861 => 8876,
    2862 => 8879,
    2863 => 8882,
    2864 => 8885,
    2865 => 8888,
    2866 => 8891,
    2867 => 8894,
    2868 => 8897,
    2869 => 8900,
    2870 => 8903,
    2871 => 8906,
    2872 => 8909,
    2873 => 8912,
    2874 => 8915,
    2875 => 8918,
    2876 => 8921,
    2877 => 8924,
    2878 => 8927,
    2879 => 8930,
    2880 => 8933,
    2881 => 8936,
    2882 => 8939,
    2883 => 8942,
    2884 => 8945,
    2885 => 8948,
    2886 => 8951,
    2887 => 8954,
    2888 => 8957,
    2889 => 8960,
    2890 => 8963,
    2891 => 8966,
    2892 => 8969,
    2893 => 8972,
    2894 => 8975,
    2895 => 8978,
    2896 => 8981,
    2897 => 8984,
    2898 => 8987,
    2899 => 8990,
    2900 => 8993,
    2901 => 8996,
    2902 => 8999,
    2903 => 9002,
    2904 => 9006,
    2905 => 9009,
    2906 => 9012,
    2907 => 9015,
    2908 => 9018,
    2909 => 9021,
    2910 => 9024,
    2911 => 9027,
    2912 => 9030,
    2913 => 9033,
    2914 => 9036,
    2915 => 9039,
    2916 => 9042,
    2917 => 9045,
    2918 => 9048,
    2919 => 9051,
    2920 => 9054,
    2921 => 9057,
    2922 => 9060,
    2923 => 9063,
    2924 => 9066,
    2925 => 9069,
    2926 => 9072,
    2927 => 9075,
    2928 => 9078,
    2929 => 9081,
    2930 => 9084,
    2931 => 9087,
    2932 => 9090,
    2933 => 9093,
    2934 => 9096,
    2935 => 9099,
    2936 => 9102,
    2937 => 9105,
    2938 => 9108,
    2939 => 9111,
    2940 => 9114,
    2941 => 9117,
    2942 => 9120,
    2943 => 9123,
    2944 => 9126,
    2945 => 9129,
    2946 => 9132,
    2947 => 9135,
    2948 => 9138,
    2949 => 9141,
    2950 => 9144,
    2951 => 9147,
    2952 => 9150,
    2953 => 9153,
    2954 => 9156,
    2955 => 9159,
    2956 => 9162,
    2957 => 9165,
    2958 => 9168,
    2959 => 9172,
    2960 => 9175,
    2961 => 9178,
    2962 => 9181,
    2963 => 9184,
    2964 => 9187,
    2965 => 9190,
    2966 => 9193,
    2967 => 9196,
    2968 => 9199,
    2969 => 9202,
    2970 => 9205,
    2971 => 9208,
    2972 => 9211,
    2973 => 9214,
    2974 => 9217,
    2975 => 9220,
    2976 => 9223,
    2977 => 9226,
    2978 => 9229,
    2979 => 9232,
    2980 => 9235,
    2981 => 9238,
    2982 => 9241,
    2983 => 9244,
    2984 => 9247,
    2985 => 9250,
    2986 => 9253,
    2987 => 9256,
    2988 => 9259,
    2989 => 9262,
    2990 => 9265,
    2991 => 9268,
    2992 => 9271,
    2993 => 9274,
    2994 => 9277,
    2995 => 9280,
    2996 => 9283,
    2997 => 9286,
    2998 => 9289,
    2999 => 9292,
    3000 => 9295,
    3001 => 9298,
    3002 => 9301,
    3003 => 9304,
    3004 => 9307,
    3005 => 9310,
    3006 => 9313,
    3007 => 9316,
    3008 => 9319,
    3009 => 9322,
    3010 => 9325,
    3011 => 9328,
    3012 => 9331,
    3013 => 9334,
    3014 => 9337,
    3015 => 9340,
    3016 => 9343,
    3017 => 9346,
    3018 => 9349,
    3019 => 9352,
    3020 => 9355,
    3021 => 9358,
    3022 => 9361,
    3023 => 9364,
    3024 => 9367,
    3025 => 9370,
    3026 => 9373,
    3027 => 9376,
    3028 => 9379,
    3029 => 9382,
    3030 => 9385,
    3031 => 9388,
    3032 => 9391,
    3033 => 9394,
    3034 => 9397,
    3035 => 9400,
    3036 => 9403,
    3037 => 9406,
    3038 => 9409,
    3039 => 9413,
    3040 => 9416,
    3041 => 9419,
    3042 => 9422,
    3043 => 9425,
    3044 => 9428,
    3045 => 9431,
    3046 => 9434,
    3047 => 9437,
    3048 => 9440,
    3049 => 9443,
    3050 => 9446,
    3051 => 9449,
    3052 => 9452,
    3053 => 9455,
    3054 => 9458,
    3055 => 9461,
    3056 => 9464,
    3057 => 9467,
    3058 => 9470,
    3059 => 9473,
    3060 => 9476,
    3061 => 9479,
    3062 => 9482,
    3063 => 9485,
    3064 => 9488,
    3065 => 9491,
    3066 => 9494,
    3067 => 9497,
    3068 => 9500,
    3069 => 9503,
    3070 => 9506,
    3071 => 9509,
    3072 => 9512,
    3073 => 9515,
    3074 => 9518,
    3075 => 9521,
    3076 => 9524,
    3077 => 9527,
    3078 => 9530,
    3079 => 9533,
    3080 => 9536,
    3081 => 9539,
    3082 => 9542,
    3083 => 9545,
    3084 => 9548,
    3085 => 9551,
    3086 => 9554,
    3087 => 9557,
    3088 => 9560,
    3089 => 9563,
    3090 => 9566,
    3091 => 9569,
    3092 => 9572,
    3093 => 9575,
    3094 => 9578,
    3095 => 9581,
    3096 => 9584,
    3097 => 9587,
    3098 => 9590,
    3099 => 9593,
    3100 => 9596,
    3101 => 9599,
    3102 => 9602,
    3103 => 9605,
    3104 => 9608,
    3105 => 9611,
    3106 => 9614,
    3107 => 9617,
    3108 => 9620,
    3109 => 9623,
    3110 => 9626,
    3111 => 9629,
    3112 => 9632,
    3113 => 9635,
    3114 => 9638,
    3115 => 9641,
    3116 => 9644,
    3117 => 9647,
    3118 => 9650,
    3119 => 9653,
    3120 => 9656,
    3121 => 9659,
    3122 => 9662,
    3123 => 9665,
    3124 => 9668,
    3125 => 9671,
    3126 => 9674,
    3127 => 9677,
    3128 => 9680,
    3129 => 9683,
    3130 => 9686,
    3131 => 9689,
    3132 => 9692,
    3133 => 9695,
    3134 => 9698,
    3135 => 9701,
    3136 => 9704,
    3137 => 9707,
    3138 => 9710,
    3139 => 9713,
    3140 => 9716,
    3141 => 9719,
    3142 => 9722,
    3143 => 9725,
    3144 => 9728,
    3145 => 9731,
    3146 => 9734,
    3147 => 9737,
    3148 => 9740,
    3149 => 9743,
    3150 => 9746,
    3151 => 9749,
    3152 => 9752,
    3153 => 9755,
    3154 => 9758,
    3155 => 9761,
    3156 => 9764,
    3157 => 9767,
    3158 => 9770,
    3159 => 9773,
    3160 => 9776,
    3161 => 9779,
    3162 => 9782,
    3163 => 9785,
    3164 => 9788,
    3165 => 9791,
    3166 => 9794,
    3167 => 9797,
    3168 => 9800,
    3169 => 9803,
    3170 => 9806,
    3171 => 9809,
    3172 => 9812,
    3173 => 9815,
    3174 => 9818,
    3175 => 9821,
    3176 => 9824,
    3177 => 9827,
    3178 => 9830,
    3179 => 9833,
    3180 => 9836,
    3181 => 9839,
    3182 => 9842,
    3183 => 9845,
    3184 => 9848,
    3185 => 9851,
    3186 => 9854,
    3187 => 9857,
    3188 => 9860,
    3189 => 9863,
    3190 => 9866,
    3191 => 9869,
    3192 => 9872,
    3193 => 9875,
    3194 => 9878,
    3195 => 9881,
    3196 => 9884,
    3197 => 9887,
    3198 => 9890,
    3199 => 9893,
    3200 => 9896,
    3201 => 9899,
    3202 => 9902,
    3203 => 9905,
    3204 => 9908,
    3205 => 9911,
    3206 => 9914,
    3207 => 9917,
    3208 => 9920,
    3209 => 9923,
    3210 => 9926,
    3211 => 9929,
    3212 => 9932,
    3213 => 9935,
    3214 => 9938,
    3215 => 9941,
    3216 => 9944,
    3217 => 9947,
    3218 => 9950,
    3219 => 9953,
    3220 => 9956,
    3221 => 9959,
    3222 => 9962,
    3223 => 9965,
    3224 => 9968,
    3225 => 9971,
    3226 => 9974,
    3227 => 9977,
    3228 => 9980,
    3229 => 9983,
    3230 => 9986,
    3231 => 9989,
    3232 => 9992,
    3233 => 9995,
    3234 => 9998,
    3235 => 10001,
    3236 => 10004,
    3237 => 10007,
    3238 => 10010,
    3239 => 10013,
    3240 => 10016,
    3241 => 10019,
    3242 => 10022,
    3243 => 10025,
    3244 => 10028,
    3245 => 10031,
    3246 => 10033,
    3247 => 10036,
    3248 => 10039,
    3249 => 10042,
    3250 => 10045,
    3251 => 10048,
    3252 => 10051,
    3253 => 10054,
    3254 => 10057,
    3255 => 10060,
    3256 => 10063,
    3257 => 10066,
    3258 => 10069,
    3259 => 10072,
    3260 => 10075,
    3261 => 10078,
    3262 => 10081,
    3263 => 10084,
    3264 => 10087,
    3265 => 10090,
    3266 => 10093,
    3267 => 10096,
    3268 => 10099,
    3269 => 10102,
    3270 => 10105,
    3271 => 10108,
    3272 => 10111,
    3273 => 10114,
    3274 => 10117,
    3275 => 10120,
    3276 => 10123,
    3277 => 10126,
    3278 => 10129,
    3279 => 10132,
    3280 => 10135,
    3281 => 10138,
    3282 => 10141,
    3283 => 10144,
    3284 => 10147,
    3285 => 10150,
    3286 => 10153,
    3287 => 10156,
    3288 => 10159,
    3289 => 10162,
    3290 => 10165,
    3291 => 10168,
    3292 => 10171,
    3293 => 10174,
    3294 => 10177,
    3295 => 10180,
    3296 => 10183,
    3297 => 10186,
    3298 => 10189,
    3299 => 10192,
    3300 => 10195,
    3301 => 10198,
    3302 => 10201,
    3303 => 10204,
    3304 => 10207,
    3305 => 10210,
    3306 => 10213,
    3307 => 10216,
    3308 => 10219,
    3309 => 10222,
    3310 => 10225,
    3311 => 10228,
    3312 => 10231,
    3313 => 10234,
    3314 => 10237,
    3315 => 10240,
    3316 => 10243,
    3317 => 10246,
    3318 => 10249,
    3319 => 10252,
    3320 => 10255,
    3321 => 10258,
    3322 => 10261,
    3323 => 10263,
    3324 => 10266,
    3325 => 10269,
    3326 => 10272,
    3327 => 10275,
    3328 => 10278,
    3329 => 10281,
    3330 => 10284,
    3331 => 10287,
    3332 => 10290,
    3333 => 10293,
    3334 => 10296,
    3335 => 10299,
    3336 => 10302,
    3337 => 10305,
    3338 => 10308,
    3339 => 10311,
    3340 => 10314,
    3341 => 10317,
    3342 => 10320,
    3343 => 10323,
    3344 => 10326,
    3345 => 10329,
    3346 => 10332,
    3347 => 10335,
    3348 => 10338,
    3349 => 10341,
    3350 => 10344,
    3351 => 10347,
    3352 => 10350,
    3353 => 10353,
    3354 => 10356,
    3355 => 10359,
    3356 => 10362,
    3357 => 10365,
    3358 => 10368,
    3359 => 10371,
    3360 => 10374,
    3361 => 10377,
    3362 => 10380,
    3363 => 10383,
    3364 => 10386,
    3365 => 10389,
    3366 => 10392,
    3367 => 10395,
    3368 => 10398,
    3369 => 10401,
    3370 => 10404,
    3371 => 10407,
    3372 => 10410,
    3373 => 10413,
    3374 => 10416,
    3375 => 10419,
    3376 => 10421,
    3377 => 10424,
    3378 => 10427,
    3379 => 10430,
    3380 => 10433,
    3381 => 10436,
    3382 => 10439,
    3383 => 10442,
    3384 => 10445,
    3385 => 10448,
    3386 => 10451,
    3387 => 10454,
    3388 => 10457,
    3389 => 10460,
    3390 => 10463,
    3391 => 10466,
    3392 => 10469,
    3393 => 10472,
    3394 => 10475,
    3395 => 10478,
    3396 => 10481,
    3397 => 10484,
    3398 => 10487,
    3399 => 10490,
    3400 => 10493,
    3401 => 10496,
    3402 => 10499,
    3403 => 10502,
    3404 => 10505,
    3405 => 10508,
    3406 => 10511,
    3407 => 10514,
    3408 => 10517,
    3409 => 10520,
    3410 => 10523,
    3411 => 10526,
    3412 => 10529,
    3413 => 10532,
    3414 => 10535,
    3415 => 10538,
    3416 => 10541,
    3417 => 10544,
    3418 => 10546,
    3419 => 10549,
    3420 => 10552,
    3421 => 10555,
    3422 => 10558,
    3423 => 10561,
    3424 => 10564,
    3425 => 10567,
    3426 => 10570,
    3427 => 10573,
    3428 => 10576,
    3429 => 10579,
    3430 => 10582,
    3431 => 10585,
    3432 => 10588,
    3433 => 10591,
    3434 => 10594,
    3435 => 10597,
    3436 => 10600,
    3437 => 10603,
    3438 => 10606,
    3439 => 10609,
    3440 => 10612,
    3441 => 10615,
    3442 => 10618,
    3443 => 10621,
    3444 => 10624,
    3445 => 10627,
    3446 => 10630,
    3447 => 10633,
    3448 => 10636,
    3449 => 10639,
    3450 => 10642,
    3451 => 10645,
    3452 => 10648,
    3453 => 10651,
    3454 => 10654,
    3455 => 10656,
    3456 => 10659,
    3457 => 10662,
    3458 => 10665,
    3459 => 10668,
    3460 => 10671,
    3461 => 10674,
    3462 => 10677,
    3463 => 10680,
    3464 => 10683,
    3465 => 10686,
    3466 => 10689,
    3467 => 10692,
    3468 => 10695,
    3469 => 10698,
    3470 => 10701,
    3471 => 10704,
    3472 => 10707,
    3473 => 10710,
    3474 => 10713,
    3475 => 10716,
    3476 => 10719,
    3477 => 10722,
    3478 => 10725,
    3479 => 10728,
    3480 => 10731,
    3481 => 10734,
    3482 => 10737,
    3483 => 10740,
    3484 => 10743,
    3485 => 10746,
    3486 => 10749,
    3487 => 10751,
    3488 => 10754,
    3489 => 10757,
    3490 => 10760,
    3491 => 10763,
    3492 => 10766,
    3493 => 10769,
    3494 => 10772,
    3495 => 10775,
    3496 => 10778,
    3497 => 10781,
    3498 => 10784,
    3499 => 10787,
    3500 => 10790,
    3501 => 10793,
    3502 => 10796,
    3503 => 10799,
    3504 => 10802,
    3505 => 10805,
    3506 => 10808,
    3507 => 10811,
    3508 => 10814,
    3509 => 10817,
    3510 => 10820,
    3511 => 10823,
    3512 => 10826,
    3513 => 10829,
    3514 => 10832,
    3515 => 10835,
    3516 => 10838,
    3517 => 10840,
    3518 => 10843,
    3519 => 10846,
    3520 => 10849,
    3521 => 10852,
    3522 => 10855,
    3523 => 10858,
    3524 => 10861,
    3525 => 10864,
    3526 => 10867,
    3527 => 10870,
    3528 => 10873,
    3529 => 10876,
    3530 => 10879,
    3531 => 10882,
    3532 => 10885,
    3533 => 10888,
    3534 => 10891,
    3535 => 10894,
    3536 => 10897,
    3537 => 10900,
    3538 => 10903,
    3539 => 10906,
    3540 => 10909,
    3541 => 10912,
    3542 => 10915,
    3543 => 10918,
    3544 => 10920,
    3545 => 10923,
    3546 => 10926,
    3547 => 10929,
    3548 => 10932,
    3549 => 10935,
    3550 => 10938,
    3551 => 10941,
    3552 => 10944,
    3553 => 10947,
    3554 => 10950,
    3555 => 10953,
    3556 => 10956,
    3557 => 10959,
    3558 => 10962,
    3559 => 10965,
    3560 => 10968,
    3561 => 10971,
    3562 => 10974,
    3563 => 10977,
    3564 => 10980,
    3565 => 10983,
    3566 => 10986,
    3567 => 10989,
    3568 => 10992,
    3569 => 10994,
    3570 => 10997,
    3571 => 11000,
    3572 => 11003,
    3573 => 11006,
    3574 => 11009,
    3575 => 11012,
    3576 => 11015,
    3577 => 11018,
    3578 => 11021,
    3579 => 11024,
    3580 => 11027,
    3581 => 11030,
    3582 => 11033,
    3583 => 11036,
    3584 => 11039,
    3585 => 11042,
    3586 => 11045,
    3587 => 11048,
    3588 => 11051,
    3589 => 11054,
    3590 => 11057,
    3591 => 11060,
    3592 => 11063,
    3593 => 11065,
    3594 => 11068,
    3595 => 11071,
    3596 => 11074,
    3597 => 11077,
    3598 => 11080,
    3599 => 11083,
    3600 => 11086,
    3601 => 11089,
    3602 => 11092,
    3603 => 11095,
    3604 => 11098,
    3605 => 11101,
    3606 => 11104,
    3607 => 11107,
    3608 => 11110,
    3609 => 11113,
    3610 => 11116,
    3611 => 11119,
    3612 => 11122,
    3613 => 11125,
    3614 => 11128,
    3615 => 11131,
    3616 => 11133,
    3617 => 11136,
    3618 => 11139,
    3619 => 11142,
    3620 => 11145,
    3621 => 11148,
    3622 => 11151,
    3623 => 11154,
    3624 => 11157,
    3625 => 11160,
    3626 => 11163,
    3627 => 11166,
    3628 => 11169,
    3629 => 11172,
    3630 => 11175,
    3631 => 11178,
    3632 => 11181,
    3633 => 11184,
    3634 => 11187,
    3635 => 11190,
    3636 => 11193,
    3637 => 11195,
    3638 => 11198,
    3639 => 11201,
    3640 => 11204,
    3641 => 11207,
    3642 => 11210,
    3643 => 11213,
    3644 => 11216,
    3645 => 11219,
    3646 => 11222,
    3647 => 11225,
    3648 => 11228,
    3649 => 11231,
    3650 => 11234,
    3651 => 11237,
    3652 => 11240,
    3653 => 11243,
    3654 => 11246,
    3655 => 11249,
    3656 => 11252,
    3657 => 11255,
    3658 => 11257,
    3659 => 11260,
    3660 => 11263,
    3661 => 11266,
    3662 => 11269,
    3663 => 11272,
    3664 => 11275,
    3665 => 11278,
    3666 => 11281,
    3667 => 11284,
    3668 => 11287,
    3669 => 11290,
    3670 => 11293,
    3671 => 11296,
    3672 => 11299,
    3673 => 11302,
    3674 => 11305,
    3675 => 11308,
    3676 => 11311,
    3677 => 11314,
    3678 => 11316,
    3679 => 11319,
    3680 => 11322,
    3681 => 11325,
    3682 => 11328,
    3683 => 11331,
    3684 => 11334,
    3685 => 11337,
    3686 => 11340,
    3687 => 11343,
    3688 => 11346,
    3689 => 11349,
    3690 => 11352,
    3691 => 11355,
    3692 => 11358,
    3693 => 11361,
    3694 => 11364,
    3695 => 11367,
    3696 => 11370,
    3697 => 11372,
    3698 => 11375,
    3699 => 11378,
    3700 => 11381,
    3701 => 11384,
    3702 => 11387,
    3703 => 11390,
    3704 => 11393,
    3705 => 11396,
    3706 => 11399,
    3707 => 11402,
    3708 => 11405,
    3709 => 11408,
    3710 => 11411,
    3711 => 11414,
    3712 => 11417,
    3713 => 11420,
    3714 => 11423,
    3715 => 11425,
    3716 => 11428,
    3717 => 11431,
    3718 => 11434,
    3719 => 11437,
    3720 => 11440,
    3721 => 11443,
    3722 => 11446,
    3723 => 11449,
    3724 => 11452,
    3725 => 11455,
    3726 => 11458,
    3727 => 11461,
    3728 => 11464,
    3729 => 11467,
    3730 => 11470,
    3731 => 11473,
    3732 => 11476,
    3733 => 11478,
    3734 => 11481,
    3735 => 11484,
    3736 => 11487,
    3737 => 11490,
    3738 => 11493,
    3739 => 11496,
    3740 => 11499,
    3741 => 11502,
    3742 => 11505,
    3743 => 11508,
    3744 => 11511,
    3745 => 11514,
    3746 => 11517,
    3747 => 11520,
    3748 => 11523,
    3749 => 11526,
    3750 => 11528,
    3751 => 11531,
    3752 => 11534,
    3753 => 11537,
    3754 => 11540,
    3755 => 11543,
    3756 => 11546,
    3757 => 11549,
    3758 => 11552,
    3759 => 11555,
    3760 => 11558,
    3761 => 11561,
    3762 => 11564,
    3763 => 11567,
    3764 => 11570,
    3765 => 11573,
    3766 => 11575,
    3767 => 11578,
    3768 => 11581,
    3769 => 11584,
    3770 => 11587,
    3771 => 11590,
    3772 => 11593,
    3773 => 11596,
    3774 => 11599,
    3775 => 11602,
    3776 => 11605,
    3777 => 11608,
    3778 => 11611,
    3779 => 11614,
    3780 => 11617,
    3781 => 11620,
    3782 => 11623,
    3783 => 11625,
    3784 => 11628,
    3785 => 11631,
    3786 => 11634,
    3787 => 11637,
    3788 => 11640,
    3789 => 11643,
    3790 => 11646,
    3791 => 11649,
    3792 => 11652,
    3793 => 11655,
    3794 => 11658,
    3795 => 11661,
    3796 => 11664,
    3797 => 11667,
    3798 => 11669,
    3799 => 11672,
    3800 => 11675,
    3801 => 11678,
    3802 => 11681,
    3803 => 11684,
    3804 => 11687,
    3805 => 11690,
    3806 => 11693,
    3807 => 11696,
    3808 => 11699,
    3809 => 11702,
    3810 => 11705,
    3811 => 11708,
    3812 => 11711,
    3813 => 11714,
    3814 => 11716,
    3815 => 11719,
    3816 => 11722,
    3817 => 11725,
    3818 => 11728,
    3819 => 11731,
    3820 => 11734,
    3821 => 11737,
    3822 => 11740,
    3823 => 11743,
    3824 => 11746,
    3825 => 11749,
    3826 => 11752,
    3827 => 11755,
    3828 => 11758,
    3829 => 11760,
    3830 => 11763,
    3831 => 11766,
    3832 => 11769,
    3833 => 11772,
    3834 => 11775,
    3835 => 11778,
    3836 => 11781,
    3837 => 11784,
    3838 => 11787,
    3839 => 11790,
    3840 => 11793,
    3841 => 11796,
    3842 => 11799,
    3843 => 11801,
    3844 => 11804,
    3845 => 11807,
    3846 => 11810,
    3847 => 11813,
    3848 => 11816,
    3849 => 11819,
    3850 => 11822,
    3851 => 11825,
    3852 => 11828,
    3853 => 11831,
    3854 => 11834,
    3855 => 11837,
    3856 => 11840,
    3857 => 11842,
    3858 => 11845,
    3859 => 11848,
    3860 => 11851,
    3861 => 11854,
    3862 => 11857,
    3863 => 11860,
    3864 => 11863,
    3865 => 11866,
    3866 => 11869,
    3867 => 11872,
    3868 => 11875,
    3869 => 11878,
    3870 => 11881,
    3871 => 11883,
    3872 => 11886,
    3873 => 11889,
    3874 => 11892,
    3875 => 11895,
    3876 => 11898,
    3877 => 11901,
    3878 => 11904,
    3879 => 11907,
    3880 => 11910,
    3881 => 11913,
    3882 => 11916,
    3883 => 11919,
    3884 => 11922,
    3885 => 11924,
    3886 => 11927,
    3887 => 11930,
    3888 => 11933,
    3889 => 11936,
    3890 => 11939,
    3891 => 11942,
    3892 => 11945,
    3893 => 11948,
    3894 => 11951,
    3895 => 11954,
    3896 => 11957,
    3897 => 11960,
    3898 => 11962,
    3899 => 11965,
    3900 => 11968,
    3901 => 11971,
    3902 => 11974,
    3903 => 11977,
    3904 => 11980,
    3905 => 11983,
    3906 => 11986,
    3907 => 11989,
    3908 => 11992,
    3909 => 11995,
    3910 => 11998,
    3911 => 12001,
    3912 => 12003,
    3913 => 12006,
    3914 => 12009,
    3915 => 12012,
    3916 => 12015,
    3917 => 12018,
    3918 => 12021,
    3919 => 12024,
    3920 => 12027,
    3921 => 12030,
    3922 => 12033,
    3923 => 12036,
    3924 => 12038,
    3925 => 12041,
    3926 => 12044,
    3927 => 12047,
    3928 => 12050,
    3929 => 12053,
    3930 => 12056,
    3931 => 12059,
    3932 => 12062,
    3933 => 12065,
    3934 => 12068,
    3935 => 12071,
    3936 => 12074,
    3937 => 12076,
    3938 => 12079,
    3939 => 12082,
    3940 => 12085,
    3941 => 12088,
    3942 => 12091,
    3943 => 12094,
    3944 => 12097,
    3945 => 12100,
    3946 => 12103,
    3947 => 12106,
    3948 => 12109,
    3949 => 12112,
    3950 => 12114,
    3951 => 12117,
    3952 => 12120,
    3953 => 12123,
    3954 => 12126,
    3955 => 12129,
    3956 => 12132,
    3957 => 12135,
    3958 => 12138,
    3959 => 12141,
    3960 => 12144,
    3961 => 12147,
    3962 => 12149,
    3963 => 12152,
    3964 => 12155,
    3965 => 12158,
    3966 => 12161,
    3967 => 12164,
    3968 => 12167,
    3969 => 12170,
    3970 => 12173,
    3971 => 12176,
    3972 => 12179,
    3973 => 12182,
    3974 => 12184,
    3975 => 12187,
    3976 => 12190,
    3977 => 12193,
    3978 => 12196,
    3979 => 12199,
    3980 => 12202,
    3981 => 12205,
    3982 => 12208,
    3983 => 12211,
    3984 => 12214,
    3985 => 12217,
    3986 => 12219,
    3987 => 12222,
    3988 => 12225,
    3989 => 12228,
    3990 => 12231,
    3991 => 12234,
    3992 => 12237,
    3993 => 12240,
    3994 => 12243,
    3995 => 12246,
    3996 => 12249,
    3997 => 12251,
    3998 => 12254,
    3999 => 12257,
    4000 => 12260,
    4001 => 12263,
    4002 => 12266,
    4003 => 12269,
    4004 => 12272,
    4005 => 12275,
    4006 => 12278,
    4007 => 12281,
    4008 => 12284,
    4009 => 12286,
    4010 => 12289,
    4011 => 12292,
    4012 => 12295,
    4013 => 12298,
    4014 => 12301,
    4015 => 12304,
    4016 => 12307,
    4017 => 12310,
    4018 => 12313,
    4019 => 12316,
    4020 => 12318,
    4021 => 12321,
    4022 => 12324,
    4023 => 12327,
    4024 => 12330,
    4025 => 12333,
    4026 => 12336,
    4027 => 12339,
    4028 => 12342,
    4029 => 12345,
    4030 => 12348,
    4031 => 12350,
    4032 => 12353,
    4033 => 12356,
    4034 => 12359,
    4035 => 12362,
    4036 => 12365,
    4037 => 12368,
    4038 => 12371,
    4039 => 12374,
    4040 => 12377,
    4041 => 12380,
    4042 => 12382,
    4043 => 12385,
    4044 => 12388,
    4045 => 12391,
    4046 => 12394,
    4047 => 12397,
    4048 => 12400,
    4049 => 12403,
    4050 => 12406,
    4051 => 12409,
    4052 => 12412,
    4053 => 12414,
    4054 => 12417,
    4055 => 12420,
    4056 => 12423,
    4057 => 12426,
    4058 => 12429,
    4059 => 12432,
    4060 => 12435,
    4061 => 12438,
    4062 => 12441,
    4063 => 12444,
    4064 => 12446,
    4065 => 12449,
    4066 => 12452,
    4067 => 12455,
    4068 => 12458,
    4069 => 12461,
    4070 => 12464,
    4071 => 12467,
    4072 => 12470,
    4073 => 12473,
    4074 => 12476,
    4075 => 12478,
    4076 => 12481,
    4077 => 12484,
    4078 => 12487,
    4079 => 12490,
    4080 => 12493,
    4081 => 12496,
    4082 => 12499,
    4083 => 12502,
    4084 => 12505,
    4085 => 12507,
    4086 => 12510,
    4087 => 12513,
    4088 => 12516,
    4089 => 12519,
    4090 => 12522,
    4091 => 12525,
    4092 => 12528,
    4093 => 12531,
    4094 => 12534,
    4095 => 12536,
    4096 => 12539,
    4097 => 12542,
    4098 => 12545,
    4099 => 12548,
    4100 => 12551,
    4101 => 12554,
    4102 => 12557,
    4103 => 12560,
    4104 => 12563,
    4105 => 12566,
    4106 => 12568,
    4107 => 12571,
    4108 => 12574,
    4109 => 12577,
    4110 => 12580,
    4111 => 12583,
    4112 => 12586,
    4113 => 12589,
    4114 => 12592,
    4115 => 12595,
    4116 => 12597,
    4117 => 12600,
    4118 => 12603,
    4119 => 12606,
    4120 => 12609,
    4121 => 12612,
    4122 => 12615,
    4123 => 12618,
    4124 => 12621,
    4125 => 12624,
    4126 => 12626,
    4127 => 12629,
    4128 => 12632,
    4129 => 12635,
    4130 => 12638,
    4131 => 12641,
    4132 => 12644,
    4133 => 12647,
    4134 => 12650,
    4135 => 12652,
    4136 => 12655,
    4137 => 12658,
    4138 => 12661,
    4139 => 12664,
    4140 => 12667,
    4141 => 12670,
    4142 => 12673,
    4143 => 12676,
    4144 => 12679,
    4145 => 12681,
    4146 => 12684,
    4147 => 12687,
    4148 => 12690,
    4149 => 12693,
    4150 => 12696,
    4151 => 12699,
    4152 => 12702,
    4153 => 12705,
    4154 => 12708,
    4155 => 12710,
    4156 => 12713,
    4157 => 12716,
    4158 => 12719,
    4159 => 12722,
    4160 => 12725,
    4161 => 12728,
    4162 => 12731,
    4163 => 12734,
    4164 => 12736,
    4165 => 12739,
    4166 => 12742,
    4167 => 12745,
    4168 => 12748,
    4169 => 12751,
    4170 => 12754,
    4171 => 12757,
    4172 => 12760,
    4173 => 12763,
    4174 => 12765,
    4175 => 12768,
    4176 => 12771,
    4177 => 12774,
    4178 => 12777,
    4179 => 12780,
    4180 => 12783,
    4181 => 12786,
    4182 => 12789,
    4183 => 12791,
    4184 => 12794,
    4185 => 12797,
    4186 => 12800,
    4187 => 12803,
    4188 => 12806,
    4189 => 12809,
    4190 => 12812,
    4191 => 12815,
    4192 => 12817,
    4193 => 12820,
    4194 => 12823,
    4195 => 12826,
    4196 => 12829,
    4197 => 12832,
    4198 => 12835,
    4199 => 12838,
    4200 => 12841,
    4201 => 12843,
    4202 => 12846,
    4203 => 12849,
    4204 => 12852,
    4205 => 12855,
    4206 => 12858,
    4207 => 12861,
    4208 => 12864,
    4209 => 12867,
    4210 => 12870,
    4211 => 12872,
    4212 => 12875,
    4213 => 12878,
    4214 => 12881,
    4215 => 12884,
    4216 => 12887,
    4217 => 12890,
    4218 => 12893,
    4219 => 12895,
    4220 => 12898,
    4221 => 12901,
    4222 => 12904,
    4223 => 12907,
    4224 => 12910,
    4225 => 12913,
    4226 => 12916,
    4227 => 12919,
    4228 => 12921,
    4229 => 12924,
    4230 => 12927,
    4231 => 12930,
    4232 => 12933,
    4233 => 12936,
    4234 => 12939,
    4235 => 12942,
    4236 => 12945,
    4237 => 12947,
    4238 => 12950,
    4239 => 12953,
    4240 => 12956,
    4241 => 12959,
    4242 => 12962,
    4243 => 12965,
    4244 => 12968,
    4245 => 12971,
    4246 => 12973,
    4247 => 12976,
    4248 => 12979,
    4249 => 12982,
    4250 => 12985,
    4251 => 12988,
    4252 => 12991,
    4253 => 12994,
    4254 => 12997,
    4255 => 12999,
    4256 => 13002,
    4257 => 13005,
    4258 => 13008,
    4259 => 13011,
    4260 => 13014,
    4261 => 13017,
    4262 => 13020,
    4263 => 13022,
    4264 => 13025,
    4265 => 13028,
    4266 => 13031,
    4267 => 13034,
    4268 => 13037,
    4269 => 13040,
    4270 => 13043,
    4271 => 13046,
    4272 => 13048,
    4273 => 13051,
    4274 => 13054,
    4275 => 13057,
    4276 => 13060,
    4277 => 13063,
    4278 => 13066,
    4279 => 13069,
    4280 => 13071,
    4281 => 13074,
    4282 => 13077,
    4283 => 13080,
    4284 => 13083,
    4285 => 13086,
    4286 => 13089,
    4287 => 13092,
    4288 => 13094,
    4289 => 13097,
    4290 => 13100,
    4291 => 13103,
    4292 => 13106,
    4293 => 13109,
    4294 => 13112,
    4295 => 13115,
    4296 => 13118,
    4297 => 13120,
    4298 => 13123,
    4299 => 13126,
    4300 => 13129,
    4301 => 13132,
    4302 => 13135,
    4303 => 13138,
    4304 => 13141,
    4305 => 13143,
    4306 => 13146,
    4307 => 13149,
    4308 => 13152,
    4309 => 13155,
    4310 => 13158,
    4311 => 13161,
    4312 => 13164,
    4313 => 13166,
    4314 => 13169,
    4315 => 13172,
    4316 => 13175,
    4317 => 13178,
    4318 => 13181,
    4319 => 13184,
    4320 => 13187,
    4321 => 13189,
    4322 => 13192,
    4323 => 13195,
    4324 => 13198,
    4325 => 13201,
    4326 => 13204,
    4327 => 13207,
    4328 => 13210,
    4329 => 13212,
    4330 => 13215,
    4331 => 13218,
    4332 => 13221,
    4333 => 13224,
    4334 => 13227,
    4335 => 13230,
    4336 => 13233,
    4337 => 13235,
    4338 => 13238,
    4339 => 13241,
    4340 => 13244,
    4341 => 13247,
    4342 => 13250,
    4343 => 13253,
    4344 => 13256,
    4345 => 13258,
    4346 => 13261,
    4347 => 13264,
    4348 => 13267,
    4349 => 13270,
    4350 => 13273,
    4351 => 13276,
    4352 => 13279,
    4353 => 13281,
    4354 => 13284,
    4355 => 13287,
    4356 => 13290,
    4357 => 13293,
    4358 => 13296,
    4359 => 13299,
    4360 => 13302,
    4361 => 13304,
    4362 => 13307,
    4363 => 13310,
    4364 => 13313,
    4365 => 13316,
    4366 => 13319,
    4367 => 13322,
    4368 => 13324,
    4369 => 13327,
    4370 => 13330,
    4371 => 13333,
    4372 => 13336,
    4373 => 13339,
    4374 => 13342,
    4375 => 13345,
    4376 => 13347,
    4377 => 13350,
    4378 => 13353,
    4379 => 13356,
    4380 => 13359,
    4381 => 13362,
    4382 => 13365,
    4383 => 13368,
    4384 => 13370,
    4385 => 13373,
    4386 => 13376,
    4387 => 13379,
    4388 => 13382,
    4389 => 13385,
    4390 => 13388,
    4391 => 13390,
    4392 => 13393,
    4393 => 13396,
    4394 => 13399,
    4395 => 13402,
    4396 => 13405,
    4397 => 13408,
    4398 => 13411,
    4399 => 13413,
    4400 => 13416,
    4401 => 13419,
    4402 => 13422,
    4403 => 13425,
    4404 => 13428,
    4405 => 13431,
    4406 => 13433,
    4407 => 13436,
    4408 => 13439,
    4409 => 13442,
    4410 => 13445,
    4411 => 13448,
    4412 => 13451,
    4413 => 13454,
    4414 => 13456,
    4415 => 13459,
    4416 => 13462,
    4417 => 13465,
    4418 => 13468,
    4419 => 13471,
    4420 => 13474,
    4421 => 13476,
    4422 => 13479,
    4423 => 13482,
    4424 => 13485,
    4425 => 13488,
    4426 => 13491,
    4427 => 13494,
    4428 => 13496,
    4429 => 13499,
    4430 => 13502,
    4431 => 13505,
    4432 => 13508,
    4433 => 13511,
    4434 => 13514,
    4435 => 13516,
    4436 => 13519,
    4437 => 13522,
    4438 => 13525,
    4439 => 13528,
    4440 => 13531,
    4441 => 13534,
    4442 => 13537,
    4443 => 13539,
    4444 => 13542,
    4445 => 13545,
    4446 => 13548,
    4447 => 13551,
    4448 => 13554,
    4449 => 13557,
    4450 => 13559,
    4451 => 13562,
    4452 => 13565,
    4453 => 13568,
    4454 => 13571,
    4455 => 13574,
    4456 => 13577,
    4457 => 13579,
    4458 => 13582,
    4459 => 13585,
    4460 => 13588,
    4461 => 13591,
    4462 => 13594,
    4463 => 13597,
    4464 => 13599,
    4465 => 13602,
    4466 => 13605,
    4467 => 13608,
    4468 => 13611,
    4469 => 13614,
    4470 => 13617,
    4471 => 13619,
    4472 => 13622,
    4473 => 13625,
    4474 => 13628,
    4475 => 13631,
    4476 => 13634,
    4477 => 13637,
    4478 => 13639,
    4479 => 13642,
    4480 => 13645,
    4481 => 13648,
    4482 => 13651,
    4483 => 13654,
    4484 => 13657,
    4485 => 13659,
    4486 => 13662,
    4487 => 13665,
    4488 => 13668,
    4489 => 13671,
    4490 => 13674,
    4491 => 13677,
    4492 => 13679,
    4493 => 13682,
    4494 => 13685,
    4495 => 13688,
    4496 => 13691,
    4497 => 13694,
    4498 => 13697,
    4499 => 13699,
    4500 => 13702,
    4501 => 13705,
    4502 => 13708,
    4503 => 13711,
    4504 => 13714,
    4505 => 13717,
    4506 => 13719,
    4507 => 13722,
    4508 => 13725,
    4509 => 13728,
    4510 => 13731,
    4511 => 13734,
    4512 => 13736,
    4513 => 13739,
    4514 => 13742,
    4515 => 13745,
    4516 => 13748,
    4517 => 13751,
    4518 => 13754,
    4519 => 13756,
    4520 => 13759,
    4521 => 13762,
    4522 => 13765,
    4523 => 13768,
    4524 => 13771,
    4525 => 13774,
    4526 => 13776,
    4527 => 13779,
    4528 => 13782,
    4529 => 13785,
    4530 => 13788,
    4531 => 13791,
    4532 => 13793,
    4533 => 13796,
    4534 => 13799,
    4535 => 13802,
    4536 => 13805,
    4537 => 13808,
    4538 => 13811,
    4539 => 13813,
    4540 => 13816,
    4541 => 13819,
    4542 => 13822,
    4543 => 13825,
    4544 => 13828,
    4545 => 13831,
    4546 => 13833,
    4547 => 13836,
    4548 => 13839,
    4549 => 13842,
    4550 => 13845,
    4551 => 13848,
    4552 => 13850,
    4553 => 13853,
    4554 => 13856,
    4555 => 13859,
    4556 => 13862,
    4557 => 13865,
    4558 => 13868,
    4559 => 13870,
    4560 => 13873,
    4561 => 13876,
    4562 => 13879,
    4563 => 13882,
    4564 => 13885,
    4565 => 13887,
    4566 => 13890,
    4567 => 13893,
    4568 => 13896,
    4569 => 13899,
    4570 => 13902,
    4571 => 13905,
    4572 => 13907,
    4573 => 13910,
    4574 => 13913,
    4575 => 13916,
    4576 => 13919,
    4577 => 13922,
    4578 => 13924,
    4579 => 13927,
    4580 => 13930,
    4581 => 13933,
    4582 => 13936,
    4583 => 13939,
    4584 => 13942,
    4585 => 13944,
    4586 => 13947,
    4587 => 13950,
    4588 => 13953,
    4589 => 13956,
    4590 => 13959,
    4591 => 13961,
    4592 => 13964,
    4593 => 13967,
    4594 => 13970,
    4595 => 13973,
    4596 => 13976,
    4597 => 13978,
    4598 => 13981,
    4599 => 13984,
    4600 => 13987,
    4601 => 13990,
    4602 => 13993,
    4603 => 13995,
    4604 => 13998,
    4605 => 14001,
    4606 => 14004,
    4607 => 14007,
    4608 => 14010,
    4609 => 14013,
    4610 => 14015,
    4611 => 14018,
    4612 => 14021,
    4613 => 14024,
    4614 => 14027,
    4615 => 14030,
    4616 => 14032,
    4617 => 14035,
    4618 => 14038,
    4619 => 14041,
    4620 => 14044,
    4621 => 14047,
    4622 => 14049,
    4623 => 14052,
    4624 => 14055,
    4625 => 14058,
    4626 => 14061,
    4627 => 14064,
    4628 => 14066,
    4629 => 14069,
    4630 => 14072,
    4631 => 14075,
    4632 => 14078,
    4633 => 14081,
    4634 => 14083,
    4635 => 14086,
    4636 => 14089,
    4637 => 14092,
    4638 => 14095,
    4639 => 14098,
    4640 => 14101,
    4641 => 14103,
    4642 => 14106,
    4643 => 14109,
    4644 => 14112,
    4645 => 14115,
    4646 => 14118,
    4647 => 14120,
    4648 => 14123,
    4649 => 14126,
    4650 => 14129,
    4651 => 14132,
    4652 => 14135,
    4653 => 14137,
    4654 => 14140,
    4655 => 14143,
    4656 => 14146,
    4657 => 14149,
    4658 => 14152,
    4659 => 14154,
    4660 => 14157,
    4661 => 14160,
    4662 => 14163,
    4663 => 14166,
    4664 => 14169,
    4665 => 14171,
    4666 => 14174,
    4667 => 14177,
    4668 => 14180,
    4669 => 14183,
    4670 => 14186,
    4671 => 14188,
    4672 => 14191,
    4673 => 14194,
    4674 => 14197,
    4675 => 14200,
    4676 => 14203,
    4677 => 14205,
    4678 => 14208,
    4679 => 14211,
    4680 => 14214,
    4681 => 14217,
    4682 => 14219,
    4683 => 14222,
    4684 => 14225,
    4685 => 14228,
    4686 => 14231,
    4687 => 14234,
    4688 => 14236,
    4689 => 14239,
    4690 => 14242,
    4691 => 14245,
    4692 => 14248,
    4693 => 14251,
    4694 => 14253,
    4695 => 14256,
    4696 => 14259,
    4697 => 14262,
    4698 => 14265,
    4699 => 14268,
    4700 => 14270,
    4701 => 14273,
    4702 => 14276,
    4703 => 14279,
    4704 => 14282,
    4705 => 14285,
    4706 => 14287,
    4707 => 14290,
    4708 => 14293,
    4709 => 14296,
    4710 => 14299,
    4711 => 14302,
    4712 => 14304,
    4713 => 14307,
    4714 => 14310,
    4715 => 14313,
    4716 => 14316,
    4717 => 14318,
    4718 => 14321,
    4719 => 14324,
    4720 => 14327,
    4721 => 14330,
    4722 => 14333,
    4723 => 14335,
    4724 => 14338,
    4725 => 14341,
    4726 => 14344,
    4727 => 14347,
    4728 => 14350,
    4729 => 14352,
    4730 => 14355,
    4731 => 14358,
    4732 => 14361,
    4733 => 14364,
    4734 => 14366,
    4735 => 14369,
    4736 => 14372,
    4737 => 14375,
    4738 => 14378,
    4739 => 14381,
    4740 => 14383,
    4741 => 14386,
    4742 => 14389,
    4743 => 14392,
    4744 => 14395,
    4745 => 14398,
    4746 => 14400,
    4747 => 14403,
    4748 => 14406,
    4749 => 14409,
    4750 => 14412,
    4751 => 14414,
    4752 => 14417,
    4753 => 14420,
    4754 => 14423,
    4755 => 14426,
    4756 => 14429,
    4757 => 14431,
    4758 => 14434,
    4759 => 14437,
    4760 => 14440,
    4761 => 14443,
    4762 => 14445,
    4763 => 14448,
    4764 => 14451,
    4765 => 14454,
    4766 => 14457,
    4767 => 14460,
    4768 => 14462,
    4769 => 14465,
    4770 => 14468,
    4771 => 14471,
    4772 => 14474,
    4773 => 14477,
    4774 => 14479,
    4775 => 14482,
    4776 => 14485,
    4777 => 14488,
    4778 => 14491,
    4779 => 14493,
    4780 => 14496,
    4781 => 14499,
    4782 => 14502,
    4783 => 14505,
    4784 => 14507,
    4785 => 14510,
    4786 => 14513,
    4787 => 14516,
    4788 => 14519,
    4789 => 14522,
    4790 => 14524,
    4791 => 14527,
    4792 => 14530,
    4793 => 14533,
    4794 => 14536,
    4795 => 14538,
    4796 => 14541,
    4797 => 14544,
    4798 => 14547,
    4799 => 14550,
    4800 => 14553,
    4801 => 14555,
    4802 => 14558,
    4803 => 14561,
    4804 => 14564,
    4805 => 14567,
    4806 => 14569,
    4807 => 14572,
    4808 => 14575,
    4809 => 14578,
    4810 => 14581,
    4811 => 14584,
    4812 => 14586,
    4813 => 14589,
    4814 => 14592,
    4815 => 14595,
    4816 => 14598,
    4817 => 14600,
    4818 => 14603,
    4819 => 14606,
    4820 => 14609,
    4821 => 14612,
    4822 => 14614,
    4823 => 14617,
    4824 => 14620,
    4825 => 14623,
    4826 => 14626,
    4827 => 14628,
    4828 => 14631,
    4829 => 14634,
    4830 => 14637,
    4831 => 14640,
    4832 => 14643,
    4833 => 14645,
    4834 => 14648,
    4835 => 14651,
    4836 => 14654,
    4837 => 14657,
    4838 => 14659,
    4839 => 14662,
    4840 => 14665,
    4841 => 14668,
    4842 => 14671,
    4843 => 14673,
    4844 => 14676,
    4845 => 14679,
    4846 => 14682,
    4847 => 14685,
    4848 => 14688,
    4849 => 14690,
    4850 => 14693,
    4851 => 14696,
    4852 => 14699,
    4853 => 14702,
    4854 => 14704,
    4855 => 14707,
    4856 => 14710,
    4857 => 14713,
    4858 => 14716,
    4859 => 14718,
    4860 => 14721,
    4861 => 14724,
    4862 => 14727,
    4863 => 14730,
    4864 => 14732,
    4865 => 14735,
    4866 => 14738,
    4867 => 14741,
    4868 => 14744,
    4869 => 14746,
    4870 => 14749,
    4871 => 14752,
    4872 => 14755,
    4873 => 14758,
    4874 => 14760,
    4875 => 14763,
    4876 => 14766,
    4877 => 14769,
    4878 => 14772,
    4879 => 14774,
    4880 => 14777,
    4881 => 14780,
    4882 => 14783,
    4883 => 14786,
    4884 => 14789,
    4885 => 14791,
    4886 => 14794,
    4887 => 14797,
    4888 => 14800,
    4889 => 14803,
    4890 => 14805,
    4891 => 14808,
    4892 => 14811,
    4893 => 14814,
    4894 => 14817,
    4895 => 14819,
    4896 => 14822,
    4897 => 14825,
    4898 => 14828,
    4899 => 14831,
    4900 => 14833,
    4901 => 14836,
    4902 => 14839,
    4903 => 14842,
    4904 => 14845,
    4905 => 14847,
    4906 => 14850,
    4907 => 14853,
    4908 => 14856,
    4909 => 14859,
    4910 => 14861,
    4911 => 14864,
    4912 => 14867,
    4913 => 14870,
    4914 => 14873,
    4915 => 14875,
    4916 => 14878,
    4917 => 14881,
    4918 => 14884,
    4919 => 14887,
    4920 => 14889,
    4921 => 14892,
    4922 => 14895,
    4923 => 14898,
    4924 => 14901,
    4925 => 14903,
    4926 => 14906,
    4927 => 14909,
    4928 => 14912,
    4929 => 14915,
    4930 => 14917,
    4931 => 14920,
    4932 => 14923,
    4933 => 14926,
    4934 => 14929,
    4935 => 14931,
    4936 => 14934,
    4937 => 14937,
    4938 => 14940,
    4939 => 14942,
    4940 => 14945,
    4941 => 14948,
    4942 => 14951,
    4943 => 14954,
    4944 => 14956,
    4945 => 14959,
    4946 => 14962,
    4947 => 14965,
    4948 => 14968,
    4949 => 14970,
    4950 => 14973,
    4951 => 14976,
    4952 => 14979,
    4953 => 14982,
    4954 => 14984,
    4955 => 14987,
    4956 => 14990,
    4957 => 14993,
    4958 => 14996,
    4959 => 14998,
    4960 => 15001,
    4961 => 15004,
    4962 => 15007,
    4963 => 15010,
    4964 => 15012,
    4965 => 15015,
    4966 => 15018,
    4967 => 15021,
    4968 => 15024,
    4969 => 15026,
    4970 => 15029,
    4971 => 15032,
    4972 => 15035,
    4973 => 15037,
    4974 => 15040,
    4975 => 15043,
    4976 => 15046,
    4977 => 15049,
    4978 => 15051,
    4979 => 15054,
    4980 => 15057,
    4981 => 15060,
    4982 => 15063,
    4983 => 15065,
    4984 => 15068,
    4985 => 15071,
    4986 => 15074,
    4987 => 15077,
    4988 => 15079,
    4989 => 15082,
    4990 => 15085,
    4991 => 15088,
    4992 => 15090,
    4993 => 15093,
    4994 => 15096,
    4995 => 15099,
    4996 => 15102,
    4997 => 15104,
    4998 => 15107,
    4999 => 15110,
    5000 => 15113,
    5001 => 15116,
    5002 => 15118,
    5003 => 15121,
    5004 => 15124,
    5005 => 15127,
    5006 => 15129,
    5007 => 15132,
    5008 => 15135,
    5009 => 15138,
    5010 => 15141,
    5011 => 15143,
    5012 => 15146,
    5013 => 15149,
    5014 => 15152,
    5015 => 15155,
    5016 => 15157,
    5017 => 15160,
    5018 => 15163,
    5019 => 15166,
    5020 => 15168,
    5021 => 15171,
    5022 => 15174,
    5023 => 15177,
    5024 => 15180,
    5025 => 15182,
    5026 => 15185,
    5027 => 15188,
    5028 => 15191,
    5029 => 15194,
    5030 => 15196,
    5031 => 15199,
    5032 => 15202,
    5033 => 15205,
    5034 => 15207,
    5035 => 15210,
    5036 => 15213,
    5037 => 15216,
    5038 => 15219,
    5039 => 15221,
    5040 => 15224,
    5041 => 15227,
    5042 => 15230,
    5043 => 15233,
    5044 => 15235,
    5045 => 15238,
    5046 => 15241,
    5047 => 15244,
    5048 => 15246,
    5049 => 15249,
    5050 => 15252,
    5051 => 15255,
    5052 => 15258,
    5053 => 15260,
    5054 => 15263,
    5055 => 15266,
    5056 => 15269,
    5057 => 15271,
    5058 => 15274,
    5059 => 15277,
    5060 => 15280,
    5061 => 15283,
    5062 => 15285,
    5063 => 15288,
    5064 => 15291,
    5065 => 15294,
    5066 => 15296,
    5067 => 15299,
    5068 => 15302,
    5069 => 15305,
    5070 => 15308,
    5071 => 15310,
    5072 => 15313,
    5073 => 15316,
    5074 => 15319,
    5075 => 15321,
    5076 => 15324,
    5077 => 15327,
    5078 => 15330,
    5079 => 15333,
    5080 => 15335,
    5081 => 15338,
    5082 => 15341,
    5083 => 15344,
    5084 => 15346,
    5085 => 15349,
    5086 => 15352,
    5087 => 15355,
    5088 => 15358,
    5089 => 15360,
    5090 => 15363,
    5091 => 15366,
    5092 => 15369,
    5093 => 15371,
    5094 => 15374,
    5095 => 15377,
    5096 => 15380,
    5097 => 15382,
    5098 => 15385,
    5099 => 15388,
    5100 => 15391,
    5101 => 15394,
    5102 => 15396,
    5103 => 15399,
    5104 => 15402,
    5105 => 15405,
    5106 => 15407,
    5107 => 15410,
    5108 => 15413,
    5109 => 15416,
    5110 => 15419,
    5111 => 15421,
    5112 => 15424,
    5113 => 15427,
    5114 => 15430,
    5115 => 15432,
    5116 => 15435,
    5117 => 15438,
    5118 => 15441,
    5119 => 15443,
    5120 => 15446,
    5121 => 15449,
    5122 => 15452,
    5123 => 15455,
    5124 => 15457,
    5125 => 15460,
    5126 => 15463,
    5127 => 15466,
    5128 => 15468,
    5129 => 15471,
    5130 => 15474,
    5131 => 15477,
    5132 => 15479,
    5133 => 15482,
    5134 => 15485,
    5135 => 15488,
    5136 => 15491,
    5137 => 15493,
    5138 => 15496,
    5139 => 15499,
    5140 => 15502,
    5141 => 15504,
    5142 => 15507,
    5143 => 15510,
    5144 => 15513,
    5145 => 15515,
    5146 => 15518,
    5147 => 15521,
    5148 => 15524,
    5149 => 15527,
    5150 => 15529,
    5151 => 15532,
    5152 => 15535,
    5153 => 15538,
    5154 => 15540,
    5155 => 15543,
    5156 => 15546,
    5157 => 15549,
    5158 => 15551,
    5159 => 15554,
    5160 => 15557,
    5161 => 15560,
    5162 => 15562,
    5163 => 15565,
    5164 => 15568,
    5165 => 15571,
    5166 => 15574,
    5167 => 15576,
    5168 => 15579,
    5169 => 15582,
    5170 => 15585,
    5171 => 15587,
    5172 => 15590,
    5173 => 15593,
    5174 => 15596,
    5175 => 15598,
    5176 => 15601,
    5177 => 15604,
    5178 => 15607,
    5179 => 15609,
    5180 => 15612,
    5181 => 15615,
    5182 => 15618,
    5183 => 15621,
    5184 => 15623,
    5185 => 15626,
    5186 => 15629,
    5187 => 15632,
    5188 => 15634,
    5189 => 15637,
    5190 => 15640,
    5191 => 15643,
    5192 => 15645,
    5193 => 15648,
    5194 => 15651,
    5195 => 15654,
    5196 => 15656,
    5197 => 15659,
    5198 => 15662,
    5199 => 15665,
    5200 => 15667,
    5201 => 15670,
    5202 => 15673,
    5203 => 15676,
    5204 => 15678,
    5205 => 15681,
    5206 => 15684,
    5207 => 15687,
    5208 => 15690,
    5209 => 15692,
    5210 => 15695,
    5211 => 15698,
    5212 => 15701,
    5213 => 15703,
    5214 => 15706,
    5215 => 15709,
    5216 => 15712,
    5217 => 15714,
    5218 => 15717,
    5219 => 15720,
    5220 => 15723,
    5221 => 15725,
    5222 => 15728,
    5223 => 15731,
    5224 => 15734,
    5225 => 15736,
    5226 => 15739,
    5227 => 15742,
    5228 => 15745,
    5229 => 15747,
    5230 => 15750,
    5231 => 15753,
    5232 => 15756,
    5233 => 15758,
    5234 => 15761,
    5235 => 15764,
    5236 => 15767,
    5237 => 15769,
    5238 => 15772,
    5239 => 15775,
    5240 => 15778,
    5241 => 15780,
    5242 => 15783,
    5243 => 15786,
    5244 => 15789,
    5245 => 15791,
    5246 => 15794,
    5247 => 15797,
    5248 => 15800,
    5249 => 15802,
    5250 => 15805,
    5251 => 15808,
    5252 => 15811,
    5253 => 15813,
    5254 => 15816,
    5255 => 15819,
    5256 => 15822,
    5257 => 15824,
    5258 => 15827,
    5259 => 15830,
    5260 => 15833,
    5261 => 15835,
    5262 => 15838,
    5263 => 15841,
    5264 => 15844,
    5265 => 15846,
    5266 => 15849,
    5267 => 15852,
    5268 => 15855,
    5269 => 15857,
    5270 => 15860,
    5271 => 15863,
    5272 => 15866,
    5273 => 15868,
    5274 => 15871,
    5275 => 15874,
    5276 => 15877,
    5277 => 15879,
    5278 => 15882,
    5279 => 15885,
    5280 => 15888,
    5281 => 15890,
    5282 => 15893,
    5283 => 15896,
    5284 => 15899,
    5285 => 15901,
    5286 => 15904,
    5287 => 15907,
    5288 => 15910,
    5289 => 15912,
    5290 => 15915,
    5291 => 15918,
    5292 => 15921,
    5293 => 15923,
    5294 => 15926,
    5295 => 15929,
    5296 => 15932,
    5297 => 15934,
    5298 => 15937,
    5299 => 15940,
    5300 => 15943,
    5301 => 15945,
    5302 => 15948,
    5303 => 15951,
    5304 => 15954,
    5305 => 15956,
    5306 => 15959,
    5307 => 15962,
    5308 => 15965,
    5309 => 15967,
    5310 => 15970,
    5311 => 15973,
    5312 => 15976,
    5313 => 15978,
    5314 => 15981,
    5315 => 15984,
    5316 => 15987,
    5317 => 15989,
    5318 => 15992,
    5319 => 15995,
    5320 => 15997,
    5321 => 16000,
    5322 => 16003,
    5323 => 16006,
    5324 => 16008,
    5325 => 16011,
    5326 => 16014,
    5327 => 16017,
    5328 => 16019,
    5329 => 16022,
    5330 => 16025,
    5331 => 16028,
    5332 => 16030,
    5333 => 16033,
    5334 => 16036,
    5335 => 16039,
    5336 => 16041,
    5337 => 16044,
    5338 => 16047,
    5339 => 16050,
    5340 => 16052,
    5341 => 16055,
    5342 => 16058,
    5343 => 16061,
    5344 => 16063,
    5345 => 16066,
    5346 => 16069,
    5347 => 16071,
    5348 => 16074,
    5349 => 16077,
    5350 => 16080,
    5351 => 16082,
    5352 => 16085,
    5353 => 16088,
    5354 => 16091,
    5355 => 16093,
    5356 => 16096,
    5357 => 16099,
    5358 => 16102,
    5359 => 16104,
    5360 => 16107,
    5361 => 16110,
    5362 => 16113,
    5363 => 16115,
    5364 => 16118,
    5365 => 16121,
    5366 => 16123,
    5367 => 16126,
    5368 => 16129,
    5369 => 16132,
    5370 => 16134,
    5371 => 16137,
    5372 => 16140,
    5373 => 16143,
    5374 => 16145,
    5375 => 16148,
    5376 => 16151,
    5377 => 16154,
    5378 => 16156,
    5379 => 16159,
    5380 => 16162,
    5381 => 16164,
    5382 => 16167,
    5383 => 16170,
    5384 => 16173,
    5385 => 16175,
    5386 => 16178,
    5387 => 16181,
    5388 => 16184,
    5389 => 16186,
    5390 => 16189,
    5391 => 16192,
    5392 => 16195,
    5393 => 16197,
    5394 => 16200,
    5395 => 16203,
    5396 => 16205,
    5397 => 16208,
    5398 => 16211,
    5399 => 16214,
    5400 => 16216,
    5401 => 16219,
    5402 => 16222,
    5403 => 16225,
    5404 => 16227,
    5405 => 16230,
    5406 => 16233,
    5407 => 16235,
    5408 => 16238,
    5409 => 16241,
    5410 => 16244,
    5411 => 16246,
    5412 => 16249,
    5413 => 16252,
    5414 => 16255,
    5415 => 16257,
    5416 => 16260,
    5417 => 16263,
    5418 => 16265,
    5419 => 16268,
    5420 => 16271,
    5421 => 16274,
    5422 => 16276,
    5423 => 16279,
    5424 => 16282,
    5425 => 16285,
    5426 => 16287,
    5427 => 16290,
    5428 => 16293,
    5429 => 16295,
    5430 => 16298,
    5431 => 16301,
    5432 => 16304,
    5433 => 16306,
    5434 => 16309,
    5435 => 16312,
    5436 => 16315,
    5437 => 16317,
    5438 => 16320,
    5439 => 16323,
    5440 => 16325,
    5441 => 16328,
    5442 => 16331,
    5443 => 16334,
    5444 => 16336,
    5445 => 16339,
    5446 => 16342,
    5447 => 16344,
    5448 => 16347,
    5449 => 16350,
    5450 => 16353,
    5451 => 16355,
    5452 => 16358,
    5453 => 16361,
    5454 => 16364,
    5455 => 16366,
    5456 => 16369,
    5457 => 16372,
    5458 => 16374,
    5459 => 16377,
    5460 => 16380,
    5461 => 16383,
    5462 => 16385,
    5463 => 16388,
    5464 => 16391,
    5465 => 16393,
    5466 => 16396,
    5467 => 16399,
    5468 => 16402,
    5469 => 16404,
    5470 => 16407,
    5471 => 16410,
    5472 => 16413,
    5473 => 16415,
    5474 => 16418,
    5475 => 16421,
    5476 => 16423,
    5477 => 16426,
    5478 => 16429,
    5479 => 16432,
    5480 => 16434,
    5481 => 16437,
    5482 => 16440,
    5483 => 16442,
    5484 => 16445,
    5485 => 16448,
    5486 => 16451,
    5487 => 16453,
    5488 => 16456,
    5489 => 16459,
    5490 => 16461,
    5491 => 16464,
    5492 => 16467,
    5493 => 16470,
    5494 => 16472,
    5495 => 16475,
    5496 => 16478,
    5497 => 16480,
    5498 => 16483,
    5499 => 16486,
    5500 => 16489,
    5501 => 16491,
    5502 => 16494,
    5503 => 16497,
    5504 => 16499,
    5505 => 16502,
    5506 => 16505,
    5507 => 16508,
    5508 => 16510,
    5509 => 16513,
    5510 => 16516,
    5511 => 16518,
    5512 => 16521,
    5513 => 16524,
    5514 => 16527,
    5515 => 16529,
    5516 => 16532,
    5517 => 16535,
    5518 => 16537,
    5519 => 16540,
    5520 => 16543,
    5521 => 16546,
    5522 => 16548,
    5523 => 16551,
    5524 => 16554,
    5525 => 16556,
    5526 => 16559,
    5527 => 16562,
    5528 => 16565,
    5529 => 16567,
    5530 => 16570,
    5531 => 16573,
    5532 => 16575,
    5533 => 16578,
    5534 => 16581,
    5535 => 16584,
    5536 => 16586,
    5537 => 16589,
    5538 => 16592,
    5539 => 16594,
    5540 => 16597,
    5541 => 16600,
    5542 => 16602,
    5543 => 16605,
    5544 => 16608,
    5545 => 16611,
    5546 => 16613,
    5547 => 16616,
    5548 => 16619,
    5549 => 16621,
    5550 => 16624,
    5551 => 16627,
    5552 => 16630,
    5553 => 16632,
    5554 => 16635,
    5555 => 16638,
    5556 => 16640,
    5557 => 16643,
    5558 => 16646,
    5559 => 16648,
    5560 => 16651,
    5561 => 16654,
    5562 => 16657,
    5563 => 16659,
    5564 => 16662,
    5565 => 16665,
    5566 => 16667,
    5567 => 16670,
    5568 => 16673,
    5569 => 16676,
    5570 => 16678,
    5571 => 16681,
    5572 => 16684,
    5573 => 16686,
    5574 => 16689,
    5575 => 16692,
    5576 => 16694,
    5577 => 16697,
    5578 => 16700,
    5579 => 16703,
    5580 => 16705,
    5581 => 16708,
    5582 => 16711,
    5583 => 16713,
    5584 => 16716,
    5585 => 16719,
    5586 => 16721,
    5587 => 16724,
    5588 => 16727,
    5589 => 16730,
    5590 => 16732,
    5591 => 16735,
    5592 => 16738,
    5593 => 16740,
    5594 => 16743,
    5595 => 16746,
    5596 => 16749,
    5597 => 16751,
    5598 => 16754,
    5599 => 16757,
    5600 => 16759,
    5601 => 16762,
    5602 => 16765,
    5603 => 16767,
    5604 => 16770,
    5605 => 16773,
    5606 => 16775,
    5607 => 16778,
    5608 => 16781,
    5609 => 16784,
    5610 => 16786,
    5611 => 16789,
    5612 => 16792,
    5613 => 16794,
    5614 => 16797,
    5615 => 16800,
    5616 => 16802,
    5617 => 16805,
    5618 => 16808,
    5619 => 16811,
    5620 => 16813,
    5621 => 16816,
    5622 => 16819,
    5623 => 16821,
    5624 => 16824,
    5625 => 16827,
    5626 => 16829,
    5627 => 16832,
    5628 => 16835,
    5629 => 16838,
    5630 => 16840,
    5631 => 16843,
    5632 => 16846,
    5633 => 16848,
    5634 => 16851,
    5635 => 16854,
    5636 => 16856,
    5637 => 16859,
    5638 => 16862,
    5639 => 16864,
    5640 => 16867,
    5641 => 16870,
    5642 => 16873,
    5643 => 16875,
    5644 => 16878,
    5645 => 16881,
    5646 => 16883,
    5647 => 16886,
    5648 => 16889,
    5649 => 16891,
    5650 => 16894,
    5651 => 16897,
    5652 => 16899,
    5653 => 16902,
    5654 => 16905,
    5655 => 16908,
    5656 => 16910,
    5657 => 16913,
    5658 => 16916,
    5659 => 16918,
    5660 => 16921,
    5661 => 16924,
    5662 => 16926,
    5663 => 16929,
    5664 => 16932,
    5665 => 16934,
    5666 => 16937,
    5667 => 16940,
    5668 => 16943,
    5669 => 16945,
    5670 => 16948,
    5671 => 16951,
    5672 => 16953,
    5673 => 16956,
    5674 => 16959,
    5675 => 16961,
    5676 => 16964,
    5677 => 16967,
    5678 => 16969,
    5679 => 16972,
    5680 => 16975,
    5681 => 16977,
    5682 => 16980,
    5683 => 16983,
    5684 => 16986,
    5685 => 16988,
    5686 => 16991,
    5687 => 16994,
    5688 => 16996,
    5689 => 16999,
    5690 => 17002,
    5691 => 17004,
    5692 => 17007,
    5693 => 17010,
    5694 => 17012,
    5695 => 17015,
    5696 => 17018,
    5697 => 17020,
    5698 => 17023,
    5699 => 17026,
    5700 => 17028,
    5701 => 17031,
    5702 => 17034,
    5703 => 17037,
    5704 => 17039,
    5705 => 17042,
    5706 => 17045,
    5707 => 17047,
    5708 => 17050,
    5709 => 17053,
    5710 => 17055,
    5711 => 17058,
    5712 => 17061,
    5713 => 17063,
    5714 => 17066,
    5715 => 17069,
    5716 => 17071,
    5717 => 17074,
    5718 => 17077,
    5719 => 17079,
    5720 => 17082,
    5721 => 17085,
    5722 => 17087,
    5723 => 17090,
    5724 => 17093,
    5725 => 17096,
    5726 => 17098,
    5727 => 17101,
    5728 => 17104,
    5729 => 17106,
    5730 => 17109,
    5731 => 17112,
    5732 => 17114,
    5733 => 17117,
    5734 => 17120,
    5735 => 17122,
    5736 => 17125,
    5737 => 17128,
    5738 => 17130,
    5739 => 17133,
    5740 => 17136,
    5741 => 17138,
    5742 => 17141,
    5743 => 17144,
    5744 => 17146,
    5745 => 17149,
    5746 => 17152,
    5747 => 17154,
    5748 => 17157,
    5749 => 17160,
    5750 => 17162,
    5751 => 17165,
    5752 => 17168,
    5753 => 17171,
    5754 => 17173,
    5755 => 17176,
    5756 => 17179,
    5757 => 17181,
    5758 => 17184,
    5759 => 17187,
    5760 => 17189,
    5761 => 17192,
    5762 => 17195,
    5763 => 17197,
    5764 => 17200,
    5765 => 17203,
    5766 => 17205,
    5767 => 17208,
    5768 => 17211,
    5769 => 17213,
    5770 => 17216,
    5771 => 17219,
    5772 => 17221,
    5773 => 17224,
    5774 => 17227,
    5775 => 17229,
    5776 => 17232,
    5777 => 17235,
    5778 => 17237,
    5779 => 17240,
    5780 => 17243,
    5781 => 17245,
    5782 => 17248,
    5783 => 17251,
    5784 => 17253,
    5785 => 17256,
    5786 => 17259,
    5787 => 17261,
    5788 => 17264,
    5789 => 17267,
    5790 => 17269,
    5791 => 17272,
    5792 => 17275,
    5793 => 17277,
    5794 => 17280,
    5795 => 17283,
    5796 => 17285,
    5797 => 17288,
    5798 => 17291,
    5799 => 17293,
    5800 => 17296,
    5801 => 17299,
    5802 => 17301,
    5803 => 17304,
    5804 => 17307,
    5805 => 17309,
    5806 => 17312,
    5807 => 17315,
    5808 => 17317,
    5809 => 17320,
    5810 => 17323,
    5811 => 17325,
    5812 => 17328,
    5813 => 17331,
    5814 => 17333,
    5815 => 17336,
    5816 => 17339,
    5817 => 17341,
    5818 => 17344,
    5819 => 17347,
    5820 => 17349,
    5821 => 17352,
    5822 => 17355,
    5823 => 17357,
    5824 => 17360,
    5825 => 17363,
    5826 => 17365,
    5827 => 17368,
    5828 => 17371,
    5829 => 17373,
    5830 => 17376,
    5831 => 17379,
    5832 => 17381,
    5833 => 17384,
    5834 => 17387,
    5835 => 17389,
    5836 => 17392,
    5837 => 17395,
    5838 => 17397,
    5839 => 17400,
    5840 => 17403,
    5841 => 17405,
    5842 => 17408,
    5843 => 17411,
    5844 => 17413,
    5845 => 17416,
    5846 => 17419,
    5847 => 17421,
    5848 => 17424,
    5849 => 17427,
    5850 => 17429,
    5851 => 17432,
    5852 => 17435,
    5853 => 17437,
    5854 => 17440,
    5855 => 17443,
    5856 => 17445,
    5857 => 17448,
    5858 => 17451,
    5859 => 17453,
    5860 => 17456,
    5861 => 17459,
    5862 => 17461,
    5863 => 17464,
    5864 => 17467,
    5865 => 17469,
    5866 => 17472,
    5867 => 17474,
    5868 => 17477,
    5869 => 17480,
    5870 => 17482,
    5871 => 17485,
    5872 => 17488,
    5873 => 17490,
    5874 => 17493,
    5875 => 17496,
    5876 => 17498,
    5877 => 17501,
    5878 => 17504,
    5879 => 17506,
    5880 => 17509,
    5881 => 17512,
    5882 => 17514,
    5883 => 17517,
    5884 => 17520,
    5885 => 17522,
    5886 => 17525,
    5887 => 17528,
    5888 => 17530,
    5889 => 17533,
    5890 => 17536,
    5891 => 17538,
    5892 => 17541,
    5893 => 17544,
    5894 => 17546,
    5895 => 17549,
    5896 => 17551,
    5897 => 17554,
    5898 => 17557,
    5899 => 17559,
    5900 => 17562,
    5901 => 17565,
    5902 => 17567,
    5903 => 17570,
    5904 => 17573,
    5905 => 17575,
    5906 => 17578,
    5907 => 17581,
    5908 => 17583,
    5909 => 17586,
    5910 => 17589,
    5911 => 17591,
    5912 => 17594,
    5913 => 17597,
    5914 => 17599,
    5915 => 17602,
    5916 => 17605,
    5917 => 17607,
    5918 => 17610,
    5919 => 17612,
    5920 => 17615,
    5921 => 17618,
    5922 => 17620,
    5923 => 17623,
    5924 => 17626,
    5925 => 17628,
    5926 => 17631,
    5927 => 17634,
    5928 => 17636,
    5929 => 17639,
    5930 => 17642,
    5931 => 17644,
    5932 => 17647,
    5933 => 17650,
    5934 => 17652,
    5935 => 17655,
    5936 => 17657,
    5937 => 17660,
    5938 => 17663,
    5939 => 17665,
    5940 => 17668,
    5941 => 17671,
    5942 => 17673,
    5943 => 17676,
    5944 => 17679,
    5945 => 17681,
    5946 => 17684,
    5947 => 17687,
    5948 => 17689,
    5949 => 17692,
    5950 => 17695,
    5951 => 17697,
    5952 => 17700,
    5953 => 17702,
    5954 => 17705,
    5955 => 17708,
    5956 => 17710,
    5957 => 17713,
    5958 => 17716,
    5959 => 17718,
    5960 => 17721,
    5961 => 17724,
    5962 => 17726,
    5963 => 17729,
    5964 => 17732,
    5965 => 17734,
    5966 => 17737,
    5967 => 17739,
    5968 => 17742,
    5969 => 17745,
    5970 => 17747,
    5971 => 17750,
    5972 => 17753,
    5973 => 17755,
    5974 => 17758,
    5975 => 17761,
    5976 => 17763,
    5977 => 17766,
    5978 => 17768,
    5979 => 17771,
    5980 => 17774,
    5981 => 17776,
    5982 => 17779,
    5983 => 17782,
    5984 => 17784,
    5985 => 17787,
    5986 => 17790,
    5987 => 17792,
    5988 => 17795,
    5989 => 17798,
    5990 => 17800,
    5991 => 17803,
    5992 => 17805,
    5993 => 17808,
    5994 => 17811,
    5995 => 17813,
    5996 => 17816,
    5997 => 17819,
    5998 => 17821,
    5999 => 17824,
    6000 => 17827,
    6001 => 17829,
    6002 => 17832,
    6003 => 17834,
    6004 => 17837,
    6005 => 17840,
    6006 => 17842,
    6007 => 17845,
    6008 => 17848,
    6009 => 17850,
    6010 => 17853,
    6011 => 17855,
    6012 => 17858,
    6013 => 17861,
    6014 => 17863,
    6015 => 17866,
    6016 => 17869,
    6017 => 17871,
    6018 => 17874,
    6019 => 17877,
    6020 => 17879,
    6021 => 17882,
    6022 => 17884,
    6023 => 17887,
    6024 => 17890,
    6025 => 17892,
    6026 => 17895,
    6027 => 17898,
    6028 => 17900,
    6029 => 17903,
    6030 => 17906,
    6031 => 17908,
    6032 => 17911,
    6033 => 17913,
    6034 => 17916,
    6035 => 17919,
    6036 => 17921,
    6037 => 17924,
    6038 => 17927,
    6039 => 17929,
    6040 => 17932,
    6041 => 17934,
    6042 => 17937,
    6043 => 17940,
    6044 => 17942,
    6045 => 17945,
    6046 => 17948,
    6047 => 17950,
    6048 => 17953,
    6049 => 17955,
    6050 => 17958,
    6051 => 17961,
    6052 => 17963,
    6053 => 17966,
    6054 => 17969,
    6055 => 17971,
    6056 => 17974,
    6057 => 17976,
    6058 => 17979,
    6059 => 17982,
    6060 => 17984,
    6061 => 17987,
    6062 => 17990,
    6063 => 17992,
    6064 => 17995,
    6065 => 17997,
    6066 => 18000,
    6067 => 18003,
    6068 => 18005,
    6069 => 18008,
    6070 => 18011,
    6071 => 18013,
    6072 => 18016,
    6073 => 18018,
    6074 => 18021,
    6075 => 18024,
    6076 => 18026,
    6077 => 18029,
    6078 => 18032,
    6079 => 18034,
    6080 => 18037,
    6081 => 18039,
    6082 => 18042,
    6083 => 18045,
    6084 => 18047,
    6085 => 18050,
    6086 => 18053,
    6087 => 18055,
    6088 => 18058,
    6089 => 18060,
    6090 => 18063,
    6091 => 18066,
    6092 => 18068,
    6093 => 18071,
    6094 => 18074,
    6095 => 18076,
    6096 => 18079,
    6097 => 18081,
    6098 => 18084,
    6099 => 18087,
    6100 => 18089,
    6101 => 18092,
    6102 => 18095,
    6103 => 18097,
    6104 => 18100,
    6105 => 18102,
    6106 => 18105,
    6107 => 18108,
    6108 => 18110,
    6109 => 18113,
    6110 => 18115,
    6111 => 18118,
    6112 => 18121,
    6113 => 18123,
    6114 => 18126,
    6115 => 18129,
    6116 => 18131,
    6117 => 18134,
    6118 => 18136,
    6119 => 18139,
    6120 => 18142,
    6121 => 18144,
    6122 => 18147,
    6123 => 18149,
    6124 => 18152,
    6125 => 18155,
    6126 => 18157,
    6127 => 18160,
    6128 => 18163,
    6129 => 18165,
    6130 => 18168,
    6131 => 18170,
    6132 => 18173,
    6133 => 18176,
    6134 => 18178,
    6135 => 18181,
    6136 => 18183,
    6137 => 18186,
    6138 => 18189,
    6139 => 18191,
    6140 => 18194,
    6141 => 18197,
    6142 => 18199,
    6143 => 18202,
    6144 => 18204,
    6145 => 18207,
    6146 => 18210,
    6147 => 18212,
    6148 => 18215,
    6149 => 18217,
    6150 => 18220,
    6151 => 18223,
    6152 => 18225,
    6153 => 18228,
    6154 => 18230,
    6155 => 18233,
    6156 => 18236,
    6157 => 18238,
    6158 => 18241,
    6159 => 18244,
    6160 => 18246,
    6161 => 18249,
    6162 => 18251,
    6163 => 18254,
    6164 => 18257,
    6165 => 18259,
    6166 => 18262,
    6167 => 18264,
    6168 => 18267,
    6169 => 18270,
    6170 => 18272,
    6171 => 18275,
    6172 => 18277,
    6173 => 18280,
    6174 => 18283,
    6175 => 18285,
    6176 => 18288,
    6177 => 18290,
    6178 => 18293,
    6179 => 18296,
    6180 => 18298,
    6181 => 18301,
    6182 => 18304,
    6183 => 18306,
    6184 => 18309,
    6185 => 18311,
    6186 => 18314,
    6187 => 18317,
    6188 => 18319,
    6189 => 18322,
    6190 => 18324,
    6191 => 18327,
    6192 => 18330,
    6193 => 18332,
    6194 => 18335,
    6195 => 18337,
    6196 => 18340,
    6197 => 18343,
    6198 => 18345,
    6199 => 18348,
    6200 => 18350,
    6201 => 18353,
    6202 => 18356,
    6203 => 18358,
    6204 => 18361,
    6205 => 18363,
    6206 => 18366,
    6207 => 18369,
    6208 => 18371,
    6209 => 18374,
    6210 => 18376,
    6211 => 18379,
    6212 => 18382,
    6213 => 18384,
    6214 => 18387,
    6215 => 18389,
    6216 => 18392,
    6217 => 18395,
    6218 => 18397,
    6219 => 18400,
    6220 => 18402,
    6221 => 18405,
    6222 => 18408,
    6223 => 18410,
    6224 => 18413,
    6225 => 18415,
    6226 => 18418,
    6227 => 18421,
    6228 => 18423,
    6229 => 18426,
    6230 => 18428,
    6231 => 18431,
    6232 => 18434,
    6233 => 18436,
    6234 => 18439,
    6235 => 18441,
    6236 => 18444,
    6237 => 18447,
    6238 => 18449,
    6239 => 18452,
    6240 => 18454,
    6241 => 18457,
    6242 => 18460,
    6243 => 18462,
    6244 => 18465,
    6245 => 18467,
    6246 => 18470,
    6247 => 18473,
    6248 => 18475,
    6249 => 18478,
    6250 => 18480,
    6251 => 18483,
    6252 => 18485,
    6253 => 18488,
    6254 => 18491,
    6255 => 18493,
    6256 => 18496,
    6257 => 18498,
    6258 => 18501,
    6259 => 18504,
    6260 => 18506,
    6261 => 18509,
    6262 => 18511,
    6263 => 18514,
    6264 => 18517,
    6265 => 18519,
    6266 => 18522,
    6267 => 18524,
    6268 => 18527,
    6269 => 18530,
    6270 => 18532,
    6271 => 18535,
    6272 => 18537,
    6273 => 18540,
    6274 => 18543,
    6275 => 18545,
    6276 => 18548,
    6277 => 18550,
    6278 => 18553,
    6279 => 18555,
    6280 => 18558,
    6281 => 18561,
    6282 => 18563,
    6283 => 18566,
    6284 => 18568,
    6285 => 18571,
    6286 => 18574,
    6287 => 18576,
    6288 => 18579,
    6289 => 18581,
    6290 => 18584,
    6291 => 18587,
    6292 => 18589,
    6293 => 18592,
    6294 => 18594,
    6295 => 18597,
    6296 => 18599,
    6297 => 18602,
    6298 => 18605,
    6299 => 18607,
    6300 => 18610,
    6301 => 18612,
    6302 => 18615,
    6303 => 18618,
    6304 => 18620,
    6305 => 18623,
    6306 => 18625,
    6307 => 18628,
    6308 => 18630,
    6309 => 18633,
    6310 => 18636,
    6311 => 18638,
    6312 => 18641,
    6313 => 18643,
    6314 => 18646,
    6315 => 18649,
    6316 => 18651,
    6317 => 18654,
    6318 => 18656,
    6319 => 18659,
    6320 => 18661,
    6321 => 18664,
    6322 => 18667,
    6323 => 18669,
    6324 => 18672,
    6325 => 18674,
    6326 => 18677,
    6327 => 18680,
    6328 => 18682,
    6329 => 18685,
    6330 => 18687,
    6331 => 18690,
    6332 => 18692,
    6333 => 18695,
    6334 => 18698,
    6335 => 18700,
    6336 => 18703,
    6337 => 18705,
    6338 => 18708,
    6339 => 18711,
    6340 => 18713,
    6341 => 18716,
    6342 => 18718,
    6343 => 18721,
    6344 => 18723,
    6345 => 18726,
    6346 => 18729,
    6347 => 18731,
    6348 => 18734,
    6349 => 18736,
    6350 => 18739,
    6351 => 18741,
    6352 => 18744,
    6353 => 18747,
    6354 => 18749,
    6355 => 18752,
    6356 => 18754,
    6357 => 18757,
    6358 => 18759,
    6359 => 18762,
    6360 => 18765,
    6361 => 18767,
    6362 => 18770,
    6363 => 18772,
    6364 => 18775,
    6365 => 18778,
    6366 => 18780,
    6367 => 18783,
    6368 => 18785,
    6369 => 18788,
    6370 => 18790,
    6371 => 18793,
    6372 => 18796,
    6373 => 18798,
    6374 => 18801,
    6375 => 18803,
    6376 => 18806,
    6377 => 18808,
    6378 => 18811,
    6379 => 18814,
    6380 => 18816,
    6381 => 18819,
    6382 => 18821,
    6383 => 18824,
    6384 => 18826,
    6385 => 18829,
    6386 => 18832,
    6387 => 18834,
    6388 => 18837,
    6389 => 18839,
    6390 => 18842,
    6391 => 18844,
    6392 => 18847,
    6393 => 18850,
    6394 => 18852,
    6395 => 18855,
    6396 => 18857,
    6397 => 18860,
    6398 => 18862,
    6399 => 18865,
    6400 => 18868,
    6401 => 18870,
    6402 => 18873,
    6403 => 18875,
    6404 => 18878,
    6405 => 18880,
    6406 => 18883,
    6407 => 18885,
    6408 => 18888,
    6409 => 18891,
    6410 => 18893,
    6411 => 18896,
    6412 => 18898,
    6413 => 18901,
    6414 => 18903,
    6415 => 18906,
    6416 => 18909,
    6417 => 18911,
    6418 => 18914,
    6419 => 18916,
    6420 => 18919,
    6421 => 18921,
    6422 => 18924,
    6423 => 18927,
    6424 => 18929,
    6425 => 18932,
    6426 => 18934,
    6427 => 18937,
    6428 => 18939,
    6429 => 18942,
    6430 => 18944,
    6431 => 18947,
    6432 => 18950,
    6433 => 18952,
    6434 => 18955,
    6435 => 18957,
    6436 => 18960,
    6437 => 18962,
    6438 => 18965,
    6439 => 18968,
    6440 => 18970,
    6441 => 18973,
    6442 => 18975,
    6443 => 18978,
    6444 => 18980,
    6445 => 18983,
    6446 => 18985,
    6447 => 18988,
    6448 => 18991,
    6449 => 18993,
    6450 => 18996,
    6451 => 18998,
    6452 => 19001,
    6453 => 19003,
    6454 => 19006,
    6455 => 19009,
    6456 => 19011,
    6457 => 19014,
    6458 => 19016,
    6459 => 19019,
    6460 => 19021,
    6461 => 19024,
    6462 => 19026,
    6463 => 19029,
    6464 => 19032,
    6465 => 19034,
    6466 => 19037,
    6467 => 19039,
    6468 => 19042,
    6469 => 19044,
    6470 => 19047,
    6471 => 19049,
    6472 => 19052,
    6473 => 19055,
    6474 => 19057,
    6475 => 19060,
    6476 => 19062,
    6477 => 19065,
    6478 => 19067,
    6479 => 19070,
    6480 => 19072,
    6481 => 19075,
    6482 => 19078,
    6483 => 19080,
    6484 => 19083,
    6485 => 19085,
    6486 => 19088,
    6487 => 19090,
    6488 => 19093,
    6489 => 19095,
    6490 => 19098,
    6491 => 19101,
    6492 => 19103,
    6493 => 19106,
    6494 => 19108,
    6495 => 19111,
    6496 => 19113,
    6497 => 19116,
    6498 => 19118,
    6499 => 19121,
    6500 => 19123,
    6501 => 19126,
    6502 => 19129,
    6503 => 19131,
    6504 => 19134,
    6505 => 19136,
    6506 => 19139,
    6507 => 19141,
    6508 => 19144,
    6509 => 19146,
    6510 => 19149,
    6511 => 19152,
    6512 => 19154,
    6513 => 19157,
    6514 => 19159,
    6515 => 19162,
    6516 => 19164,
    6517 => 19167,
    6518 => 19169,
    6519 => 19172,
    6520 => 19174,
    6521 => 19177,
    6522 => 19180,
    6523 => 19182,
    6524 => 19185,
    6525 => 19187,
    6526 => 19190,
    6527 => 19192,
    6528 => 19195,
    6529 => 19197,
    6530 => 19200,
    6531 => 19202,
    6532 => 19205,
    6533 => 19208,
    6534 => 19210,
    6535 => 19213,
    6536 => 19215,
    6537 => 19218,
    6538 => 19220,
    6539 => 19223,
    6540 => 19225,
    6541 => 19228,
    6542 => 19230,
    6543 => 19233,
    6544 => 19236,
    6545 => 19238,
    6546 => 19241,
    6547 => 19243,
    6548 => 19246,
    6549 => 19248,
    6550 => 19251,
    6551 => 19253,
    6552 => 19256,
    6553 => 19258,
    6554 => 19261,
    6555 => 19264,
    6556 => 19266,
    6557 => 19269,
    6558 => 19271,
    6559 => 19274,
    6560 => 19276,
    6561 => 19279,
    6562 => 19281,
    6563 => 19284,
    6564 => 19286,
    6565 => 19289,
    6566 => 19291,
    6567 => 19294,
    6568 => 19297,
    6569 => 19299,
    6570 => 19302,
    6571 => 19304,
    6572 => 19307,
    6573 => 19309,
    6574 => 19312,
    6575 => 19314,
    6576 => 19317,
    6577 => 19319,
    6578 => 19322,
    6579 => 19324,
    6580 => 19327,
    6581 => 19330,
    6582 => 19332,
    6583 => 19335,
    6584 => 19337,
    6585 => 19340,
    6586 => 19342,
    6587 => 19345,
    6588 => 19347,
    6589 => 19350,
    6590 => 19352,
    6591 => 19355,
    6592 => 19357,
    6593 => 19360,
    6594 => 19362,
    6595 => 19365,
    6596 => 19368,
    6597 => 19370,
    6598 => 19373,
    6599 => 19375,
    6600 => 19378,
    6601 => 19380,
    6602 => 19383,
    6603 => 19385,
    6604 => 19388,
    6605 => 19390,
    6606 => 19393,
    6607 => 19395,
    6608 => 19398,
    6609 => 19400,
    6610 => 19403,
    6611 => 19406,
    6612 => 19408,
    6613 => 19411,
    6614 => 19413,
    6615 => 19416,
    6616 => 19418,
    6617 => 19421,
    6618 => 19423,
    6619 => 19426,
    6620 => 19428,
    6621 => 19431,
    6622 => 19433,
    6623 => 19436,
    6624 => 19438,
    6625 => 19441,
    6626 => 19444,
    6627 => 19446,
    6628 => 19449,
    6629 => 19451,
    6630 => 19454,
    6631 => 19456,
    6632 => 19459,
    6633 => 19461,
    6634 => 19464,
    6635 => 19466,
    6636 => 19469,
    6637 => 19471,
    6638 => 19474,
    6639 => 19476,
    6640 => 19479,
    6641 => 19481,
    6642 => 19484,
    6643 => 19486,
    6644 => 19489,
    6645 => 19492,
    6646 => 19494,
    6647 => 19497,
    6648 => 19499,
    6649 => 19502,
    6650 => 19504,
    6651 => 19507,
    6652 => 19509,
    6653 => 19512,
    6654 => 19514,
    6655 => 19517,
    6656 => 19519,
    6657 => 19522,
    6658 => 19524,
    6659 => 19527,
    6660 => 19529,
    6661 => 19532,
    6662 => 19534,
    6663 => 19537,
    6664 => 19539,
    6665 => 19542,
    6666 => 19545,
    6667 => 19547,
    6668 => 19550,
    6669 => 19552,
    6670 => 19555,
    6671 => 19557,
    6672 => 19560,
    6673 => 19562,
    6674 => 19565,
    6675 => 19567,
    6676 => 19570,
    6677 => 19572,
    6678 => 19575,
    6679 => 19577,
    6680 => 19580,
    6681 => 19582,
    6682 => 19585,
    6683 => 19587,
    6684 => 19590,
    6685 => 19592,
    6686 => 19595,
    6687 => 19597,
    6688 => 19600,
    6689 => 19602,
    6690 => 19605,
    6691 => 19607,
    6692 => 19610,
    6693 => 19613,
    6694 => 19615,
    6695 => 19618,
    6696 => 19620,
    6697 => 19623,
    6698 => 19625,
    6699 => 19628,
    6700 => 19630,
    6701 => 19633,
    6702 => 19635,
    6703 => 19638,
    6704 => 19640,
    6705 => 19643,
    6706 => 19645,
    6707 => 19648,
    6708 => 19650,
    6709 => 19653,
    6710 => 19655,
    6711 => 19658,
    6712 => 19660,
    6713 => 19663,
    6714 => 19665,
    6715 => 19668,
    6716 => 19670,
    6717 => 19673,
    6718 => 19675,
    6719 => 19678,
    6720 => 19680,
    6721 => 19683,
    6722 => 19685,
    6723 => 19688,
    6724 => 19690,
    6725 => 19693,
    6726 => 19695,
    6727 => 19698,
    6728 => 19700,
    6729 => 19703,
    6730 => 19706,
    6731 => 19708,
    6732 => 19711,
    6733 => 19713,
    6734 => 19716,
    6735 => 19718,
    6736 => 19721,
    6737 => 19723,
    6738 => 19726,
    6739 => 19728,
    6740 => 19731,
    6741 => 19733,
    6742 => 19736,
    6743 => 19738,
    6744 => 19741,
    6745 => 19743,
    6746 => 19746,
    6747 => 19748,
    6748 => 19751,
    6749 => 19753,
    6750 => 19756,
    6751 => 19758,
    6752 => 19761,
    6753 => 19763,
    6754 => 19766,
    6755 => 19768,
    6756 => 19771,
    6757 => 19773,
    6758 => 19776,
    6759 => 19778,
    6760 => 19781,
    6761 => 19783,
    6762 => 19786,
    6763 => 19788,
    6764 => 19791,
    6765 => 19793,
    6766 => 19796,
    6767 => 19798,
    6768 => 19801,
    6769 => 19803,
    6770 => 19806,
    6771 => 19808,
    6772 => 19811,
    6773 => 19813,
    6774 => 19816,
    6775 => 19818,
    6776 => 19821,
    6777 => 19823,
    6778 => 19826,
    6779 => 19828,
    6780 => 19831,
    6781 => 19833,
    6782 => 19836,
    6783 => 19838,
    6784 => 19841,
    6785 => 19843,
    6786 => 19846,
    6787 => 19848,
    6788 => 19851,
    6789 => 19853,
    6790 => 19856,
    6791 => 19858,
    6792 => 19861,
    6793 => 19863,
    6794 => 19866,
    6795 => 19868,
    6796 => 19871,
    6797 => 19873,
    6798 => 19876,
    6799 => 19878,
    6800 => 19881,
    6801 => 19883,
    6802 => 19886,
    6803 => 19888,
    6804 => 19891,
    6805 => 19893,
    6806 => 19896,
    6807 => 19898,
    6808 => 19901,
    6809 => 19903,
    6810 => 19906,
    6811 => 19908,
    6812 => 19911,
    6813 => 19913,
    6814 => 19916,
    6815 => 19918,
    6816 => 19921,
    6817 => 19923,
    6818 => 19926,
    6819 => 19928,
    6820 => 19931,
    6821 => 19933,
    6822 => 19936,
    6823 => 19938,
    6824 => 19941,
    6825 => 19943,
    6826 => 19946,
    6827 => 19948,
    6828 => 19951,
    6829 => 19953,
    6830 => 19956,
    6831 => 19958,
    6832 => 19961,
    6833 => 19963,
    6834 => 19966,
    6835 => 19968,
    6836 => 19971,
    6837 => 19973,
    6838 => 19976,
    6839 => 19978,
    6840 => 19981,
    6841 => 19983,
    6842 => 19985,
    6843 => 19988,
    6844 => 19990,
    6845 => 19993,
    6846 => 19995,
    6847 => 19998,
    6848 => 20000,
    6849 => 20003,
    6850 => 20005,
    6851 => 20008,
    6852 => 20010,
    6853 => 20013,
    6854 => 20015,
    6855 => 20018,
    6856 => 20020,
    6857 => 20023,
    6858 => 20025,
    6859 => 20028,
    6860 => 20030,
    6861 => 20033,
    6862 => 20035,
    6863 => 20038,
    6864 => 20040,
    6865 => 20043,
    6866 => 20045,
    6867 => 20048,
    6868 => 20050,
    6869 => 20053,
    6870 => 20055,
    6871 => 20058,
    6872 => 20060,
    6873 => 20063,
    6874 => 20065,
    6875 => 20068,
    6876 => 20070,
    6877 => 20072,
    6878 => 20075,
    6879 => 20077,
    6880 => 20080,
    6881 => 20082,
    6882 => 20085,
    6883 => 20087,
    6884 => 20090,
    6885 => 20092,
    6886 => 20095,
    6887 => 20097,
    6888 => 20100,
    6889 => 20102,
    6890 => 20105,
    6891 => 20107,
    6892 => 20110,
    6893 => 20112,
    6894 => 20115,
    6895 => 20117,
    6896 => 20120,
    6897 => 20122,
    6898 => 20125,
    6899 => 20127,
    6900 => 20130,
    6901 => 20132,
    6902 => 20135,
    6903 => 20137,
    6904 => 20139,
    6905 => 20142,
    6906 => 20144,
    6907 => 20147,
    6908 => 20149,
    6909 => 20152,
    6910 => 20154,
    6911 => 20157,
    6912 => 20159,
    6913 => 20162,
    6914 => 20164,
    6915 => 20167,
    6916 => 20169,
    6917 => 20172,
    6918 => 20174,
    6919 => 20177,
    6920 => 20179,
    6921 => 20182,
    6922 => 20184,
    6923 => 20187,
    6924 => 20189,
    6925 => 20191,
    6926 => 20194,
    6927 => 20196,
    6928 => 20199,
    6929 => 20201,
    6930 => 20204,
    6931 => 20206,
    6932 => 20209,
    6933 => 20211,
    6934 => 20214,
    6935 => 20216,
    6936 => 20219,
    6937 => 20221,
    6938 => 20224,
    6939 => 20226,
    6940 => 20229,
    6941 => 20231,
    6942 => 20234,
    6943 => 20236,
    6944 => 20238,
    6945 => 20241,
    6946 => 20243,
    6947 => 20246,
    6948 => 20248,
    6949 => 20251,
    6950 => 20253,
    6951 => 20256,
    6952 => 20258,
    6953 => 20261,
    6954 => 20263,
    6955 => 20266,
    6956 => 20268,
    6957 => 20271,
    6958 => 20273,
    6959 => 20275,
    6960 => 20278,
    6961 => 20280,
    6962 => 20283,
    6963 => 20285,
    6964 => 20288,
    6965 => 20290,
    6966 => 20293,
    6967 => 20295,
    6968 => 20298,
    6969 => 20300,
    6970 => 20303,
    6971 => 20305,
    6972 => 20308,
    6973 => 20310,
    6974 => 20312,
    6975 => 20315,
    6976 => 20317,
    6977 => 20320,
    6978 => 20322,
    6979 => 20325,
    6980 => 20327,
    6981 => 20330,
    6982 => 20332,
    6983 => 20335,
    6984 => 20337,
    6985 => 20340,
    6986 => 20342,
    6987 => 20345,
    6988 => 20347,
    6989 => 20349,
    6990 => 20352,
    6991 => 20354,
    6992 => 20357,
    6993 => 20359,
    6994 => 20362,
    6995 => 20364,
    6996 => 20367,
    6997 => 20369,
    6998 => 20372,
    6999 => 20374,
    7000 => 20377,
    7001 => 20379,
    7002 => 20381,
    7003 => 20384,
    7004 => 20386,
    7005 => 20389,
    7006 => 20391,
    7007 => 20394,
    7008 => 20396,
    7009 => 20399,
    7010 => 20401,
    7011 => 20404,
    7012 => 20406,
    7013 => 20408,
    7014 => 20411,
    7015 => 20413,
    7016 => 20416,
    7017 => 20418,
    7018 => 20421,
    7019 => 20423,
    7020 => 20426,
    7021 => 20428,
    7022 => 20431,
    7023 => 20433,
    7024 => 20436,
    7025 => 20438,
    7026 => 20440,
    7027 => 20443,
    7028 => 20445,
    7029 => 20448,
    7030 => 20450,
    7031 => 20453,
    7032 => 20455,
    7033 => 20458,
    7034 => 20460,
    7035 => 20463,
    7036 => 20465,
    7037 => 20467,
    7038 => 20470,
    7039 => 20472,
    7040 => 20475,
    7041 => 20477,
    7042 => 20480,
    7043 => 20482,
    7044 => 20485,
    7045 => 20487,
    7046 => 20489,
    7047 => 20492,
    7048 => 20494,
    7049 => 20497,
    7050 => 20499,
    7051 => 20502,
    7052 => 20504,
    7053 => 20507,
    7054 => 20509,
    7055 => 20512,
    7056 => 20514,
    7057 => 20516,
    7058 => 20519,
    7059 => 20521,
    7060 => 20524,
    7061 => 20526,
    7062 => 20529,
    7063 => 20531,
    7064 => 20534,
    7065 => 20536,
    7066 => 20538,
    7067 => 20541,
    7068 => 20543,
    7069 => 20546,
    7070 => 20548,
    7071 => 20551,
    7072 => 20553,
    7073 => 20556,
    7074 => 20558,
    7075 => 20560,
    7076 => 20563,
    7077 => 20565,
    7078 => 20568,
    7079 => 20570,
    7080 => 20573,
    7081 => 20575,
    7082 => 20578,
    7083 => 20580,
    7084 => 20583,
    7085 => 20585,
    7086 => 20587,
    7087 => 20590,
    7088 => 20592,
    7089 => 20595,
    7090 => 20597,
    7091 => 20600,
    7092 => 20602,
    7093 => 20604,
    7094 => 20607,
    7095 => 20609,
    7096 => 20612,
    7097 => 20614,
    7098 => 20617,
    7099 => 20619,
    7100 => 20622,
    7101 => 20624,
    7102 => 20626,
    7103 => 20629,
    7104 => 20631,
    7105 => 20634,
    7106 => 20636,
    7107 => 20639,
    7108 => 20641,
    7109 => 20644,
    7110 => 20646,
    7111 => 20648,
    7112 => 20651,
    7113 => 20653,
    7114 => 20656,
    7115 => 20658,
    7116 => 20661,
    7117 => 20663,
    7118 => 20666,
    7119 => 20668,
    7120 => 20670,
    7121 => 20673,
    7122 => 20675,
    7123 => 20678,
    7124 => 20680,
    7125 => 20683,
    7126 => 20685,
    7127 => 20687,
    7128 => 20690,
    7129 => 20692,
    7130 => 20695,
    7131 => 20697,
    7132 => 20700,
    7133 => 20702,
    7134 => 20704,
    7135 => 20707,
    7136 => 20709,
    7137 => 20712,
    7138 => 20714,
    7139 => 20717,
    7140 => 20719,
    7141 => 20722,
    7142 => 20724,
    7143 => 20726,
    7144 => 20729,
    7145 => 20731,
    7146 => 20734,
    7147 => 20736,
    7148 => 20739,
    7149 => 20741,
    7150 => 20743,
    7151 => 20746,
    7152 => 20748,
    7153 => 20751,
    7154 => 20753,
    7155 => 20756,
    7156 => 20758,
    7157 => 20760,
    7158 => 20763,
    7159 => 20765,
    7160 => 20768,
    7161 => 20770,
    7162 => 20773,
    7163 => 20775,
    7164 => 20777,
    7165 => 20780,
    7166 => 20782,
    7167 => 20785,
    7168 => 20787,
    7169 => 20790,
    7170 => 20792,
    7171 => 20794,
    7172 => 20797,
    7173 => 20799,
    7174 => 20802,
    7175 => 20804,
    7176 => 20807,
    7177 => 20809,
    7178 => 20811,
    7179 => 20814,
    7180 => 20816,
    7181 => 20819,
    7182 => 20821,
    7183 => 20824,
    7184 => 20826,
    7185 => 20828,
    7186 => 20831,
    7187 => 20833,
    7188 => 20836,
    7189 => 20838,
    7190 => 20841,
    7191 => 20843,
    7192 => 20845,
    7193 => 20848,
    7194 => 20850,
    7195 => 20853,
    7196 => 20855,
    7197 => 20858,
    7198 => 20860,
    7199 => 20862,
    7200 => 20865,
    7201 => 20867,
    7202 => 20870,
    7203 => 20872,
    7204 => 20874,
    7205 => 20877,
    7206 => 20879,
    7207 => 20882,
    7208 => 20884,
    7209 => 20887,
    7210 => 20889,
    7211 => 20891,
    7212 => 20894,
    7213 => 20896,
    7214 => 20899,
    7215 => 20901,
    7216 => 20904,
    7217 => 20906,
    7218 => 20908,
    7219 => 20911,
    7220 => 20913,
    7221 => 20916,
    7222 => 20918,
    7223 => 20920,
    7224 => 20923,
    7225 => 20925,
    7226 => 20928,
    7227 => 20930,
    7228 => 20933,
    7229 => 20935,
    7230 => 20937,
    7231 => 20940,
    7232 => 20942,
    7233 => 20945,
    7234 => 20947,
    7235 => 20949,
    7236 => 20952,
    7237 => 20954,
    7238 => 20957,
    7239 => 20959,
    7240 => 20962,
    7241 => 20964,
    7242 => 20966,
    7243 => 20969,
    7244 => 20971,
    7245 => 20974,
    7246 => 20976,
    7247 => 20978,
    7248 => 20981,
    7249 => 20983,
    7250 => 20986,
    7251 => 20988,
    7252 => 20990,
    7253 => 20993,
    7254 => 20995,
    7255 => 20998,
    7256 => 21000,
    7257 => 21003,
    7258 => 21005,
    7259 => 21007,
    7260 => 21010,
    7261 => 21012,
    7262 => 21015,
    7263 => 21017,
    7264 => 21019,
    7265 => 21022,
    7266 => 21024,
    7267 => 21027,
    7268 => 21029,
    7269 => 21031,
    7270 => 21034,
    7271 => 21036,
    7272 => 21039,
    7273 => 21041,
    7274 => 21043,
    7275 => 21046,
    7276 => 21048,
    7277 => 21051,
    7278 => 21053,
    7279 => 21056,
    7280 => 21058,
    7281 => 21060,
    7282 => 21063,
    7283 => 21065,
    7284 => 21068,
    7285 => 21070,
    7286 => 21072,
    7287 => 21075,
    7288 => 21077,
    7289 => 21080,
    7290 => 21082,
    7291 => 21084,
    7292 => 21087,
    7293 => 21089,
    7294 => 21092,
    7295 => 21094,
    7296 => 21096,
    7297 => 21099,
    7298 => 21101,
    7299 => 21104,
    7300 => 21106,
    7301 => 21108,
    7302 => 21111,
    7303 => 21113,
    7304 => 21116,
    7305 => 21118,
    7306 => 21120,
    7307 => 21123,
    7308 => 21125,
    7309 => 21128,
    7310 => 21130,
    7311 => 21132,
    7312 => 21135,
    7313 => 21137,
    7314 => 21140,
    7315 => 21142,
    7316 => 21144,
    7317 => 21147,
    7318 => 21149,
    7319 => 21152,
    7320 => 21154,
    7321 => 21156,
    7322 => 21159,
    7323 => 21161,
    7324 => 21164,
    7325 => 21166,
    7326 => 21168,
    7327 => 21171,
    7328 => 21173,
    7329 => 21176,
    7330 => 21178,
    7331 => 21180,
    7332 => 21183,
    7333 => 21185,
    7334 => 21188,
    7335 => 21190,
    7336 => 21192,
    7337 => 21195,
    7338 => 21197,
    7339 => 21200,
    7340 => 21202,
    7341 => 21204,
    7342 => 21207,
    7343 => 21209,
    7344 => 21212,
    7345 => 21214,
    7346 => 21216,
    7347 => 21219,
    7348 => 21221,
    7349 => 21224,
    7350 => 21226,
    7351 => 21228,
    7352 => 21231,
    7353 => 21233,
    7354 => 21236,
    7355 => 21238,
    7356 => 21240,
    7357 => 21243,
    7358 => 21245,
    7359 => 21247,
    7360 => 21250,
    7361 => 21252,
    7362 => 21255,
    7363 => 21257,
    7364 => 21259,
    7365 => 21262,
    7366 => 21264,
    7367 => 21267,
    7368 => 21269,
    7369 => 21271,
    7370 => 21274,
    7371 => 21276,
    7372 => 21279,
    7373 => 21281,
    7374 => 21283,
    7375 => 21286,
    7376 => 21288,
    7377 => 21290,
    7378 => 21293,
    7379 => 21295,
    7380 => 21298,
    7381 => 21300,
    7382 => 21302,
    7383 => 21305,
    7384 => 21307,
    7385 => 21310,
    7386 => 21312,
    7387 => 21314,
    7388 => 21317,
    7389 => 21319,
    7390 => 21322,
    7391 => 21324,
    7392 => 21326,
    7393 => 21329,
    7394 => 21331,
    7395 => 21333,
    7396 => 21336,
    7397 => 21338,
    7398 => 21341,
    7399 => 21343,
    7400 => 21345,
    7401 => 21348,
    7402 => 21350,
    7403 => 21353,
    7404 => 21355,
    7405 => 21357,
    7406 => 21360,
    7407 => 21362,
    7408 => 21364,
    7409 => 21367,
    7410 => 21369,
    7411 => 21372,
    7412 => 21374,
    7413 => 21376,
    7414 => 21379,
    7415 => 21381,
    7416 => 21383,
    7417 => 21386,
    7418 => 21388,
    7419 => 21391,
    7420 => 21393,
    7421 => 21395,
    7422 => 21398,
    7423 => 21400,
    7424 => 21403,
    7425 => 21405,
    7426 => 21407,
    7427 => 21410,
    7428 => 21412,
    7429 => 21414,
    7430 => 21417,
    7431 => 21419,
    7432 => 21422,
    7433 => 21424,
    7434 => 21426,
    7435 => 21429,
    7436 => 21431,
    7437 => 21433,
    7438 => 21436,
    7439 => 21438,
    7440 => 21441,
    7441 => 21443,
    7442 => 21445,
    7443 => 21448,
    7444 => 21450,
    7445 => 21452,
    7446 => 21455,
    7447 => 21457,
    7448 => 21460,
    7449 => 21462,
    7450 => 21464,
    7451 => 21467,
    7452 => 21469,
    7453 => 21471,
    7454 => 21474,
    7455 => 21476,
    7456 => 21479,
    7457 => 21481,
    7458 => 21483,
    7459 => 21486,
    7460 => 21488,
    7461 => 21490,
    7462 => 21493,
    7463 => 21495,
    7464 => 21498,
    7465 => 21500,
    7466 => 21502,
    7467 => 21505,
    7468 => 21507,
    7469 => 21509,
    7470 => 21512,
    7471 => 21514,
    7472 => 21516,
    7473 => 21519,
    7474 => 21521,
    7475 => 21524,
    7476 => 21526,
    7477 => 21528,
    7478 => 21531,
    7479 => 21533,
    7480 => 21535,
    7481 => 21538,
    7482 => 21540,
    7483 => 21543,
    7484 => 21545,
    7485 => 21547,
    7486 => 21550,
    7487 => 21552,
    7488 => 21554,
    7489 => 21557,
    7490 => 21559,
    7491 => 21561,
    7492 => 21564,
    7493 => 21566,
    7494 => 21569,
    7495 => 21571,
    7496 => 21573,
    7497 => 21576,
    7498 => 21578,
    7499 => 21580,
    7500 => 21583,
    7501 => 21585,
    7502 => 21587,
    7503 => 21590,
    7504 => 21592,
    7505 => 21595,
    7506 => 21597,
    7507 => 21599,
    7508 => 21602,
    7509 => 21604,
    7510 => 21606,
    7511 => 21609,
    7512 => 21611,
    7513 => 21613,
    7514 => 21616,
    7515 => 21618,
    7516 => 21621,
    7517 => 21623,
    7518 => 21625,
    7519 => 21628,
    7520 => 21630,
    7521 => 21632,
    7522 => 21635,
    7523 => 21637,
    7524 => 21639,
    7525 => 21642,
    7526 => 21644,
    7527 => 21646,
    7528 => 21649,
    7529 => 21651,
    7530 => 21654,
    7531 => 21656,
    7532 => 21658,
    7533 => 21661,
    7534 => 21663,
    7535 => 21665,
    7536 => 21668,
    7537 => 21670,
    7538 => 21672,
    7539 => 21675,
    7540 => 21677,
    7541 => 21679,
    7542 => 21682,
    7543 => 21684,
    7544 => 21687,
    7545 => 21689,
    7546 => 21691,
    7547 => 21694,
    7548 => 21696,
    7549 => 21698,
    7550 => 21701,
    7551 => 21703,
    7552 => 21705,
    7553 => 21708,
    7554 => 21710,
    7555 => 21712,
    7556 => 21715,
    7557 => 21717,
    7558 => 21719,
    7559 => 21722,
    7560 => 21724,
    7561 => 21727,
    7562 => 21729,
    7563 => 21731,
    7564 => 21734,
    7565 => 21736,
    7566 => 21738,
    7567 => 21741,
    7568 => 21743,
    7569 => 21745,
    7570 => 21748,
    7571 => 21750,
    7572 => 21752,
    7573 => 21755,
    7574 => 21757,
    7575 => 21759,
    7576 => 21762,
    7577 => 21764,
    7578 => 21766,
    7579 => 21769,
    7580 => 21771,
    7581 => 21774,
    7582 => 21776,
    7583 => 21778,
    7584 => 21781,
    7585 => 21783,
    7586 => 21785,
    7587 => 21788,
    7588 => 21790,
    7589 => 21792,
    7590 => 21795,
    7591 => 21797,
    7592 => 21799,
    7593 => 21802,
    7594 => 21804,
    7595 => 21806,
    7596 => 21809,
    7597 => 21811,
    7598 => 21813,
    7599 => 21816,
    7600 => 21818,
    7601 => 21820,
    7602 => 21823,
    7603 => 21825,
    7604 => 21827,
    7605 => 21830,
    7606 => 21832,
    7607 => 21835,
    7608 => 21837,
    7609 => 21839,
    7610 => 21842,
    7611 => 21844,
    7612 => 21846,
    7613 => 21849,
    7614 => 21851,
    7615 => 21853,
    7616 => 21856,
    7617 => 21858,
    7618 => 21860,
    7619 => 21863,
    7620 => 21865,
    7621 => 21867,
    7622 => 21870,
    7623 => 21872,
    7624 => 21874,
    7625 => 21877,
    7626 => 21879,
    7627 => 21881,
    7628 => 21884,
    7629 => 21886,
    7630 => 21888,
    7631 => 21891,
    7632 => 21893,
    7633 => 21895,
    7634 => 21898,
    7635 => 21900,
    7636 => 21902,
    7637 => 21905,
    7638 => 21907,
    7639 => 21909,
    7640 => 21912,
    7641 => 21914,
    7642 => 21916,
    7643 => 21919,
    7644 => 21921,
    7645 => 21923,
    7646 => 21926,
    7647 => 21928,
    7648 => 21930,
    7649 => 21933,
    7650 => 21935,
    7651 => 21937,
    7652 => 21940,
    7653 => 21942,
    7654 => 21944,
    7655 => 21947,
    7656 => 21949,
    7657 => 21951,
    7658 => 21954,
    7659 => 21956,
    7660 => 21958,
    7661 => 21961,
    7662 => 21963,
    7663 => 21965,
    7664 => 21968,
    7665 => 21970,
    7666 => 21972,
    7667 => 21975,
    7668 => 21977,
    7669 => 21979,
    7670 => 21982,
    7671 => 21984,
    7672 => 21986,
    7673 => 21989,
    7674 => 21991,
    7675 => 21993,
    7676 => 21996,
    7677 => 21998,
    7678 => 22000,
    7679 => 22003,
    7680 => 22005,
    7681 => 22007,
    7682 => 22010,
    7683 => 22012,
    7684 => 22014,
    7685 => 22017,
    7686 => 22019,
    7687 => 22021,
    7688 => 22024,
    7689 => 22026,
    7690 => 22028,
    7691 => 22031,
    7692 => 22033,
    7693 => 22035,
    7694 => 22038,
    7695 => 22040,
    7696 => 22042,
    7697 => 22045,
    7698 => 22047,
    7699 => 22049,
    7700 => 22051,
    7701 => 22054,
    7702 => 22056,
    7703 => 22058,
    7704 => 22061,
    7705 => 22063,
    7706 => 22065,
    7707 => 22068,
    7708 => 22070,
    7709 => 22072,
    7710 => 22075,
    7711 => 22077,
    7712 => 22079,
    7713 => 22082,
    7714 => 22084,
    7715 => 22086,
    7716 => 22089,
    7717 => 22091,
    7718 => 22093,
    7719 => 22096,
    7720 => 22098,
    7721 => 22100,
    7722 => 22103,
    7723 => 22105,
    7724 => 22107,
    7725 => 22110,
    7726 => 22112,
    7727 => 22114,
    7728 => 22116,
    7729 => 22119,
    7730 => 22121,
    7731 => 22123,
    7732 => 22126,
    7733 => 22128,
    7734 => 22130,
    7735 => 22133,
    7736 => 22135,
    7737 => 22137,
    7738 => 22140,
    7739 => 22142,
    7740 => 22144,
    7741 => 22147,
    7742 => 22149,
    7743 => 22151,
    7744 => 22154,
    7745 => 22156,
    7746 => 22158,
    7747 => 22160,
    7748 => 22163,
    7749 => 22165,
    7750 => 22167,
    7751 => 22170,
    7752 => 22172,
    7753 => 22174,
    7754 => 22177,
    7755 => 22179,
    7756 => 22181,
    7757 => 22184,
    7758 => 22186,
    7759 => 22188,
    7760 => 22191,
    7761 => 22193,
    7762 => 22195,
    7763 => 22197,
    7764 => 22200,
    7765 => 22202,
    7766 => 22204,
    7767 => 22207,
    7768 => 22209,
    7769 => 22211,
    7770 => 22214,
    7771 => 22216,
    7772 => 22218,
    7773 => 22221,
    7774 => 22223,
    7775 => 22225,
    7776 => 22227,
    7777 => 22230,
    7778 => 22232,
    7779 => 22234,
    7780 => 22237,
    7781 => 22239,
    7782 => 22241,
    7783 => 22244,
    7784 => 22246,
    7785 => 22248,
    7786 => 22251,
    7787 => 22253,
    7788 => 22255,
    7789 => 22257,
    7790 => 22260,
    7791 => 22262,
    7792 => 22264,
    7793 => 22267,
    7794 => 22269,
    7795 => 22271,
    7796 => 22274,
    7797 => 22276,
    7798 => 22278,
    7799 => 22281,
    7800 => 22283,
    7801 => 22285,
    7802 => 22287,
    7803 => 22290,
    7804 => 22292,
    7805 => 22294,
    7806 => 22297,
    7807 => 22299,
    7808 => 22301,
    7809 => 22304,
    7810 => 22306,
    7811 => 22308,
    7812 => 22310,
    7813 => 22313,
    7814 => 22315,
    7815 => 22317,
    7816 => 22320,
    7817 => 22322,
    7818 => 22324,
    7819 => 22327,
    7820 => 22329,
    7821 => 22331,
    7822 => 22333,
    7823 => 22336,
    7824 => 22338,
    7825 => 22340,
    7826 => 22343,
    7827 => 22345,
    7828 => 22347,
    7829 => 22350,
    7830 => 22352,
    7831 => 22354,
    7832 => 22356,
    7833 => 22359,
    7834 => 22361,
    7835 => 22363,
    7836 => 22366,
    7837 => 22368,
    7838 => 22370,
    7839 => 22373,
    7840 => 22375,
    7841 => 22377,
    7842 => 22379,
    7843 => 22382,
    7844 => 22384,
    7845 => 22386,
    7846 => 22389,
    7847 => 22391,
    7848 => 22393,
    7849 => 22395,
    7850 => 22398,
    7851 => 22400,
    7852 => 22402,
    7853 => 22405,
    7854 => 22407,
    7855 => 22409,
    7856 => 22411,
    7857 => 22414,
    7858 => 22416,
    7859 => 22418,
    7860 => 22421,
    7861 => 22423,
    7862 => 22425,
    7863 => 22428,
    7864 => 22430,
    7865 => 22432,
    7866 => 22434,
    7867 => 22437,
    7868 => 22439,
    7869 => 22441,
    7870 => 22444,
    7871 => 22446,
    7872 => 22448,
    7873 => 22450,
    7874 => 22453,
    7875 => 22455,
    7876 => 22457,
    7877 => 22460,
    7878 => 22462,
    7879 => 22464,
    7880 => 22466,
    7881 => 22469,
    7882 => 22471,
    7883 => 22473,
    7884 => 22476,
    7885 => 22478,
    7886 => 22480,
    7887 => 22482,
    7888 => 22485,
    7889 => 22487,
    7890 => 22489,
    7891 => 22492,
    7892 => 22494,
    7893 => 22496,
    7894 => 22498,
    7895 => 22501,
    7896 => 22503,
    7897 => 22505,
    7898 => 22508,
    7899 => 22510,
    7900 => 22512,
    7901 => 22514,
    7902 => 22517,
    7903 => 22519,
    7904 => 22521,
    7905 => 22524,
    7906 => 22526,
    7907 => 22528,
    7908 => 22530,
    7909 => 22533,
    7910 => 22535,
    7911 => 22537,
    7912 => 22540,
    7913 => 22542,
    7914 => 22544,
    7915 => 22546,
    7916 => 22549,
    7917 => 22551,
    7918 => 22553,
    7919 => 22555,
    7920 => 22558,
    7921 => 22560,
    7922 => 22562,
    7923 => 22565,
    7924 => 22567,
    7925 => 22569,
    7926 => 22571,
    7927 => 22574,
    7928 => 22576,
    7929 => 22578,
    7930 => 22581,
    7931 => 22583,
    7932 => 22585,
    7933 => 22587,
    7934 => 22590,
    7935 => 22592,
    7936 => 22594,
    7937 => 22596,
    7938 => 22599,
    7939 => 22601,
    7940 => 22603,
    7941 => 22606,
    7942 => 22608,
    7943 => 22610,
    7944 => 22612,
    7945 => 22615,
    7946 => 22617,
    7947 => 22619,
    7948 => 22621,
    7949 => 22624,
    7950 => 22626,
    7951 => 22628,
    7952 => 22631,
    7953 => 22633,
    7954 => 22635,
    7955 => 22637,
    7956 => 22640,
    7957 => 22642,
    7958 => 22644,
    7959 => 22646,
    7960 => 22649,
    7961 => 22651,
    7962 => 22653,
    7963 => 22656,
    7964 => 22658,
    7965 => 22660,
    7966 => 22662,
    7967 => 22665,
    7968 => 22667,
    7969 => 22669,
    7970 => 22671,
    7971 => 22674,
    7972 => 22676,
    7973 => 22678,
    7974 => 22680,
    7975 => 22683,
    7976 => 22685,
    7977 => 22687,
    7978 => 22690,
    7979 => 22692,
    7980 => 22694,
    7981 => 22696,
    7982 => 22699,
    7983 => 22701,
    7984 => 22703,
    7985 => 22705,
    7986 => 22708,
    7987 => 22710,
    7988 => 22712,
    7989 => 22714,
    7990 => 22717,
    7991 => 22719,
    7992 => 22721,
    7993 => 22724,
    7994 => 22726,
    7995 => 22728,
    7996 => 22730,
    7997 => 22733,
    7998 => 22735,
    7999 => 22737,
    8000 => 22739,
    8001 => 22742,
    8002 => 22744,
    8003 => 22746,
    8004 => 22748,
    8005 => 22751,
    8006 => 22753,
    8007 => 22755,
    8008 => 22757,
    8009 => 22760,
    8010 => 22762,
    8011 => 22764,
    8012 => 22766,
    8013 => 22769,
    8014 => 22771,
    8015 => 22773,
    8016 => 22776,
    8017 => 22778,
    8018 => 22780,
    8019 => 22782,
    8020 => 22785,
    8021 => 22787,
    8022 => 22789,
    8023 => 22791,
    8024 => 22794,
    8025 => 22796,
    8026 => 22798,
    8027 => 22800,
    8028 => 22803,
    8029 => 22805,
    8030 => 22807,
    8031 => 22809,
    8032 => 22812,
    8033 => 22814,
    8034 => 22816,
    8035 => 22818,
    8036 => 22821,
    8037 => 22823,
    8038 => 22825,
    8039 => 22827,
    8040 => 22830,
    8041 => 22832,
    8042 => 22834,
    8043 => 22836,
    8044 => 22839,
    8045 => 22841,
    8046 => 22843,
    8047 => 22845,
    8048 => 22848,
    8049 => 22850,
    8050 => 22852,
    8051 => 22854,
    8052 => 22857,
    8053 => 22859,
    8054 => 22861,
    8055 => 22863,
    8056 => 22866,
    8057 => 22868,
    8058 => 22870,
    8059 => 22872,
    8060 => 22875,
    8061 => 22877,
    8062 => 22879,
    8063 => 22881,
    8064 => 22884,
    8065 => 22886,
    8066 => 22888,
    8067 => 22890,
    8068 => 22893,
    8069 => 22895,
    8070 => 22897,
    8071 => 22899,
    8072 => 22902,
    8073 => 22904,
    8074 => 22906,
    8075 => 22908,
    8076 => 22911,
    8077 => 22913,
    8078 => 22915,
    8079 => 22917,
    8080 => 22920,
    8081 => 22922,
    8082 => 22924,
    8083 => 22926,
    8084 => 22929,
    8085 => 22931,
    8086 => 22933,
    8087 => 22935,
    8088 => 22938,
    8089 => 22940,
    8090 => 22942,
    8091 => 22944,
    8092 => 22947,
    8093 => 22949,
    8094 => 22951,
    8095 => 22953,
    8096 => 22956,
    8097 => 22958,
    8098 => 22960,
    8099 => 22962,
    8100 => 22965,
    8101 => 22967,
    8102 => 22969,
    8103 => 22971,
    8104 => 22973,
    8105 => 22976,
    8106 => 22978,
    8107 => 22980,
    8108 => 22982,
    8109 => 22985,
    8110 => 22987,
    8111 => 22989,
    8112 => 22991,
    8113 => 22994,
    8114 => 22996,
    8115 => 22998,
    8116 => 23000,
    8117 => 23003,
    8118 => 23005,
    8119 => 23007,
    8120 => 23009,
    8121 => 23012,
    8122 => 23014,
    8123 => 23016,
    8124 => 23018,
    8125 => 23020,
    8126 => 23023,
    8127 => 23025,
    8128 => 23027,
    8129 => 23029,
    8130 => 23032,
    8131 => 23034,
    8132 => 23036,
    8133 => 23038,
    8134 => 23041,
    8135 => 23043,
    8136 => 23045,
    8137 => 23047,
    8138 => 23050,
    8139 => 23052,
    8140 => 23054,
    8141 => 23056,
    8142 => 23058,
    8143 => 23061,
    8144 => 23063,
    8145 => 23065,
    8146 => 23067,
    8147 => 23070,
    8148 => 23072,
    8149 => 23074,
    8150 => 23076,
    8151 => 23079,
    8152 => 23081,
    8153 => 23083,
    8154 => 23085,
    8155 => 23087,
    8156 => 23090,
    8157 => 23092,
    8158 => 23094,
    8159 => 23096,
    8160 => 23099,
    8161 => 23101,
    8162 => 23103,
    8163 => 23105,
    8164 => 23107,
    8165 => 23110,
    8166 => 23112,
    8167 => 23114,
    8168 => 23116,
    8169 => 23119,
    8170 => 23121,
    8171 => 23123,
    8172 => 23125,
    8173 => 23128,
    8174 => 23130,
    8175 => 23132,
    8176 => 23134,
    8177 => 23136,
    8178 => 23139,
    8179 => 23141,
    8180 => 23143,
    8181 => 23145,
    8182 => 23148,
    8183 => 23150,
    8184 => 23152,
    8185 => 23154,
    8186 => 23156,
    8187 => 23159,
    8188 => 23161,
    8189 => 23163,
    8190 => 23165,
    8191 => 23168,
    8192 => 23170,
    8193 => 23172,
    8194 => 23174,
    8195 => 23176,
    8196 => 23179,
    8197 => 23181,
    8198 => 23183,
    8199 => 23185,
    8200 => 23188,
    8201 => 23190,
    8202 => 23192,
    8203 => 23194,
    8204 => 23196,
    8205 => 23199,
    8206 => 23201,
    8207 => 23203,
    8208 => 23205,
    8209 => 23208,
    8210 => 23210,
    8211 => 23212,
    8212 => 23214,
    8213 => 23216,
    8214 => 23219,
    8215 => 23221,
    8216 => 23223,
    8217 => 23225,
    8218 => 23227,
    8219 => 23230,
    8220 => 23232,
    8221 => 23234,
    8222 => 23236,
    8223 => 23239,
    8224 => 23241,
    8225 => 23243,
    8226 => 23245,
    8227 => 23247,
    8228 => 23250,
    8229 => 23252,
    8230 => 23254,
    8231 => 23256,
    8232 => 23258,
    8233 => 23261,
    8234 => 23263,
    8235 => 23265,
    8236 => 23267,
    8237 => 23270,
    8238 => 23272,
    8239 => 23274,
    8240 => 23276,
    8241 => 23278,
    8242 => 23281,
    8243 => 23283,
    8244 => 23285,
    8245 => 23287,
    8246 => 23289,
    8247 => 23292,
    8248 => 23294,
    8249 => 23296,
    8250 => 23298,
    8251 => 23300,
    8252 => 23303,
    8253 => 23305,
    8254 => 23307,
    8255 => 23309,
    8256 => 23311,
    8257 => 23314,
    8258 => 23316,
    8259 => 23318,
    8260 => 23320,
    8261 => 23323,
    8262 => 23325,
    8263 => 23327,
    8264 => 23329,
    8265 => 23331,
    8266 => 23334,
    8267 => 23336,
    8268 => 23338,
    8269 => 23340,
    8270 => 23342,
    8271 => 23345,
    8272 => 23347,
    8273 => 23349,
    8274 => 23351,
    8275 => 23353,
    8276 => 23356,
    8277 => 23358,
    8278 => 23360,
    8279 => 23362,
    8280 => 23364,
    8281 => 23367,
    8282 => 23369,
    8283 => 23371,
    8284 => 23373,
    8285 => 23375,
    8286 => 23378,
    8287 => 23380,
    8288 => 23382,
    8289 => 23384,
    8290 => 23386,
    8291 => 23389,
    8292 => 23391,
    8293 => 23393,
    8294 => 23395,
    8295 => 23397,
    8296 => 23400,
    8297 => 23402,
    8298 => 23404,
    8299 => 23406,
    8300 => 23408,
    8301 => 23411,
    8302 => 23413,
    8303 => 23415,
    8304 => 23417,
    8305 => 23419,
    8306 => 23422,
    8307 => 23424,
    8308 => 23426,
    8309 => 23428,
    8310 => 23430,
    8311 => 23433,
    8312 => 23435,
    8313 => 23437,
    8314 => 23439,
    8315 => 23441,
    8316 => 23444,
    8317 => 23446,
    8318 => 23448,
    8319 => 23450,
    8320 => 23452,
    8321 => 23455,
    8322 => 23457,
    8323 => 23459,
    8324 => 23461,
    8325 => 23463,
    8326 => 23466,
    8327 => 23468,
    8328 => 23470,
    8329 => 23472,
    8330 => 23474,
    8331 => 23476,
    8332 => 23479,
    8333 => 23481,
    8334 => 23483,
    8335 => 23485,
    8336 => 23487,
    8337 => 23490,
    8338 => 23492,
    8339 => 23494,
    8340 => 23496,
    8341 => 23498,
    8342 => 23501,
    8343 => 23503,
    8344 => 23505,
    8345 => 23507,
    8346 => 23509,
    8347 => 23512,
    8348 => 23514,
    8349 => 23516,
    8350 => 23518,
    8351 => 23520,
    8352 => 23522,
    8353 => 23525,
    8354 => 23527,
    8355 => 23529,
    8356 => 23531,
    8357 => 23533,
    8358 => 23536,
    8359 => 23538,
    8360 => 23540,
    8361 => 23542,
    8362 => 23544,
    8363 => 23546,
    8364 => 23549,
    8365 => 23551,
    8366 => 23553,
    8367 => 23555,
    8368 => 23557,
    8369 => 23560,
    8370 => 23562,
    8371 => 23564,
    8372 => 23566,
    8373 => 23568,
    8374 => 23571,
    8375 => 23573,
    8376 => 23575,
    8377 => 23577,
    8378 => 23579,
    8379 => 23581,
    8380 => 23584,
    8381 => 23586,
    8382 => 23588,
    8383 => 23590,
    8384 => 23592,
    8385 => 23595,
    8386 => 23597,
    8387 => 23599,
    8388 => 23601,
    8389 => 23603,
    8390 => 23605,
    8391 => 23608,
    8392 => 23610,
    8393 => 23612,
    8394 => 23614,
    8395 => 23616,
    8396 => 23618,
    8397 => 23621,
    8398 => 23623,
    8399 => 23625,
    8400 => 23627,
    8401 => 23629,
    8402 => 23632,
    8403 => 23634,
    8404 => 23636,
    8405 => 23638,
    8406 => 23640,
    8407 => 23642,
    8408 => 23645,
    8409 => 23647,
    8410 => 23649,
    8411 => 23651,
    8412 => 23653,
    8413 => 23655,
    8414 => 23658,
    8415 => 23660,
    8416 => 23662,
    8417 => 23664,
    8418 => 23666,
    8419 => 23668,
    8420 => 23671,
    8421 => 23673,
    8422 => 23675,
    8423 => 23677,
    8424 => 23679,
    8425 => 23682,
    8426 => 23684,
    8427 => 23686,
    8428 => 23688,
    8429 => 23690,
    8430 => 23692,
    8431 => 23695,
    8432 => 23697,
    8433 => 23699,
    8434 => 23701,
    8435 => 23703,
    8436 => 23705,
    8437 => 23708,
    8438 => 23710,
    8439 => 23712,
    8440 => 23714,
    8441 => 23716,
    8442 => 23718,
    8443 => 23721,
    8444 => 23723,
    8445 => 23725,
    8446 => 23727,
    8447 => 23729,
    8448 => 23731,
    8449 => 23734,
    8450 => 23736,
    8451 => 23738,
    8452 => 23740,
    8453 => 23742,
    8454 => 23744,
    8455 => 23747,
    8456 => 23749,
    8457 => 23751,
    8458 => 23753,
    8459 => 23755,
    8460 => 23757,
    8461 => 23760,
    8462 => 23762,
    8463 => 23764,
    8464 => 23766,
    8465 => 23768,
    8466 => 23770,
    8467 => 23773,
    8468 => 23775,
    8469 => 23777,
    8470 => 23779,
    8471 => 23781,
    8472 => 23783,
    8473 => 23785,
    8474 => 23788,
    8475 => 23790,
    8476 => 23792,
    8477 => 23794,
    8478 => 23796,
    8479 => 23798,
    8480 => 23801,
    8481 => 23803,
    8482 => 23805,
    8483 => 23807,
    8484 => 23809,
    8485 => 23811,
    8486 => 23814,
    8487 => 23816,
    8488 => 23818,
    8489 => 23820,
    8490 => 23822,
    8491 => 23824,
    8492 => 23827,
    8493 => 23829,
    8494 => 23831,
    8495 => 23833,
    8496 => 23835,
    8497 => 23837,
    8498 => 23839,
    8499 => 23842,
    8500 => 23844,
    8501 => 23846,
    8502 => 23848,
    8503 => 23850,
    8504 => 23852,
    8505 => 23855,
    8506 => 23857,
    8507 => 23859,
    8508 => 23861,
    8509 => 23863,
    8510 => 23865,
    8511 => 23867,
    8512 => 23870,
    8513 => 23872,
    8514 => 23874,
    8515 => 23876,
    8516 => 23878,
    8517 => 23880,
    8518 => 23883,
    8519 => 23885,
    8520 => 23887,
    8521 => 23889,
    8522 => 23891,
    8523 => 23893,
    8524 => 23895,
    8525 => 23898,
    8526 => 23900,
    8527 => 23902,
    8528 => 23904,
    8529 => 23906,
    8530 => 23908,
    8531 => 23910,
    8532 => 23913,
    8533 => 23915,
    8534 => 23917,
    8535 => 23919,
    8536 => 23921,
    8537 => 23923,
    8538 => 23925,
    8539 => 23928,
    8540 => 23930,
    8541 => 23932,
    8542 => 23934,
    8543 => 23936,
    8544 => 23938,
    8545 => 23940,
    8546 => 23943,
    8547 => 23945,
    8548 => 23947,
    8549 => 23949,
    8550 => 23951,
    8551 => 23953,
    8552 => 23956,
    8553 => 23958,
    8554 => 23960,
    8555 => 23962,
    8556 => 23964,
    8557 => 23966,
    8558 => 23968,
    8559 => 23971,
    8560 => 23973,
    8561 => 23975,
    8562 => 23977,
    8563 => 23979,
    8564 => 23981,
    8565 => 23983,
    8566 => 23985,
    8567 => 23988,
    8568 => 23990,
    8569 => 23992,
    8570 => 23994,
    8571 => 23996,
    8572 => 23998,
    8573 => 24000,
    8574 => 24003,
    8575 => 24005,
    8576 => 24007,
    8577 => 24009,
    8578 => 24011,
    8579 => 24013,
    8580 => 24015,
    8581 => 24018,
    8582 => 24020,
    8583 => 24022,
    8584 => 24024,
    8585 => 24026,
    8586 => 24028,
    8587 => 24030,
    8588 => 24033,
    8589 => 24035,
    8590 => 24037,
    8591 => 24039,
    8592 => 24041,
    8593 => 24043,
    8594 => 24045,
    8595 => 24047,
    8596 => 24050,
    8597 => 24052,
    8598 => 24054,
    8599 => 24056,
    8600 => 24058,
    8601 => 24060,
    8602 => 24062,
    8603 => 24065,
    8604 => 24067,
    8605 => 24069,
    8606 => 24071,
    8607 => 24073,
    8608 => 24075,
    8609 => 24077,
    8610 => 24079,
    8611 => 24082,
    8612 => 24084,
    8613 => 24086,
    8614 => 24088,
    8615 => 24090,
    8616 => 24092,
    8617 => 24094,
    8618 => 24096,
    8619 => 24099,
    8620 => 24101,
    8621 => 24103,
    8622 => 24105,
    8623 => 24107,
    8624 => 24109,
    8625 => 24111,
    8626 => 24114,
    8627 => 24116,
    8628 => 24118,
    8629 => 24120,
    8630 => 24122,
    8631 => 24124,
    8632 => 24126,
    8633 => 24128,
    8634 => 24131,
    8635 => 24133,
    8636 => 24135,
    8637 => 24137,
    8638 => 24139,
    8639 => 24141,
    8640 => 24143,
    8641 => 24145,
    8642 => 24148,
    8643 => 24150,
    8644 => 24152,
    8645 => 24154,
    8646 => 24156,
    8647 => 24158,
    8648 => 24160,
    8649 => 24162,
    8650 => 24164,
    8651 => 24167,
    8652 => 24169,
    8653 => 24171,
    8654 => 24173,
    8655 => 24175,
    8656 => 24177,
    8657 => 24179,
    8658 => 24181,
    8659 => 24184,
    8660 => 24186,
    8661 => 24188,
    8662 => 24190,
    8663 => 24192,
    8664 => 24194,
    8665 => 24196,
    8666 => 24198,
    8667 => 24201,
    8668 => 24203,
    8669 => 24205,
    8670 => 24207,
    8671 => 24209,
    8672 => 24211,
    8673 => 24213,
    8674 => 24215,
    8675 => 24217,
    8676 => 24220,
    8677 => 24222,
    8678 => 24224,
    8679 => 24226,
    8680 => 24228,
    8681 => 24230,
    8682 => 24232,
    8683 => 24234,
    8684 => 24237,
    8685 => 24239,
    8686 => 24241,
    8687 => 24243,
    8688 => 24245,
    8689 => 24247,
    8690 => 24249,
    8691 => 24251,
    8692 => 24253,
    8693 => 24256,
    8694 => 24258,
    8695 => 24260,
    8696 => 24262,
    8697 => 24264,
    8698 => 24266,
    8699 => 24268,
    8700 => 24270,
    8701 => 24272,
    8702 => 24275,
    8703 => 24277,
    8704 => 24279,
    8705 => 24281,
    8706 => 24283,
    8707 => 24285,
    8708 => 24287,
    8709 => 24289,
    8710 => 24291,
    8711 => 24294,
    8712 => 24296,
    8713 => 24298,
    8714 => 24300,
    8715 => 24302,
    8716 => 24304,
    8717 => 24306,
    8718 => 24308,
    8719 => 24310,
    8720 => 24312,
    8721 => 24315,
    8722 => 24317,
    8723 => 24319,
    8724 => 24321,
    8725 => 24323,
    8726 => 24325,
    8727 => 24327,
    8728 => 24329,
    8729 => 24331,
    8730 => 24334,
    8731 => 24336,
    8732 => 24338,
    8733 => 24340,
    8734 => 24342,
    8735 => 24344,
    8736 => 24346,
    8737 => 24348,
    8738 => 24350,
    8739 => 24352,
    8740 => 24355,
    8741 => 24357,
    8742 => 24359,
    8743 => 24361,
    8744 => 24363,
    8745 => 24365,
    8746 => 24367,
    8747 => 24369,
    8748 => 24371,
    8749 => 24373,
    8750 => 24376,
    8751 => 24378,
    8752 => 24380,
    8753 => 24382,
    8754 => 24384,
    8755 => 24386,
    8756 => 24388,
    8757 => 24390,
    8758 => 24392,
    8759 => 24394,
    8760 => 24397,
    8761 => 24399,
    8762 => 24401,
    8763 => 24403,
    8764 => 24405,
    8765 => 24407,
    8766 => 24409,
    8767 => 24411,
    8768 => 24413,
    8769 => 24415,
    8770 => 24417,
    8771 => 24420,
    8772 => 24422,
    8773 => 24424,
    8774 => 24426,
    8775 => 24428,
    8776 => 24430,
    8777 => 24432,
    8778 => 24434,
    8779 => 24436,
    8780 => 24438,
    8781 => 24441,
    8782 => 24443,
    8783 => 24445,
    8784 => 24447,
    8785 => 24449,
    8786 => 24451,
    8787 => 24453,
    8788 => 24455,
    8789 => 24457,
    8790 => 24459,
    8791 => 24461,
    8792 => 24464,
    8793 => 24466,
    8794 => 24468,
    8795 => 24470,
    8796 => 24472,
    8797 => 24474,
    8798 => 24476,
    8799 => 24478,
    8800 => 24480,
    8801 => 24482,
    8802 => 24484,
    8803 => 24487,
    8804 => 24489,
    8805 => 24491,
    8806 => 24493,
    8807 => 24495,
    8808 => 24497,
    8809 => 24499,
    8810 => 24501,
    8811 => 24503,
    8812 => 24505,
    8813 => 24507,
    8814 => 24509,
    8815 => 24512,
    8816 => 24514,
    8817 => 24516,
    8818 => 24518,
    8819 => 24520,
    8820 => 24522,
    8821 => 24524,
    8822 => 24526,
    8823 => 24528,
    8824 => 24530,
    8825 => 24532,
    8826 => 24534,
    8827 => 24537,
    8828 => 24539,
    8829 => 24541,
    8830 => 24543,
    8831 => 24545,
    8832 => 24547,
    8833 => 24549,
    8834 => 24551,
    8835 => 24553,
    8836 => 24555,
    8837 => 24557,
    8838 => 24559,
    8839 => 24562,
    8840 => 24564,
    8841 => 24566,
    8842 => 24568,
    8843 => 24570,
    8844 => 24572,
    8845 => 24574,
    8846 => 24576,
    8847 => 24578,
    8848 => 24580,
    8849 => 24582,
    8850 => 24584,
    8851 => 24586,
    8852 => 24589,
    8853 => 24591,
    8854 => 24593,
    8855 => 24595,
    8856 => 24597,
    8857 => 24599,
    8858 => 24601,
    8859 => 24603,
    8860 => 24605,
    8861 => 24607,
    8862 => 24609,
    8863 => 24611,
    8864 => 24613,
    8865 => 24616,
    8866 => 24618,
    8867 => 24620,
    8868 => 24622,
    8869 => 24624,
    8870 => 24626,
    8871 => 24628,
    8872 => 24630,
    8873 => 24632,
    8874 => 24634,
    8875 => 24636,
    8876 => 24638,
    8877 => 24640,
    8878 => 24642,
    8879 => 24645,
    8880 => 24647,
    8881 => 24649,
    8882 => 24651,
    8883 => 24653,
    8884 => 24655,
    8885 => 24657,
    8886 => 24659,
    8887 => 24661,
    8888 => 24663,
    8889 => 24665,
    8890 => 24667,
    8891 => 24669,
    8892 => 24671,
    8893 => 24673,
    8894 => 24676,
    8895 => 24678,
    8896 => 24680,
    8897 => 24682,
    8898 => 24684,
    8899 => 24686,
    8900 => 24688,
    8901 => 24690,
    8902 => 24692,
    8903 => 24694,
    8904 => 24696,
    8905 => 24698,
    8906 => 24700,
    8907 => 24702,
    8908 => 24704,
    8909 => 24707,
    8910 => 24709,
    8911 => 24711,
    8912 => 24713,
    8913 => 24715,
    8914 => 24717,
    8915 => 24719,
    8916 => 24721,
    8917 => 24723,
    8918 => 24725,
    8919 => 24727,
    8920 => 24729,
    8921 => 24731,
    8922 => 24733,
    8923 => 24735,
    8924 => 24737,
    8925 => 24740,
    8926 => 24742,
    8927 => 24744,
    8928 => 24746,
    8929 => 24748,
    8930 => 24750,
    8931 => 24752,
    8932 => 24754,
    8933 => 24756,
    8934 => 24758,
    8935 => 24760,
    8936 => 24762,
    8937 => 24764,
    8938 => 24766,
    8939 => 24768,
    8940 => 24770,
    8941 => 24772,
    8942 => 24774,
    8943 => 24777,
    8944 => 24779,
    8945 => 24781,
    8946 => 24783,
    8947 => 24785,
    8948 => 24787,
    8949 => 24789,
    8950 => 24791,
    8951 => 24793,
    8952 => 24795,
    8953 => 24797,
    8954 => 24799,
    8955 => 24801,
    8956 => 24803,
    8957 => 24805,
    8958 => 24807,
    8959 => 24809,
    8960 => 24811,
    8961 => 24814,
    8962 => 24816,
    8963 => 24818,
    8964 => 24820,
    8965 => 24822,
    8966 => 24824,
    8967 => 24826,
    8968 => 24828,
    8969 => 24830,
    8970 => 24832,
    8971 => 24834,
    8972 => 24836,
    8973 => 24838,
    8974 => 24840,
    8975 => 24842,
    8976 => 24844,
    8977 => 24846,
    8978 => 24848,
    8979 => 24850,
    8980 => 24852,
    8981 => 24855,
    8982 => 24857,
    8983 => 24859,
    8984 => 24861,
    8985 => 24863,
    8986 => 24865,
    8987 => 24867,
    8988 => 24869,
    8989 => 24871,
    8990 => 24873,
    8991 => 24875,
    8992 => 24877,
    8993 => 24879,
    8994 => 24881,
    8995 => 24883,
    8996 => 24885,
    8997 => 24887,
    8998 => 24889,
    8999 => 24891,
    9000 => 24893,
    9001 => 24895,
    9002 => 24897,
    9003 => 24899,
    9004 => 24902,
    9005 => 24904,
    9006 => 24906,
    9007 => 24908,
    9008 => 24910,
    9009 => 24912,
    9010 => 24914,
    9011 => 24916,
    9012 => 24918,
    9013 => 24920,
    9014 => 24922,
    9015 => 24924,
    9016 => 24926,
    9017 => 24928,
    9018 => 24930,
    9019 => 24932,
    9020 => 24934,
    9021 => 24936,
    9022 => 24938,
    9023 => 24940,
    9024 => 24942,
    9025 => 24944,
    9026 => 24946,
    9027 => 24948,
    9028 => 24950,
    9029 => 24953,
    9030 => 24955,
    9031 => 24957,
    9032 => 24959,
    9033 => 24961,
    9034 => 24963,
    9035 => 24965,
    9036 => 24967,
    9037 => 24969,
    9038 => 24971,
    9039 => 24973,
    9040 => 24975,
    9041 => 24977,
    9042 => 24979,
    9043 => 24981,
    9044 => 24983,
    9045 => 24985,
    9046 => 24987,
    9047 => 24989,
    9048 => 24991,
    9049 => 24993,
    9050 => 24995,
    9051 => 24997,
    9052 => 24999,
    9053 => 25001,
    9054 => 25003,
    9055 => 25005,
    9056 => 25007,
    9057 => 25009,
    9058 => 25011,
    9059 => 25013,
    9060 => 25016,
    9061 => 25018,
    9062 => 25020,
    9063 => 25022,
    9064 => 25024,
    9065 => 25026,
    9066 => 25028,
    9067 => 25030,
    9068 => 25032,
    9069 => 25034,
    9070 => 25036,
    9071 => 25038,
    9072 => 25040,
    9073 => 25042,
    9074 => 25044,
    9075 => 25046,
    9076 => 25048,
    9077 => 25050,
    9078 => 25052,
    9079 => 25054,
    9080 => 25056,
    9081 => 25058,
    9082 => 25060,
    9083 => 25062,
    9084 => 25064,
    9085 => 25066,
    9086 => 25068,
    9087 => 25070,
    9088 => 25072,
    9089 => 25074,
    9090 => 25076,
    9091 => 25078,
    9092 => 25080,
    9093 => 25082,
    9094 => 25084,
    9095 => 25086,
    9096 => 25088,
    9097 => 25090,
    9098 => 25092,
    9099 => 25094,
    9100 => 25096,
    9101 => 25099,
    9102 => 25101,
    9103 => 25103,
    9104 => 25105,
    9105 => 25107,
    9106 => 25109,
    9107 => 25111,
    9108 => 25113,
    9109 => 25115,
    9110 => 25117,
    9111 => 25119,
    9112 => 25121,
    9113 => 25123,
    9114 => 25125,
    9115 => 25127,
    9116 => 25129,
    9117 => 25131,
    9118 => 25133,
    9119 => 25135,
    9120 => 25137,
    9121 => 25139,
    9122 => 25141,
    9123 => 25143,
    9124 => 25145,
    9125 => 25147,
    9126 => 25149,
    9127 => 25151,
    9128 => 25153,
    9129 => 25155,
    9130 => 25157,
    9131 => 25159,
    9132 => 25161,
    9133 => 25163,
    9134 => 25165,
    9135 => 25167,
    9136 => 25169,
    9137 => 25171,
    9138 => 25173,
    9139 => 25175,
    9140 => 25177,
    9141 => 25179,
    9142 => 25181,
    9143 => 25183,
    9144 => 25185,
    9145 => 25187,
    9146 => 25189,
    9147 => 25191,
    9148 => 25193,
    9149 => 25195,
    9150 => 25197,
    9151 => 25199,
    9152 => 25201,
    9153 => 25203,
    9154 => 25205,
    9155 => 25207,
    9156 => 25209,
    9157 => 25211,
    9158 => 25213,
    9159 => 25215,
    9160 => 25217,
    9161 => 25219,
    9162 => 25221,
    9163 => 25223,
    9164 => 25225,
    9165 => 25227,
    9166 => 25229,
    9167 => 25231,
    9168 => 25233,
    9169 => 25235,
    9170 => 25237,
    9171 => 25239,
    9172 => 25241,
    9173 => 25243,
    9174 => 25245,
    9175 => 25247,
    9176 => 25249,
    9177 => 25251,
    9178 => 25253,
    9179 => 25255,
    9180 => 25257,
    9181 => 25259,
    9182 => 25261,
    9183 => 25263,
    9184 => 25265,
    9185 => 25267,
    9186 => 25269,
    9187 => 25271,
    9188 => 25273,
    9189 => 25275,
    9190 => 25277,
    9191 => 25279,
    9192 => 25281,
    9193 => 25283,
    9194 => 25285,
    9195 => 25287,
    9196 => 25289,
    9197 => 25291,
    9198 => 25293,
    9199 => 25295,
    9200 => 25297,
    9201 => 25299,
    9202 => 25301,
    9203 => 25303,
    9204 => 25305,
    9205 => 25307,
    9206 => 25309,
    9207 => 25311,
    9208 => 25313,
    9209 => 25315,
    9210 => 25317,
    9211 => 25319,
    9212 => 25321,
    9213 => 25323,
    9214 => 25325,
    9215 => 25327,
    9216 => 25329,
    9217 => 25331,
    9218 => 25333,
    9219 => 25335,
    9220 => 25337,
    9221 => 25339,
    9222 => 25341,
    9223 => 25343,
    9224 => 25345,
    9225 => 25347,
    9226 => 25349,
    9227 => 25351,
    9228 => 25353,
    9229 => 25355,
    9230 => 25357,
    9231 => 25359,
    9232 => 25361,
    9233 => 25363,
    9234 => 25365,
    9235 => 25367,
    9236 => 25369,
    9237 => 25371,
    9238 => 25373,
    9239 => 25375,
    9240 => 25377,
    9241 => 25379,
    9242 => 25381,
    9243 => 25383,
    9244 => 25385,
    9245 => 25387,
    9246 => 25389,
    9247 => 25391,
    9248 => 25393,
    9249 => 25395,
    9250 => 25397,
    9251 => 25399,
    9252 => 25401,
    9253 => 25403,
    9254 => 25405,
    9255 => 25407,
    9256 => 25409,
    9257 => 25411,
    9258 => 25413,
    9259 => 25415,
    9260 => 25417,
    9261 => 25419,
    9262 => 25421,
    9263 => 25423,
    9264 => 25425,
    9265 => 25427,
    9266 => 25429,
    9267 => 25431,
    9268 => 25433,
    9269 => 25435,
    9270 => 25437,
    9271 => 25438,
    9272 => 25440,
    9273 => 25442,
    9274 => 25444,
    9275 => 25446,
    9276 => 25448,
    9277 => 25450,
    9278 => 25452,
    9279 => 25454,
    9280 => 25456,
    9281 => 25458,
    9282 => 25460,
    9283 => 25462,
    9284 => 25464,
    9285 => 25466,
    9286 => 25468,
    9287 => 25470,
    9288 => 25472,
    9289 => 25474,
    9290 => 25476,
    9291 => 25478,
    9292 => 25480,
    9293 => 25482,
    9294 => 25484,
    9295 => 25486,
    9296 => 25488,
    9297 => 25490,
    9298 => 25492,
    9299 => 25494,
    9300 => 25496,
    9301 => 25498,
    9302 => 25500,
    9303 => 25502,
    9304 => 25504,
    9305 => 25506,
    9306 => 25508,
    9307 => 25510,
    9308 => 25512,
    9309 => 25514,
    9310 => 25516,
    9311 => 25518,
    9312 => 25519,
    9313 => 25521,
    9314 => 25523,
    9315 => 25525,
    9316 => 25527,
    9317 => 25529,
    9318 => 25531,
    9319 => 25533,
    9320 => 25535,
    9321 => 25537,
    9322 => 25539,
    9323 => 25541,
    9324 => 25543,
    9325 => 25545,
    9326 => 25547,
    9327 => 25549,
    9328 => 25551,
    9329 => 25553,
    9330 => 25555,
    9331 => 25557,
    9332 => 25559,
    9333 => 25561,
    9334 => 25563,
    9335 => 25565,
    9336 => 25567,
    9337 => 25569,
    9338 => 25571,
    9339 => 25573,
    9340 => 25575,
    9341 => 25577,
    9342 => 25578,
    9343 => 25580,
    9344 => 25582,
    9345 => 25584,
    9346 => 25586,
    9347 => 25588,
    9348 => 25590,
    9349 => 25592,
    9350 => 25594,
    9351 => 25596,
    9352 => 25598,
    9353 => 25600,
    9354 => 25602,
    9355 => 25604,
    9356 => 25606,
    9357 => 25608,
    9358 => 25610,
    9359 => 25612,
    9360 => 25614,
    9361 => 25616,
    9362 => 25618,
    9363 => 25620,
    9364 => 25622,
    9365 => 25624,
    9366 => 25626,
    9367 => 25628,
    9368 => 25629,
    9369 => 25631,
    9370 => 25633,
    9371 => 25635,
    9372 => 25637,
    9373 => 25639,
    9374 => 25641,
    9375 => 25643,
    9376 => 25645,
    9377 => 25647,
    9378 => 25649,
    9379 => 25651,
    9380 => 25653,
    9381 => 25655,
    9382 => 25657,
    9383 => 25659,
    9384 => 25661,
    9385 => 25663,
    9386 => 25665,
    9387 => 25667,
    9388 => 25669,
    9389 => 25671,
    9390 => 25672,
    9391 => 25674,
    9392 => 25676,
    9393 => 25678,
    9394 => 25680,
    9395 => 25682,
    9396 => 25684,
    9397 => 25686,
    9398 => 25688,
    9399 => 25690,
    9400 => 25692,
    9401 => 25694,
    9402 => 25696,
    9403 => 25698,
    9404 => 25700,
    9405 => 25702,
    9406 => 25704,
    9407 => 25706,
    9408 => 25708,
    9409 => 25710,
    9410 => 25711,
    9411 => 25713,
    9412 => 25715,
    9413 => 25717,
    9414 => 25719,
    9415 => 25721,
    9416 => 25723,
    9417 => 25725,
    9418 => 25727,
    9419 => 25729,
    9420 => 25731,
    9421 => 25733,
    9422 => 25735,
    9423 => 25737,
    9424 => 25739,
    9425 => 25741,
    9426 => 25743,
    9427 => 25745,
    9428 => 25746,
    9429 => 25748,
    9430 => 25750,
    9431 => 25752,
    9432 => 25754,
    9433 => 25756,
    9434 => 25758,
    9435 => 25760,
    9436 => 25762,
    9437 => 25764,
    9438 => 25766,
    9439 => 25768,
    9440 => 25770,
    9441 => 25772,
    9442 => 25774,
    9443 => 25776,
    9444 => 25778,
    9445 => 25779,
    9446 => 25781,
    9447 => 25783,
    9448 => 25785,
    9449 => 25787,
    9450 => 25789,
    9451 => 25791,
    9452 => 25793,
    9453 => 25795,
    9454 => 25797,
    9455 => 25799,
    9456 => 25801,
    9457 => 25803,
    9458 => 25805,
    9459 => 25807,
    9460 => 25809,
    9461 => 25810,
    9462 => 25812,
    9463 => 25814,
    9464 => 25816,
    9465 => 25818,
    9466 => 25820,
    9467 => 25822,
    9468 => 25824,
    9469 => 25826,
    9470 => 25828,
    9471 => 25830,
    9472 => 25832,
    9473 => 25834,
    9474 => 25836,
    9475 => 25838,
    9476 => 25839,
    9477 => 25841,
    9478 => 25843,
    9479 => 25845,
    9480 => 25847,
    9481 => 25849,
    9482 => 25851,
    9483 => 25853,
    9484 => 25855,
    9485 => 25857,
    9486 => 25859,
    9487 => 25861,
    9488 => 25863,
    9489 => 25865,
    9490 => 25866,
    9491 => 25868,
    9492 => 25870,
    9493 => 25872,
    9494 => 25874,
    9495 => 25876,
    9496 => 25878,
    9497 => 25880,
    9498 => 25882,
    9499 => 25884,
    9500 => 25886,
    9501 => 25888,
    9502 => 25890,
    9503 => 25892,
    9504 => 25893,
    9505 => 25895,
    9506 => 25897,
    9507 => 25899,
    9508 => 25901,
    9509 => 25903,
    9510 => 25905,
    9511 => 25907,
    9512 => 25909,
    9513 => 25911,
    9514 => 25913,
    9515 => 25915,
    9516 => 25917,
    9517 => 25918,
    9518 => 25920,
    9519 => 25922,
    9520 => 25924,
    9521 => 25926,
    9522 => 25928,
    9523 => 25930,
    9524 => 25932,
    9525 => 25934,
    9526 => 25936,
    9527 => 25938,
    9528 => 25940,
    9529 => 25942,
    9530 => 25943,
    9531 => 25945,
    9532 => 25947,
    9533 => 25949,
    9534 => 25951,
    9535 => 25953,
    9536 => 25955,
    9537 => 25957,
    9538 => 25959,
    9539 => 25961,
    9540 => 25963,
    9541 => 25965,
    9542 => 25966,
    9543 => 25968,
    9544 => 25970,
    9545 => 25972,
    9546 => 25974,
    9547 => 25976,
    9548 => 25978,
    9549 => 25980,
    9550 => 25982,
    9551 => 25984,
    9552 => 25986,
    9553 => 25988,
    9554 => 25989,
    9555 => 25991,
    9556 => 25993,
    9557 => 25995,
    9558 => 25997,
    9559 => 25999,
    9560 => 26001,
    9561 => 26003,
    9562 => 26005,
    9563 => 26007,
    9564 => 26009,
    9565 => 26010,
    9566 => 26012,
    9567 => 26014,
    9568 => 26016,
    9569 => 26018,
    9570 => 26020,
    9571 => 26022,
    9572 => 26024,
    9573 => 26026,
    9574 => 26028,
    9575 => 26030,
    9576 => 26031,
    9577 => 26033,
    9578 => 26035,
    9579 => 26037,
    9580 => 26039,
    9581 => 26041,
    9582 => 26043,
    9583 => 26045,
    9584 => 26047,
    9585 => 26049,
    9586 => 26051,
    9587 => 26052,
    9588 => 26054,
    9589 => 26056,
    9590 => 26058,
    9591 => 26060,
    9592 => 26062,
    9593 => 26064,
    9594 => 26066,
    9595 => 26068,
    9596 => 26070,
    9597 => 26071,
    9598 => 26073,
    9599 => 26075,
    9600 => 26077,
    9601 => 26079,
    9602 => 26081,
    9603 => 26083,
    9604 => 26085,
    9605 => 26087,
    9606 => 26089,
    9607 => 26090,
    9608 => 26092,
    9609 => 26094,
    9610 => 26096,
    9611 => 26098,
    9612 => 26100,
    9613 => 26102,
    9614 => 26104,
    9615 => 26106,
    9616 => 26108,
    9617 => 26109,
    9618 => 26111,
    9619 => 26113,
    9620 => 26115,
    9621 => 26117,
    9622 => 26119,
    9623 => 26121,
    9624 => 26123,
    9625 => 26125,
    9626 => 26127,
    9627 => 26128,
    9628 => 26130,
    9629 => 26132,
    9630 => 26134,
    9631 => 26136,
    9632 => 26138,
    9633 => 26140,
    9634 => 26142,
    9635 => 26144,
    9636 => 26146,
    9637 => 26147,
    9638 => 26149,
    9639 => 26151,
    9640 => 26153,
    9641 => 26155,
    9642 => 26157,
    9643 => 26159,
    9644 => 26161,
    9645 => 26163,
    9646 => 26164,
    9647 => 26166,
    9648 => 26168,
    9649 => 26170,
    9650 => 26172,
    9651 => 26174,
    9652 => 26176,
    9653 => 26178,
    9654 => 26180,
    9655 => 26181,
    9656 => 26183,
    9657 => 26185,
    9658 => 26187,
    9659 => 26189,
    9660 => 26191,
    9661 => 26193,
    9662 => 26195,
    9663 => 26197,
    9664 => 26198,
    9665 => 26200,
    9666 => 26202,
    9667 => 26204,
    9668 => 26206,
    9669 => 26208,
    9670 => 26210,
    9671 => 26212,
    9672 => 26214,
    9673 => 26215,
    9674 => 26217,
    9675 => 26219,
    9676 => 26221,
    9677 => 26223,
    9678 => 26225,
    9679 => 26227,
    9680 => 26229,
    9681 => 26230,
    9682 => 26232,
    9683 => 26234,
    9684 => 26236,
    9685 => 26238,
    9686 => 26240,
    9687 => 26242,
    9688 => 26244,
    9689 => 26246,
    9690 => 26247,
    9691 => 26249,
    9692 => 26251,
    9693 => 26253,
    9694 => 26255,
    9695 => 26257,
    9696 => 26259,
    9697 => 26261,
    9698 => 26262,
    9699 => 26264,
    9700 => 26266,
    9701 => 26268,
    9702 => 26270,
    9703 => 26272,
    9704 => 26274,
    9705 => 26276,
    9706 => 26277,
    9707 => 26279,
    9708 => 26281,
    9709 => 26283,
    9710 => 26285,
    9711 => 26287,
    9712 => 26289,
    9713 => 26291,
    9714 => 26292,
    9715 => 26294,
    9716 => 26296,
    9717 => 26298,
    9718 => 26300,
    9719 => 26302,
    9720 => 26304,
    9721 => 26306,
    9722 => 26307,
    9723 => 26309,
    9724 => 26311,
    9725 => 26313,
    9726 => 26315,
    9727 => 26317,
    9728 => 26319,
    9729 => 26321,
    9730 => 26322,
    9731 => 26324,
    9732 => 26326,
    9733 => 26328,
    9734 => 26330,
    9735 => 26332,
    9736 => 26334,
    9737 => 26336,
    9738 => 26337,
    9739 => 26339,
    9740 => 26341,
    9741 => 26343,
    9742 => 26345,
    9743 => 26347,
    9744 => 26349,
    9745 => 26350,
    9746 => 26352,
    9747 => 26354,
    9748 => 26356,
    9749 => 26358,
    9750 => 26360,
    9751 => 26362,
    9752 => 26364,
    9753 => 26365,
    9754 => 26367,
    9755 => 26369,
    9756 => 26371,
    9757 => 26373,
    9758 => 26375,
    9759 => 26377,
    9760 => 26378,
    9761 => 26380,
    9762 => 26382,
    9763 => 26384,
    9764 => 26386,
    9765 => 26388,
    9766 => 26390,
    9767 => 26392,
    9768 => 26393,
    9769 => 26395,
    9770 => 26397,
    9771 => 26399,
    9772 => 26401,
    9773 => 26403,
    9774 => 26405,
    9775 => 26406,
    9776 => 26408,
    9777 => 26410,
    9778 => 26412,
    9779 => 26414,
    9780 => 26416,
    9781 => 26418,
    9782 => 26419,
    9783 => 26421,
    9784 => 26423,
    9785 => 26425,
    9786 => 26427,
    9787 => 26429,
    9788 => 26431,
    9789 => 26432,
    9790 => 26434,
    9791 => 26436,
    9792 => 26438,
    9793 => 26440,
    9794 => 26442,
    9795 => 26444,
    9796 => 26445,
    9797 => 26447,
    9798 => 26449,
    9799 => 26451,
    9800 => 26453,
    9801 => 26455,
    9802 => 26457,
    9803 => 26458,
    9804 => 26460,
    9805 => 26462,
    9806 => 26464,
    9807 => 26466,
    9808 => 26468,
    9809 => 26469,
    9810 => 26471,
    9811 => 26473,
    9812 => 26475,
    9813 => 26477,
    9814 => 26479,
    9815 => 26481,
    9816 => 26482,
    9817 => 26484,
    9818 => 26486,
    9819 => 26488,
    9820 => 26490,
    9821 => 26492,
    9822 => 26494,
    9823 => 26495,
    9824 => 26497,
    9825 => 26499,
    9826 => 26501,
    9827 => 26503,
    9828 => 26505,
    9829 => 26506,
    9830 => 26508,
    9831 => 26510,
    9832 => 26512,
    9833 => 26514,
    9834 => 26516,
    9835 => 26518,
    9836 => 26519,
    9837 => 26521,
    9838 => 26523,
    9839 => 26525,
    9840 => 26527,
    9841 => 26529,
    9842 => 26530,
    9843 => 26532,
    9844 => 26534,
    9845 => 26536,
    9846 => 26538,
    9847 => 26540,
    9848 => 26542,
    9849 => 26543,
    9850 => 26545,
    9851 => 26547,
    9852 => 26549,
    9853 => 26551,
    9854 => 26553,
    9855 => 26554,
    9856 => 26556,
    9857 => 26558,
    9858 => 26560,
    9859 => 26562,
    9860 => 26564,
    9861 => 26565,
    9862 => 26567,
    9863 => 26569,
    9864 => 26571,
    9865 => 26573,
    9866 => 26575,
    9867 => 26576,
    9868 => 26578,
    9869 => 26580,
    9870 => 26582,
    9871 => 26584,
    9872 => 26586,
    9873 => 26588,
    9874 => 26589,
    9875 => 26591,
    9876 => 26593,
    9877 => 26595,
    9878 => 26597,
    9879 => 26599,
    9880 => 26600,
    9881 => 26602,
    9882 => 26604,
    9883 => 26606,
    9884 => 26608,
    9885 => 26610,
    9886 => 26611,
    9887 => 26613,
    9888 => 26615,
    9889 => 26617,
    9890 => 26619,
    9891 => 26621,
    9892 => 26622,
    9893 => 26624,
    9894 => 26626,
    9895 => 26628,
    9896 => 26630,
    9897 => 26631,
    9898 => 26633,
    9899 => 26635,
    9900 => 26637,
    9901 => 26639,
    9902 => 26641,
    9903 => 26642,
    9904 => 26644,
    9905 => 26646,
    9906 => 26648,
    9907 => 26650,
    9908 => 26652,
    9909 => 26653,
    9910 => 26655,
    9911 => 26657,
    9912 => 26659,
    9913 => 26661,
    9914 => 26663,
    9915 => 26664,
    9916 => 26666,
    9917 => 26668,
    9918 => 26670,
    9919 => 26672,
    9920 => 26674,
    9921 => 26675,
    9922 => 26677,
    9923 => 26679,
    9924 => 26681,
    9925 => 26683,
    9926 => 26684,
    9927 => 26686,
    9928 => 26688,
    9929 => 26690,
    9930 => 26692,
    9931 => 26694,
    9932 => 26695,
    9933 => 26697,
    9934 => 26699,
    9935 => 26701,
    9936 => 26703,
    9937 => 26705,
    9938 => 26706,
    9939 => 26708,
    9940 => 26710,
    9941 => 26712,
    9942 => 26714,
    9943 => 26715,
    9944 => 26717,
    9945 => 26719,
    9946 => 26721,
    9947 => 26723,
    9948 => 26725,
    9949 => 26726,
    9950 => 26728,
    9951 => 26730,
    9952 => 26732,
    9953 => 26734,
    9954 => 26735,
    9955 => 26737,
    9956 => 26739,
    9957 => 26741,
    9958 => 26743,
    9959 => 26745,
    9960 => 26746,
    9961 => 26748,
    9962 => 26750,
    9963 => 26752,
    9964 => 26754,
    9965 => 26755,
    9966 => 26757,
    9967 => 26759,
    9968 => 26761,
    9969 => 26763,
    9970 => 26764,
    9971 => 26766,
    9972 => 26768,
    9973 => 26770,
    9974 => 26772,
    9975 => 26774,
    9976 => 26775,
    9977 => 26777,
    9978 => 26779,
    9979 => 26781,
    9980 => 26783,
    9981 => 26784,
    9982 => 26786,
    9983 => 26788,
    9984 => 26790,
    9985 => 26792,
    9986 => 26793,
    9987 => 26795,
    9988 => 26797,
    9989 => 26799,
    9990 => 26801,
    9991 => 26802,
    9992 => 26804,
    9993 => 26806,
    9994 => 26808,
    9995 => 26810,
    9996 => 26811,
    9997 => 26813,
    9998 => 26815,
    9999 => 26817,
    10000 => 26819,
    10001 => 26821,
    10002 => 26822,
    10003 => 26824,
    10004 => 26826,
    10005 => 26828,
    10006 => 26830,
    10007 => 26831,
    10008 => 26833,
    10009 => 26835,
    10010 => 26837,
    10011 => 26839,
    10012 => 26840,
    10013 => 26842,
    10014 => 26844,
    10015 => 26846,
    10016 => 26848,
    10017 => 26849,
    10018 => 26851,
    10019 => 26853,
    10020 => 26855,
    10021 => 26857,
    10022 => 26858,
    10023 => 26860,
    10024 => 26862,
    10025 => 26864,
    10026 => 26866,
    10027 => 26867,
    10028 => 26869,
    10029 => 26871,
    10030 => 26873,
    10031 => 26875,
    10032 => 26876,
    10033 => 26878,
    10034 => 26880,
    10035 => 26882,
    10036 => 26884,
    10037 => 26885,
    10038 => 26887,
    10039 => 26889,
    10040 => 26891,
    10041 => 26893,
    10042 => 26894,
    10043 => 26896,
    10044 => 26898,
    10045 => 26900,
    10046 => 26901,
    10047 => 26903,
    10048 => 26905,
    10049 => 26907,
    10050 => 26909,
    10051 => 26910,
    10052 => 26912,
    10053 => 26914,
    10054 => 26916,
    10055 => 26918,
    10056 => 26919,
    10057 => 26921,
    10058 => 26923,
    10059 => 26925,
    10060 => 26927,
    10061 => 26928,
    10062 => 26930,
    10063 => 26932,
    10064 => 26934,
    10065 => 26936,
    10066 => 26937,
    10067 => 26939,
    10068 => 26941,
    10069 => 26943,
    10070 => 26944,
    10071 => 26946,
    10072 => 26948,
    10073 => 26950,
    10074 => 26952,
    10075 => 26953,
    10076 => 26955,
    10077 => 26957,
    10078 => 26959,
    10079 => 26961,
    10080 => 26962,
    10081 => 26964,
    10082 => 26966,
    10083 => 26968,
    10084 => 26969,
    10085 => 26971,
    10086 => 26973,
    10087 => 26975,
    10088 => 26977,
    10089 => 26978,
    10090 => 26980,
    10091 => 26982,
    10092 => 26984,
    10093 => 26986,
    10094 => 26987,
    10095 => 26989,
    10096 => 26991,
    10097 => 26993,
    10098 => 26994,
    10099 => 26996,
    10100 => 26998,
    10101 => 27000,
    10102 => 27002,
    10103 => 27003,
    10104 => 27005,
    10105 => 27007,
    10106 => 27009,
    10107 => 27010,
    10108 => 27012,
    10109 => 27014,
    10110 => 27016,
    10111 => 27018,
    10112 => 27019,
    10113 => 27021,
    10114 => 27023,
    10115 => 27025,
    10116 => 27026,
    10117 => 27028,
    10118 => 27030,
    10119 => 27032,
    10120 => 27034,
    10121 => 27035,
    10122 => 27037,
    10123 => 27039,
    10124 => 27041,
    10125 => 27042,
    10126 => 27044,
    10127 => 27046,
    10128 => 27048,
    10129 => 27049,
    10130 => 27051,
    10131 => 27053,
    10132 => 27055,
    10133 => 27057,
    10134 => 27058,
    10135 => 27060,
    10136 => 27062,
    10137 => 27064,
    10138 => 27065,
    10139 => 27067,
    10140 => 27069,
    10141 => 27071,
    10142 => 27073,
    10143 => 27074,
    10144 => 27076,
    10145 => 27078,
    10146 => 27080,
    10147 => 27081,
    10148 => 27083,
    10149 => 27085,
    10150 => 27087,
    10151 => 27088,
    10152 => 27090,
    10153 => 27092,
    10154 => 27094,
    10155 => 27096,
    10156 => 27097,
    10157 => 27099,
    10158 => 27101,
    10159 => 27103,
    10160 => 27104,
    10161 => 27106,
    10162 => 27108,
    10163 => 27110,
    10164 => 27111,
    10165 => 27113,
    10166 => 27115,
    10167 => 27117,
    10168 => 27118,
    10169 => 27120,
    10170 => 27122,
    10171 => 27124,
    10172 => 27126,
    10173 => 27127,
    10174 => 27129,
    10175 => 27131,
    10176 => 27133,
    10177 => 27134,
    10178 => 27136,
    10179 => 27138,
    10180 => 27140,
    10181 => 27141,
    10182 => 27143,
    10183 => 27145,
    10184 => 27147,
    10185 => 27148,
    10186 => 27150,
    10187 => 27152,
    10188 => 27154,
    10189 => 27155,
    10190 => 27157,
    10191 => 27159,
    10192 => 27161,
    10193 => 27162,
    10194 => 27164,
    10195 => 27166,
    10196 => 27168,
    10197 => 27169,
    10198 => 27171,
    10199 => 27173,
    10200 => 27175,
    10201 => 27177,
    10202 => 27178,
    10203 => 27180,
    10204 => 27182,
    10205 => 27184,
    10206 => 27185,
    10207 => 27187,
    10208 => 27189,
    10209 => 27191,
    10210 => 27192,
    10211 => 27194,
    10212 => 27196,
    10213 => 27198,
    10214 => 27199,
    10215 => 27201,
    10216 => 27203,
    10217 => 27205,
    10218 => 27206,
    10219 => 27208,
    10220 => 27210,
    10221 => 27212,
    10222 => 27213,
    10223 => 27215,
    10224 => 27217,
    10225 => 27219,
    10226 => 27220,
    10227 => 27222,
    10228 => 27224,
    10229 => 27226,
    10230 => 27227,
    10231 => 27229,
    10232 => 27231,
    10233 => 27233,
    10234 => 27234,
    10235 => 27236,
    10236 => 27238,
    10237 => 27240,
    10238 => 27241,
    10239 => 27243,
    10240 => 27245,
    10241 => 27247,
    10242 => 27248,
    10243 => 27250,
    10244 => 27252,
    10245 => 27253,
    10246 => 27255,
    10247 => 27257,
    10248 => 27259,
    10249 => 27260,
    10250 => 27262,
    10251 => 27264,
    10252 => 27266,
    10253 => 27267,
    10254 => 27269,
    10255 => 27271,
    10256 => 27273,
    10257 => 27274,
    10258 => 27276,
    10259 => 27278,
    10260 => 27280,
    10261 => 27281,
    10262 => 27283,
    10263 => 27285,
    10264 => 27287,
    10265 => 27288,
    10266 => 27290,
    10267 => 27292,
    10268 => 27294,
    10269 => 27295,
    10270 => 27297,
    10271 => 27299,
    10272 => 27300,
    10273 => 27302,
    10274 => 27304,
    10275 => 27306,
    10276 => 27307,
    10277 => 27309,
    10278 => 27311,
    10279 => 27313,
    10280 => 27314,
    10281 => 27316,
    10282 => 27318,
    10283 => 27320,
    10284 => 27321,
    10285 => 27323,
    10286 => 27325,
    10287 => 27327,
    10288 => 27328,
    10289 => 27330,
    10290 => 27332,
    10291 => 27333,
    10292 => 27335,
    10293 => 27337,
    10294 => 27339,
    10295 => 27340,
    10296 => 27342,
    10297 => 27344,
    10298 => 27346,
    10299 => 27347,
    10300 => 27349,
    10301 => 27351,
    10302 => 27352,
    10303 => 27354,
    10304 => 27356,
    10305 => 27358,
    10306 => 27359,
    10307 => 27361,
    10308 => 27363,
    10309 => 27365,
    10310 => 27366,
    10311 => 27368,
    10312 => 27370,
    10313 => 27372,
    10314 => 27373,
    10315 => 27375,
    10316 => 27377,
    10317 => 27378,
    10318 => 27380,
    10319 => 27382,
    10320 => 27384,
    10321 => 27385,
    10322 => 27387,
    10323 => 27389,
    10324 => 27390,
    10325 => 27392,
    10326 => 27394,
    10327 => 27396,
    10328 => 27397,
    10329 => 27399,
    10330 => 27401,
    10331 => 27403,
    10332 => 27404,
    10333 => 27406,
    10334 => 27408,
    10335 => 27409,
    10336 => 27411,
    10337 => 27413,
    10338 => 27415,
    10339 => 27416,
    10340 => 27418,
    10341 => 27420,
    10342 => 27421,
    10343 => 27423,
    10344 => 27425,
    10345 => 27427,
    10346 => 27428,
    10347 => 27430,
    10348 => 27432,
    10349 => 27434,
    10350 => 27435,
    10351 => 27437,
    10352 => 27439,
    10353 => 27440,
    10354 => 27442,
    10355 => 27444,
    10356 => 27446,
    10357 => 27447,
    10358 => 27449,
    10359 => 27451,
    10360 => 27452,
    10361 => 27454,
    10362 => 27456,
    10363 => 27458,
    10364 => 27459,
    10365 => 27461,
    10366 => 27463,
    10367 => 27464,
    10368 => 27466,
    10369 => 27468,
    10370 => 27470,
    10371 => 27471,
    10372 => 27473,
    10373 => 27475,
    10374 => 27476,
    10375 => 27478,
    10376 => 27480,
    10377 => 27482,
    10378 => 27483,
    10379 => 27485,
    10380 => 27487,
    10381 => 27488,
    10382 => 27490,
    10383 => 27492,
    10384 => 27493,
    10385 => 27495,
    10386 => 27497,
    10387 => 27499,
    10388 => 27500,
    10389 => 27502,
    10390 => 27504,
    10391 => 27505,
    10392 => 27507,
    10393 => 27509,
    10394 => 27511,
    10395 => 27512,
    10396 => 27514,
    10397 => 27516,
    10398 => 27517,
    10399 => 27519,
    10400 => 27521,
    10401 => 27523,
    10402 => 27524,
    10403 => 27526,
    10404 => 27528,
    10405 => 27529,
    10406 => 27531,
    10407 => 27533,
    10408 => 27534,
    10409 => 27536,
    10410 => 27538,
    10411 => 27540,
    10412 => 27541,
    10413 => 27543,
    10414 => 27545,
    10415 => 27546,
    10416 => 27548,
    10417 => 27550,
    10418 => 27551,
    10419 => 27553,
    10420 => 27555,
    10421 => 27557,
    10422 => 27558,
    10423 => 27560,
    10424 => 27562,
    10425 => 27563,
    10426 => 27565,
    10427 => 27567,
    10428 => 27568,
    10429 => 27570,
    10430 => 27572,
    10431 => 27574,
    10432 => 27575,
    10433 => 27577,
    10434 => 27579,
    10435 => 27580,
    10436 => 27582,
    10437 => 27584,
    10438 => 27585,
    10439 => 27587,
    10440 => 27589,
    10441 => 27590,
    10442 => 27592,
    10443 => 27594,
    10444 => 27596,
    10445 => 27597,
    10446 => 27599,
    10447 => 27601,
    10448 => 27602,
    10449 => 27604,
    10450 => 27606,
    10451 => 27607,
    10452 => 27609,
    10453 => 27611,
    10454 => 27613,
    10455 => 27614,
    10456 => 27616,
    10457 => 27618,
    10458 => 27619,
    10459 => 27621,
    10460 => 27623,
    10461 => 27624,
    10462 => 27626,
    10463 => 27628,
    10464 => 27629,
    10465 => 27631,
    10466 => 27633,
    10467 => 27634,
    10468 => 27636,
    10469 => 27638,
    10470 => 27640,
    10471 => 27641,
    10472 => 27643,
    10473 => 27645,
    10474 => 27646,
    10475 => 27648,
    10476 => 27650,
    10477 => 27651,
    10478 => 27653,
    10479 => 27655,
    10480 => 27656,
    10481 => 27658,
    10482 => 27660,
    10483 => 27661,
    10484 => 27663,
    10485 => 27665,
    10486 => 27666,
    10487 => 27668,
    10488 => 27670,
    10489 => 27672,
    10490 => 27673,
    10491 => 27675,
    10492 => 27677,
    10493 => 27678,
    10494 => 27680,
    10495 => 27682,
    10496 => 27683,
    10497 => 27685,
    10498 => 27687,
    10499 => 27688,
    10500 => 27690,
    10501 => 27692,
    10502 => 27693,
    10503 => 27695,
    10504 => 27697,
    10505 => 27698,
    10506 => 27700,
    10507 => 27702,
    10508 => 27703,
    10509 => 27705,
    10510 => 27707,
    10511 => 27708,
    10512 => 27710,
    10513 => 27712,
    10514 => 27714,
    10515 => 27715,
    10516 => 27717,
    10517 => 27719,
    10518 => 27720,
    10519 => 27722,
    10520 => 27724,
    10521 => 27725,
    10522 => 27727,
    10523 => 27729,
    10524 => 27730,
    10525 => 27732,
    10526 => 27734,
    10527 => 27735,
    10528 => 27737,
    10529 => 27739,
    10530 => 27740,
    10531 => 27742,
    10532 => 27744,
    10533 => 27745,
    10534 => 27747,
    10535 => 27749,
    10536 => 27750,
    10537 => 27752,
    10538 => 27754,
    10539 => 27755,
    10540 => 27757,
    10541 => 27759,
    10542 => 27760,
    10543 => 27762,
    10544 => 27764,
    10545 => 27765,
    10546 => 27767,
    10547 => 27769,
    10548 => 27770,
    10549 => 27772,
    10550 => 27774,
    10551 => 27775,
    10552 => 27777,
    10553 => 27779,
    10554 => 27780,
    10555 => 27782,
    10556 => 27784,
    10557 => 27785,
    10558 => 27787,
    10559 => 27789,
    10560 => 27790,
    10561 => 27792,
    10562 => 27794,
    10563 => 27795,
    10564 => 27797,
    10565 => 27799,
    10566 => 27800,
    10567 => 27802,
    10568 => 27804,
    10569 => 27805,
    10570 => 27807,
    10571 => 27809,
    10572 => 27810,
    10573 => 27812,
    10574 => 27814,
    10575 => 27815,
    10576 => 27817,
    10577 => 27819,
    10578 => 27820,
    10579 => 27822,
    10580 => 27824,
    10581 => 27825,
    10582 => 27827,
    10583 => 27829,
    10584 => 27830,
    10585 => 27832,
    10586 => 27834,
    10587 => 27835,
    10588 => 27837,
    10589 => 27839,
    10590 => 27840,
    10591 => 27842,
    10592 => 27843,
    10593 => 27845,
    10594 => 27847,
    10595 => 27848,
    10596 => 27850,
    10597 => 27852,
    10598 => 27853,
    10599 => 27855,
    10600 => 27857,
    10601 => 27858,
    10602 => 27860,
    10603 => 27862,
    10604 => 27863,
    10605 => 27865,
    10606 => 27867,
    10607 => 27868,
    10608 => 27870,
    10609 => 27872,
    10610 => 27873,
    10611 => 27875,
    10612 => 27877,
    10613 => 27878,
    10614 => 27880,
    10615 => 27882,
    10616 => 27883,
    10617 => 27885,
    10618 => 27886,
    10619 => 27888,
    10620 => 27890,
    10621 => 27891,
    10622 => 27893,
    10623 => 27895,
    10624 => 27896,
    10625 => 27898,
    10626 => 27900,
    10627 => 27901,
    10628 => 27903,
    10629 => 27905,
    10630 => 27906,
    10631 => 27908,
    10632 => 27910,
    10633 => 27911,
    10634 => 27913,
    10635 => 27914,
    10636 => 27916,
    10637 => 27918,
    10638 => 27919,
    10639 => 27921,
    10640 => 27923,
    10641 => 27924,
    10642 => 27926,
    10643 => 27928,
    10644 => 27929,
    10645 => 27931,
    10646 => 27933,
    10647 => 27934,
    10648 => 27936,
    10649 => 27937,
    10650 => 27939,
    10651 => 27941,
    10652 => 27942,
    10653 => 27944,
    10654 => 27946,
    10655 => 27947,
    10656 => 27949,
    10657 => 27951,
    10658 => 27952,
    10659 => 27954,
    10660 => 27956,
    10661 => 27957,
    10662 => 27959,
    10663 => 27960,
    10664 => 27962,
    10665 => 27964,
    10666 => 27965,
    10667 => 27967,
    10668 => 27969,
    10669 => 27970,
    10670 => 27972,
    10671 => 27974,
    10672 => 27975,
    10673 => 27977,
    10674 => 27978,
    10675 => 27980,
    10676 => 27982,
    10677 => 27983,
    10678 => 27985,
    10679 => 27987,
    10680 => 27988,
    10681 => 27990,
    10682 => 27992,
    10683 => 27993,
    10684 => 27995,
    10685 => 27996,
    10686 => 27998,
    10687 => 28000,
    10688 => 28001,
    10689 => 28003,
    10690 => 28005,
    10691 => 28006,
    10692 => 28008,
    10693 => 28009,
    10694 => 28011,
    10695 => 28013,
    10696 => 28014,
    10697 => 28016,
    10698 => 28018,
    10699 => 28019,
    10700 => 28021,
    10701 => 28022,
    10702 => 28024,
    10703 => 28026,
    10704 => 28027,
    10705 => 28029,
    10706 => 28031,
    10707 => 28032,
    10708 => 28034,
    10709 => 28036,
    10710 => 28037,
    10711 => 28039,
    10712 => 28040,
    10713 => 28042,
    10714 => 28044,
    10715 => 28045,
    10716 => 28047,
    10717 => 28049,
    10718 => 28050,
    10719 => 28052,
    10720 => 28053,
    10721 => 28055,
    10722 => 28057,
    10723 => 28058,
    10724 => 28060,
    10725 => 28061,
    10726 => 28063,
    10727 => 28065,
    10728 => 28066,
    10729 => 28068,
    10730 => 28070,
    10731 => 28071,
    10732 => 28073,
    10733 => 28074,
    10734 => 28076,
    10735 => 28078,
    10736 => 28079,
    10737 => 28081,
    10738 => 28083,
    10739 => 28084,
    10740 => 28086,
    10741 => 28087,
    10742 => 28089,
    10743 => 28091,
    10744 => 28092,
    10745 => 28094,
    10746 => 28095,
    10747 => 28097,
    10748 => 28099,
    10749 => 28100,
    10750 => 28102,
    10751 => 28104,
    10752 => 28105,
    10753 => 28107,
    10754 => 28108,
    10755 => 28110,
    10756 => 28112,
    10757 => 28113,
    10758 => 28115,
    10759 => 28116,
    10760 => 28118,
    10761 => 28120,
    10762 => 28121,
    10763 => 28123,
    10764 => 28125,
    10765 => 28126,
    10766 => 28128,
    10767 => 28129,
    10768 => 28131,
    10769 => 28133,
    10770 => 28134,
    10771 => 28136,
    10772 => 28137,
    10773 => 28139,
    10774 => 28141,
    10775 => 28142,
    10776 => 28144,
    10777 => 28145,
    10778 => 28147,
    10779 => 28149,
    10780 => 28150,
    10781 => 28152,
    10782 => 28154,
    10783 => 28155,
    10784 => 28157,
    10785 => 28158,
    10786 => 28160,
    10787 => 28162,
    10788 => 28163,
    10789 => 28165,
    10790 => 28166,
    10791 => 28168,
    10792 => 28170,
    10793 => 28171,
    10794 => 28173,
    10795 => 28174,
    10796 => 28176,
    10797 => 28178,
    10798 => 28179,
    10799 => 28181,
    10800 => 28182,
    10801 => 28184,
    10802 => 28186,
    10803 => 28187,
    10804 => 28189,
    10805 => 28190,
    10806 => 28192,
    10807 => 28194,
    10808 => 28195,
    10809 => 28197,
    10810 => 28198,
    10811 => 28200,
    10812 => 28202,
    10813 => 28203,
    10814 => 28205,
    10815 => 28206,
    10816 => 28208,
    10817 => 28210,
    10818 => 28211,
    10819 => 28213,
    10820 => 28214,
    10821 => 28216,
    10822 => 28218,
    10823 => 28219,
    10824 => 28221,
    10825 => 28222,
    10826 => 28224,
    10827 => 28226,
    10828 => 28227,
    10829 => 28229,
    10830 => 28230,
    10831 => 28232,
    10832 => 28234,
    10833 => 28235,
    10834 => 28237,
    10835 => 28238,
    10836 => 28240,
    10837 => 28242,
    10838 => 28243,
    10839 => 28245,
    10840 => 28246,
    10841 => 28248,
    10842 => 28249,
    10843 => 28251,
    10844 => 28253,
    10845 => 28254,
    10846 => 28256,
    10847 => 28257,
    10848 => 28259,
    10849 => 28261,
    10850 => 28262,
    10851 => 28264,
    10852 => 28265,
    10853 => 28267,
    10854 => 28269,
    10855 => 28270,
    10856 => 28272,
    10857 => 28273,
    10858 => 28275,
    10859 => 28277,
    10860 => 28278,
    10861 => 28280,
    10862 => 28281,
    10863 => 28283,
    10864 => 28284,
    10865 => 28286,
    10866 => 28288,
    10867 => 28289,
    10868 => 28291,
    10869 => 28292,
    10870 => 28294,
    10871 => 28296,
    10872 => 28297,
    10873 => 28299,
    10874 => 28300,
    10875 => 28302,
    10876 => 28303,
    10877 => 28305,
    10878 => 28307,
    10879 => 28308,
    10880 => 28310,
    10881 => 28311,
    10882 => 28313,
    10883 => 28315,
    10884 => 28316,
    10885 => 28318,
    10886 => 28319,
    10887 => 28321,
    10888 => 28322,
    10889 => 28324,
    10890 => 28326,
    10891 => 28327,
    10892 => 28329,
    10893 => 28330,
    10894 => 28332,
    10895 => 28333,
    10896 => 28335,
    10897 => 28337,
    10898 => 28338,
    10899 => 28340,
    10900 => 28341,
    10901 => 28343,
    10902 => 28345,
    10903 => 28346,
    10904 => 28348,
    10905 => 28349,
    10906 => 28351,
    10907 => 28352,
    10908 => 28354,
    10909 => 28356,
    10910 => 28357,
    10911 => 28359,
    10912 => 28360,
    10913 => 28362,
    10914 => 28363,
    10915 => 28365,
    10916 => 28367,
    10917 => 28368,
    10918 => 28370,
    10919 => 28371,
    10920 => 28373,
    10921 => 28374,
    10922 => 28376,
    10923 => 28378,
    10924 => 28379,
    10925 => 28381,
    10926 => 28382,
    10927 => 28384,
    10928 => 28385,
    10929 => 28387,
    10930 => 28389,
    10931 => 28390,
    10932 => 28392,
    10933 => 28393,
    10934 => 28395,
    10935 => 28396,
    10936 => 28398,
    10937 => 28400,
    10938 => 28401,
    10939 => 28403,
    10940 => 28404,
    10941 => 28406,
    10942 => 28407,
    10943 => 28409,
    10944 => 28411,
    10945 => 28412,
    10946 => 28414,
    10947 => 28415,
    10948 => 28417,
    10949 => 28418,
    10950 => 28420,
    10951 => 28421,
    10952 => 28423,
    10953 => 28425,
    10954 => 28426,
    10955 => 28428,
    10956 => 28429,
    10957 => 28431,
    10958 => 28432,
    10959 => 28434,
    10960 => 28436,
    10961 => 28437,
    10962 => 28439,
    10963 => 28440,
    10964 => 28442,
    10965 => 28443,
    10966 => 28445,
    10967 => 28446,
    10968 => 28448,
    10969 => 28450,
    10970 => 28451,
    10971 => 28453,
    10972 => 28454,
    10973 => 28456,
    10974 => 28457,
    10975 => 28459,
    10976 => 28460,
    10977 => 28462,
    10978 => 28464,
    10979 => 28465,
    10980 => 28467,
    10981 => 28468,
    10982 => 28470,
    10983 => 28471,
    10984 => 28473,
    10985 => 28474,
    10986 => 28476,
    10987 => 28478,
    10988 => 28479,
    10989 => 28481,
    10990 => 28482,
    10991 => 28484,
    10992 => 28485,
    10993 => 28487,
    10994 => 28488,
    10995 => 28490,
    10996 => 28492,
    10997 => 28493,
    10998 => 28495,
    10999 => 28496,
    11000 => 28498,
    11001 => 28499,
    11002 => 28501,
    11003 => 28502,
    11004 => 28504,
    11005 => 28505,
    11006 => 28507,
    11007 => 28509,
    11008 => 28510,
    11009 => 28512,
    11010 => 28513,
    11011 => 28515,
    11012 => 28516,
    11013 => 28518,
    11014 => 28519,
    11015 => 28521,
    11016 => 28523,
    11017 => 28524,
    11018 => 28526,
    11019 => 28527,
    11020 => 28529,
    11021 => 28530,
    11022 => 28532,
    11023 => 28533,
    11024 => 28535,
    11025 => 28536,
    11026 => 28538,
    11027 => 28540,
    11028 => 28541,
    11029 => 28543,
    11030 => 28544,
    11031 => 28546,
    11032 => 28547,
    11033 => 28549,
    11034 => 28550,
    11035 => 28552,
    11036 => 28553,
    11037 => 28555,
    11038 => 28556,
    11039 => 28558,
    11040 => 28560,
    11041 => 28561,
    11042 => 28563,
    11043 => 28564,
    11044 => 28566,
    11045 => 28567,
    11046 => 28569,
    11047 => 28570,
    11048 => 28572,
    11049 => 28573,
    11050 => 28575,
    11051 => 28576,
    11052 => 28578,
    11053 => 28580,
    11054 => 28581,
    11055 => 28583,
    11056 => 28584,
    11057 => 28586,
    11058 => 28587,
    11059 => 28589,
    11060 => 28590,
    11061 => 28592,
    11062 => 28593,
    11063 => 28595,
    11064 => 28596,
    11065 => 28598,
    11066 => 28600,
    11067 => 28601,
    11068 => 28603,
    11069 => 28604,
    11070 => 28606,
    11071 => 28607,
    11072 => 28609,
    11073 => 28610,
    11074 => 28612,
    11075 => 28613,
    11076 => 28615,
    11077 => 28616,
    11078 => 28618,
    11079 => 28619,
    11080 => 28621,
    11081 => 28622,
    11082 => 28624,
    11083 => 28626,
    11084 => 28627,
    11085 => 28629,
    11086 => 28630,
    11087 => 28632,
    11088 => 28633,
    11089 => 28635,
    11090 => 28636,
    11091 => 28638,
    11092 => 28639,
    11093 => 28641,
    11094 => 28642,
    11095 => 28644,
    11096 => 28645,
    11097 => 28647,
    11098 => 28648,
    11099 => 28650,
    11100 => 28651,
    11101 => 28653,
    11102 => 28655,
    11103 => 28656,
    11104 => 28658,
    11105 => 28659,
    11106 => 28661,
    11107 => 28662,
    11108 => 28664,
    11109 => 28665,
    11110 => 28667,
    11111 => 28668,
    11112 => 28670,
    11113 => 28671,
    11114 => 28673,
    11115 => 28674,
    11116 => 28676,
    11117 => 28677,
    11118 => 28679,
    11119 => 28680,
    11120 => 28682,
    11121 => 28683,
    11122 => 28685,
    11123 => 28686,
    11124 => 28688,
    11125 => 28690,
    11126 => 28691,
    11127 => 28693,
    11128 => 28694,
    11129 => 28696,
    11130 => 28697,
    11131 => 28699,
    11132 => 28700,
    11133 => 28702,
    11134 => 28703,
    11135 => 28705,
    11136 => 28706,
    11137 => 28708,
    11138 => 28709,
    11139 => 28711,
    11140 => 28712,
    11141 => 28714,
    11142 => 28715,
    11143 => 28717,
    11144 => 28718,
    11145 => 28720,
    11146 => 28721,
    11147 => 28723,
    11148 => 28724,
    11149 => 28726,
    11150 => 28727,
    11151 => 28729,
    11152 => 28730,
    11153 => 28732,
    11154 => 28733,
    11155 => 28735,
    11156 => 28736,
    11157 => 28738,
    11158 => 28739,
    11159 => 28741,
    11160 => 28742,
    11161 => 28744,
    11162 => 28745,
    11163 => 28747,
    11164 => 28748,
    11165 => 28750,
    11166 => 28752,
    11167 => 28753,
    11168 => 28755,
    11169 => 28756,
    11170 => 28758,
    11171 => 28759,
    11172 => 28761,
    11173 => 28762,
    11174 => 28764,
    11175 => 28765,
    11176 => 28767,
    11177 => 28768,
    11178 => 28770,
    11179 => 28771,
    11180 => 28773,
    11181 => 28774,
    11182 => 28776,
    11183 => 28777,
    11184 => 28779,
    11185 => 28780,
    11186 => 28782,
    11187 => 28783,
    11188 => 28785,
    11189 => 28786,
    11190 => 28788,
    11191 => 28789,
    11192 => 28791,
    11193 => 28792,
    11194 => 28794,
    11195 => 28795,
    11196 => 28797,
    11197 => 28798,
    11198 => 28800,
    11199 => 28801,
    11200 => 28803,
    11201 => 28804,
    11202 => 28806,
    11203 => 28807,
    11204 => 28809,
    11205 => 28810,
    11206 => 28812,
    11207 => 28813,
    11208 => 28815,
    11209 => 28816,
    11210 => 28818,
    11211 => 28819,
    11212 => 28821,
    11213 => 28822,
    11214 => 28824,
    11215 => 28825,
    11216 => 28827,
    11217 => 28828,
    11218 => 28830,
    11219 => 28831,
    11220 => 28832,
    11221 => 28834,
    11222 => 28835,
    11223 => 28837,
    11224 => 28838,
    11225 => 28840,
    11226 => 28841,
    11227 => 28843,
    11228 => 28844,
    11229 => 28846,
    11230 => 28847,
    11231 => 28849,
    11232 => 28850,
    11233 => 28852,
    11234 => 28853,
    11235 => 28855,
    11236 => 28856,
    11237 => 28858,
    11238 => 28859,
    11239 => 28861,
    11240 => 28862,
    11241 => 28864,
    11242 => 28865,
    11243 => 28867,
    11244 => 28868,
    11245 => 28870,
    11246 => 28871,
    11247 => 28873,
    11248 => 28874,
    11249 => 28876,
    11250 => 28877,
    11251 => 28879,
    11252 => 28880,
    11253 => 28882,
    11254 => 28883,
    11255 => 28885,
    11256 => 28886,
    11257 => 28888,
    11258 => 28889,
    11259 => 28891,
    11260 => 28892,
    11261 => 28893,
    11262 => 28895,
    11263 => 28896,
    11264 => 28898,
    11265 => 28899,
    11266 => 28901,
    11267 => 28902,
    11268 => 28904,
    11269 => 28905,
    11270 => 28907,
    11271 => 28908,
    11272 => 28910,
    11273 => 28911,
    11274 => 28913,
    11275 => 28914,
    11276 => 28916,
    11277 => 28917,
    11278 => 28919,
    11279 => 28920,
    11280 => 28922,
    11281 => 28923,
    11282 => 28925,
    11283 => 28926,
    11284 => 28927,
    11285 => 28929,
    11286 => 28930,
    11287 => 28932,
    11288 => 28933,
    11289 => 28935,
    11290 => 28936,
    11291 => 28938,
    11292 => 28939,
    11293 => 28941,
    11294 => 28942,
    11295 => 28944,
    11296 => 28945,
    11297 => 28947,
    11298 => 28948,
    11299 => 28950,
    11300 => 28951,
    11301 => 28953,
    11302 => 28954,
    11303 => 28955,
    11304 => 28957,
    11305 => 28958,
    11306 => 28960,
    11307 => 28961,
    11308 => 28963,
    11309 => 28964,
    11310 => 28966,
    11311 => 28967,
    11312 => 28969,
    11313 => 28970,
    11314 => 28972,
    11315 => 28973,
    11316 => 28975,
    11317 => 28976,
    11318 => 28977,
    11319 => 28979,
    11320 => 28980,
    11321 => 28982,
    11322 => 28983,
    11323 => 28985,
    11324 => 28986,
    11325 => 28988,
    11326 => 28989,
    11327 => 28991,
    11328 => 28992,
    11329 => 28994,
    11330 => 28995,
    11331 => 28997,
    11332 => 28998,
    11333 => 28999,
    11334 => 29001,
    11335 => 29002,
    11336 => 29004,
    11337 => 29005,
    11338 => 29007,
    11339 => 29008,
    11340 => 29010,
    11341 => 29011,
    11342 => 29013,
    11343 => 29014,
    11344 => 29016,
    11345 => 29017,
    11346 => 29018,
    11347 => 29020,
    11348 => 29021,
    11349 => 29023,
    11350 => 29024,
    11351 => 29026,
    11352 => 29027,
    11353 => 29029,
    11354 => 29030,
    11355 => 29032,
    11356 => 29033,
    11357 => 29034,
    11358 => 29036,
    11359 => 29037,
    11360 => 29039,
    11361 => 29040,
    11362 => 29042,
    11363 => 29043,
    11364 => 29045,
    11365 => 29046,
    11366 => 29048,
    11367 => 29049,
    11368 => 29050,
    11369 => 29052,
    11370 => 29053,
    11371 => 29055,
    11372 => 29056,
    11373 => 29058,
    11374 => 29059,
    11375 => 29061,
    11376 => 29062,
    11377 => 29064,
    11378 => 29065,
    11379 => 29066,
    11380 => 29068,
    11381 => 29069,
    11382 => 29071,
    11383 => 29072,
    11384 => 29074,
    11385 => 29075,
    11386 => 29077,
    11387 => 29078,
    11388 => 29079,
    11389 => 29081,
    11390 => 29082,
    11391 => 29084,
    11392 => 29085,
    11393 => 29087,
    11394 => 29088,
    11395 => 29090,
    11396 => 29091,
    11397 => 29093,
    11398 => 29094,
    11399 => 29095,
    11400 => 29097,
    11401 => 29098,
    11402 => 29100,
    11403 => 29101,
    11404 => 29103,
    11405 => 29104,
    11406 => 29106,
    11407 => 29107,
    11408 => 29108,
    11409 => 29110,
    11410 => 29111,
    11411 => 29113,
    11412 => 29114,
    11413 => 29116,
    11414 => 29117,
    11415 => 29118,
    11416 => 29120,
    11417 => 29121,
    11418 => 29123,
    11419 => 29124,
    11420 => 29126,
    11421 => 29127,
    11422 => 29129,
    11423 => 29130,
    11424 => 29131,
    11425 => 29133,
    11426 => 29134,
    11427 => 29136,
    11428 => 29137,
    11429 => 29139,
    11430 => 29140,
    11431 => 29142,
    11432 => 29143,
    11433 => 29144,
    11434 => 29146,
    11435 => 29147,
    11436 => 29149,
    11437 => 29150,
    11438 => 29152,
    11439 => 29153,
    11440 => 29154,
    11441 => 29156,
    11442 => 29157,
    11443 => 29159,
    11444 => 29160,
    11445 => 29162,
    11446 => 29163,
    11447 => 29164,
    11448 => 29166,
    11449 => 29167,
    11450 => 29169,
    11451 => 29170,
    11452 => 29172,
    11453 => 29173,
    11454 => 29174,
    11455 => 29176,
    11456 => 29177,
    11457 => 29179,
    11458 => 29180,
    11459 => 29182,
    11460 => 29183,
    11461 => 29184,
    11462 => 29186,
    11463 => 29187,
    11464 => 29189,
    11465 => 29190,
    11466 => 29192,
    11467 => 29193,
    11468 => 29194,
    11469 => 29196,
    11470 => 29197,
    11471 => 29199,
    11472 => 29200,
    11473 => 29202,
    11474 => 29203,
    11475 => 29204,
    11476 => 29206,
    11477 => 29207,
    11478 => 29209,
    11479 => 29210,
    11480 => 29212,
    11481 => 29213,
    11482 => 29214,
    11483 => 29216,
    11484 => 29217,
    11485 => 29219,
    11486 => 29220,
    11487 => 29222,
    11488 => 29223,
    11489 => 29224,
    11490 => 29226,
    11491 => 29227,
    11492 => 29229,
    11493 => 29230,
    11494 => 29231,
    11495 => 29233,
    11496 => 29234,
    11497 => 29236,
    11498 => 29237,
    11499 => 29239,
    11500 => 29240,
    11501 => 29241,
    11502 => 29243,
    11503 => 29244,
    11504 => 29246,
    11505 => 29247,
    11506 => 29248,
    11507 => 29250,
    11508 => 29251,
    11509 => 29253,
    11510 => 29254,
    11511 => 29256,
    11512 => 29257,
    11513 => 29258,
    11514 => 29260,
    11515 => 29261,
    11516 => 29263,
    11517 => 29264,
    11518 => 29265,
    11519 => 29267,
    11520 => 29268,
    11521 => 29270,
    11522 => 29271,
    11523 => 29273,
    11524 => 29274,
    11525 => 29275,
    11526 => 29277,
    11527 => 29278,
    11528 => 29280,
    11529 => 29281,
    11530 => 29282,
    11531 => 29284,
    11532 => 29285,
    11533 => 29287,
    11534 => 29288,
    11535 => 29289,
    11536 => 29291,
    11537 => 29292,
    11538 => 29294,
    11539 => 29295,
    11540 => 29296,
    11541 => 29298,
    11542 => 29299,
    11543 => 29301,
    11544 => 29302,
    11545 => 29304,
    11546 => 29305,
    11547 => 29306,
    11548 => 29308,
    11549 => 29309,
    11550 => 29311,
    11551 => 29312,
    11552 => 29313,
    11553 => 29315,
    11554 => 29316,
    11555 => 29318,
    11556 => 29319,
    11557 => 29320,
    11558 => 29322,
    11559 => 29323,
    11560 => 29325,
    11561 => 29326,
    11562 => 29327,
    11563 => 29329,
    11564 => 29330,
    11565 => 29332,
    11566 => 29333,
    11567 => 29334,
    11568 => 29336,
    11569 => 29337,
    11570 => 29339,
    11571 => 29340,
    11572 => 29341,
    11573 => 29343,
    11574 => 29344,
    11575 => 29346,
    11576 => 29347,
    11577 => 29348,
    11578 => 29350,
    11579 => 29351,
    11580 => 29353,
    11581 => 29354,
    11582 => 29355,
    11583 => 29357,
    11584 => 29358,
    11585 => 29360,
    11586 => 29361,
    11587 => 29362,
    11588 => 29364,
    11589 => 29365,
    11590 => 29366,
    11591 => 29368,
    11592 => 29369,
    11593 => 29371,
    11594 => 29372,
    11595 => 29373,
    11596 => 29375,
    11597 => 29376,
    11598 => 29378,
    11599 => 29379,
    11600 => 29380,
    11601 => 29382,
    11602 => 29383,
    11603 => 29385,
    11604 => 29386,
    11605 => 29387,
    11606 => 29389,
    11607 => 29390,
    11608 => 29392,
    11609 => 29393,
    11610 => 29394,
    11611 => 29396,
    11612 => 29397,
    11613 => 29398,
    11614 => 29400,
    11615 => 29401,
    11616 => 29403,
    11617 => 29404,
    11618 => 29405,
    11619 => 29407,
    11620 => 29408,
    11621 => 29410,
    11622 => 29411,
    11623 => 29412,
    11624 => 29414,
    11625 => 29415,
    11626 => 29416,
    11627 => 29418,
    11628 => 29419,
    11629 => 29421,
    11630 => 29422,
    11631 => 29423,
    11632 => 29425,
    11633 => 29426,
    11634 => 29428,
    11635 => 29429,
    11636 => 29430,
    11637 => 29432,
    11638 => 29433,
    11639 => 29434,
    11640 => 29436,
    11641 => 29437,
    11642 => 29439,
    11643 => 29440,
    11644 => 29441,
    11645 => 29443,
    11646 => 29444,
    11647 => 29445,
    11648 => 29447,
    11649 => 29448,
    11650 => 29450,
    11651 => 29451,
    11652 => 29452,
    11653 => 29454,
    11654 => 29455,
    11655 => 29457,
    11656 => 29458,
    11657 => 29459,
    11658 => 29461,
    11659 => 29462,
    11660 => 29463,
    11661 => 29465,
    11662 => 29466,
    11663 => 29468,
    11664 => 29469,
    11665 => 29470,
    11666 => 29472,
    11667 => 29473,
    11668 => 29474,
    11669 => 29476,
    11670 => 29477,
    11671 => 29478,
    11672 => 29480,
    11673 => 29481,
    11674 => 29483,
    11675 => 29484,
    11676 => 29485,
    11677 => 29487,
    11678 => 29488,
    11679 => 29489,
    11680 => 29491,
    11681 => 29492,
    11682 => 29494,
    11683 => 29495,
    11684 => 29496,
    11685 => 29498,
    11686 => 29499,
    11687 => 29500,
    11688 => 29502,
    11689 => 29503,
    11690 => 29504,
    11691 => 29506,
    11692 => 29507,
    11693 => 29509,
    11694 => 29510,
    11695 => 29511,
    11696 => 29513,
    11697 => 29514,
    11698 => 29515,
    11699 => 29517,
    11700 => 29518,
    11701 => 29520,
    11702 => 29521,
    11703 => 29522,
    11704 => 29524,
    11705 => 29525,
    11706 => 29526,
    11707 => 29528,
    11708 => 29529,
    11709 => 29530,
    11710 => 29532,
    11711 => 29533,
    11712 => 29534,
    11713 => 29536,
    11714 => 29537,
    11715 => 29539,
    11716 => 29540,
    11717 => 29541,
    11718 => 29543,
    11719 => 29544,
    11720 => 29545,
    11721 => 29547,
    11722 => 29548,
    11723 => 29549,
    11724 => 29551,
    11725 => 29552,
    11726 => 29554,
    11727 => 29555,
    11728 => 29556,
    11729 => 29558,
    11730 => 29559,
    11731 => 29560,
    11732 => 29562,
    11733 => 29563,
    11734 => 29564,
    11735 => 29566,
    11736 => 29567,
    11737 => 29568,
    11738 => 29570,
    11739 => 29571,
    11740 => 29572,
    11741 => 29574,
    11742 => 29575,
    11743 => 29577,
    11744 => 29578,
    11745 => 29579,
    11746 => 29581,
    11747 => 29582,
    11748 => 29583,
    11749 => 29585,
    11750 => 29586,
    11751 => 29587,
    11752 => 29589,
    11753 => 29590,
    11754 => 29591,
    11755 => 29593,
    11756 => 29594,
    11757 => 29595,
    11758 => 29597,
    11759 => 29598,
    11760 => 29599,
    11761 => 29601,
    11762 => 29602,
    11763 => 29604,
    11764 => 29605,
    11765 => 29606,
    11766 => 29608,
    11767 => 29609,
    11768 => 29610,
    11769 => 29612,
    11770 => 29613,
    11771 => 29614,
    11772 => 29616,
    11773 => 29617,
    11774 => 29618,
    11775 => 29620,
    11776 => 29621,
    11777 => 29622,
    11778 => 29624,
    11779 => 29625,
    11780 => 29626,
    11781 => 29628,
    11782 => 29629,
    11783 => 29630,
    11784 => 29632,
    11785 => 29633,
    11786 => 29634,
    11787 => 29636,
    11788 => 29637,
    11789 => 29638,
    11790 => 29640,
    11791 => 29641,
    11792 => 29642,
    11793 => 29644,
    11794 => 29645,
    11795 => 29646,
    11796 => 29648,
    11797 => 29649,
    11798 => 29651,
    11799 => 29652,
    11800 => 29653,
    11801 => 29655,
    11802 => 29656,
    11803 => 29657,
    11804 => 29659,
    11805 => 29660,
    11806 => 29661,
    11807 => 29663,
    11808 => 29664,
    11809 => 29665,
    11810 => 29667,
    11811 => 29668,
    11812 => 29669,
    11813 => 29671,
    11814 => 29672,
    11815 => 29673,
    11816 => 29675,
    11817 => 29676,
    11818 => 29677,
    11819 => 29679,
    11820 => 29680,
    11821 => 29681,
    11822 => 29683,
    11823 => 29684,
    11824 => 29685,
    11825 => 29687,
    11826 => 29688,
    11827 => 29689,
    11828 => 29690,
    11829 => 29692,
    11830 => 29693,
    11831 => 29694,
    11832 => 29696,
    11833 => 29697,
    11834 => 29698,
    11835 => 29700,
    11836 => 29701,
    11837 => 29702,
    11838 => 29704,
    11839 => 29705,
    11840 => 29706,
    11841 => 29708,
    11842 => 29709,
    11843 => 29710,
    11844 => 29712,
    11845 => 29713,
    11846 => 29714,
    11847 => 29716,
    11848 => 29717,
    11849 => 29718,
    11850 => 29720,
    11851 => 29721,
    11852 => 29722,
    11853 => 29724,
    11854 => 29725,
    11855 => 29726,
    11856 => 29728,
    11857 => 29729,
    11858 => 29730,
    11859 => 29732,
    11860 => 29733,
    11861 => 29734,
    11862 => 29736,
    11863 => 29737,
    11864 => 29738,
    11865 => 29739,
    11866 => 29741,
    11867 => 29742,
    11868 => 29743,
    11869 => 29745,
    11870 => 29746,
    11871 => 29747,
    11872 => 29749,
    11873 => 29750,
    11874 => 29751,
    11875 => 29753,
    11876 => 29754,
    11877 => 29755,
    11878 => 29757,
    11879 => 29758,
    11880 => 29759,
    11881 => 29761,
    11882 => 29762,
    11883 => 29763,
    11884 => 29764,
    11885 => 29766,
    11886 => 29767,
    11887 => 29768,
    11888 => 29770,
    11889 => 29771,
    11890 => 29772,
    11891 => 29774,
    11892 => 29775,
    11893 => 29776,
    11894 => 29778,
    11895 => 29779,
    11896 => 29780,
    11897 => 29782,
    11898 => 29783,
    11899 => 29784,
    11900 => 29785,
    11901 => 29787,
    11902 => 29788,
    11903 => 29789,
    11904 => 29791,
    11905 => 29792,
    11906 => 29793,
    11907 => 29795,
    11908 => 29796,
    11909 => 29797,
    11910 => 29799,
    11911 => 29800,
    11912 => 29801,
    11913 => 29802,
    11914 => 29804,
    11915 => 29805,
    11916 => 29806,
    11917 => 29808,
    11918 => 29809,
    11919 => 29810,
    11920 => 29812,
    11921 => 29813,
    11922 => 29814,
    11923 => 29816,
    11924 => 29817,
    11925 => 29818,
    11926 => 29819,
    11927 => 29821,
    11928 => 29822,
    11929 => 29823,
    11930 => 29825,
    11931 => 29826,
    11932 => 29827,
    11933 => 29829,
    11934 => 29830,
    11935 => 29831,
    11936 => 29832,
    11937 => 29834,
    11938 => 29835,
    11939 => 29836,
    11940 => 29838,
    11941 => 29839,
    11942 => 29840,
    11943 => 29842,
    11944 => 29843,
    11945 => 29844,
    11946 => 29845,
    11947 => 29847,
    11948 => 29848,
    11949 => 29849,
    11950 => 29851,
    11951 => 29852,
    11952 => 29853,
    11953 => 29854,
    11954 => 29856,
    11955 => 29857,
    11956 => 29858,
    11957 => 29860,
    11958 => 29861,
    11959 => 29862,
    11960 => 29864,
    11961 => 29865,
    11962 => 29866,
    11963 => 29867,
    11964 => 29869,
    11965 => 29870,
    11966 => 29871,
    11967 => 29873,
    11968 => 29874,
    11969 => 29875,
    11970 => 29876,
    11971 => 29878,
    11972 => 29879,
    11973 => 29880,
    11974 => 29882,
    11975 => 29883,
    11976 => 29884,
    11977 => 29885,
    11978 => 29887,
    11979 => 29888,
    11980 => 29889,
    11981 => 29891,
    11982 => 29892,
    11983 => 29893,
    11984 => 29894,
    11985 => 29896,
    11986 => 29897,
    11987 => 29898,
    11988 => 29900,
    11989 => 29901,
    11990 => 29902,
    11991 => 29903,
    11992 => 29905,
    11993 => 29906,
    11994 => 29907,
    11995 => 29909,
    11996 => 29910,
    11997 => 29911,
    11998 => 29912,
    11999 => 29914,
    12000 => 29915,
    12001 => 29916,
    12002 => 29918,
    12003 => 29919,
    12004 => 29920,
    12005 => 29921,
    12006 => 29923,
    12007 => 29924,
    12008 => 29925,
    12009 => 29927,
    12010 => 29928,
    12011 => 29929,
    12012 => 29930,
    12013 => 29932,
    12014 => 29933,
    12015 => 29934,
    12016 => 29936,
    12017 => 29937,
    12018 => 29938,
    12019 => 29939,
    12020 => 29941,
    12021 => 29942,
    12022 => 29943,
    12023 => 29944,
    12024 => 29946,
    12025 => 29947,
    12026 => 29948,
    12027 => 29950,
    12028 => 29951,
    12029 => 29952,
    12030 => 29953,
    12031 => 29955,
    12032 => 29956,
    12033 => 29957,
    12034 => 29958,
    12035 => 29960,
    12036 => 29961,
    12037 => 29962,
    12038 => 29964,
    12039 => 29965,
    12040 => 29966,
    12041 => 29967,
    12042 => 29969,
    12043 => 29970,
    12044 => 29971,
    12045 => 29972,
    12046 => 29974,
    12047 => 29975,
    12048 => 29976,
    12049 => 29978,
    12050 => 29979,
    12051 => 29980,
    12052 => 29981,
    12053 => 29983,
    12054 => 29984,
    12055 => 29985,
    12056 => 29986,
    12057 => 29988,
    12058 => 29989,
    12059 => 29990,
    12060 => 29991,
    12061 => 29993,
    12062 => 29994,
    12063 => 29995,
    12064 => 29997,
    12065 => 29998,
    12066 => 29999,
    12067 => 30000,
    12068 => 30002,
    12069 => 30003,
    12070 => 30004,
    12071 => 30005,
    12072 => 30007,
    12073 => 30008,
    12074 => 30009,
    12075 => 30010,
    12076 => 30012,
    12077 => 30013,
    12078 => 30014,
    12079 => 30015,
    12080 => 30017,
    12081 => 30018,
    12082 => 30019,
    12083 => 30020,
    12084 => 30022,
    12085 => 30023,
    12086 => 30024,
    12087 => 30026,
    12088 => 30027,
    12089 => 30028,
    12090 => 30029,
    12091 => 30031,
    12092 => 30032,
    12093 => 30033,
    12094 => 30034,
    12095 => 30036,
    12096 => 30037,
    12097 => 30038,
    12098 => 30039,
    12099 => 30041,
    12100 => 30042,
    12101 => 30043,
    12102 => 30044,
    12103 => 30046,
    12104 => 30047,
    12105 => 30048,
    12106 => 30049,
    12107 => 30051,
    12108 => 30052,
    12109 => 30053,
    12110 => 30054,
    12111 => 30056,
    12112 => 30057,
    12113 => 30058,
    12114 => 30059,
    12115 => 30061,
    12116 => 30062,
    12117 => 30063,
    12118 => 30064,
    12119 => 30066,
    12120 => 30067,
    12121 => 30068,
    12122 => 30069,
    12123 => 30071,
    12124 => 30072,
    12125 => 30073,
    12126 => 30074,
    12127 => 30076,
    12128 => 30077,
    12129 => 30078,
    12130 => 30079,
    12131 => 30081,
    12132 => 30082,
    12133 => 30083,
    12134 => 30084,
    12135 => 30086,
    12136 => 30087,
    12137 => 30088,
    12138 => 30089,
    12139 => 30091,
    12140 => 30092,
    12141 => 30093,
    12142 => 30094,
    12143 => 30096,
    12144 => 30097,
    12145 => 30098,
    12146 => 30099,
    12147 => 30100,
    12148 => 30102,
    12149 => 30103,
    12150 => 30104,
    12151 => 30105,
    12152 => 30107,
    12153 => 30108,
    12154 => 30109,
    12155 => 30110,
    12156 => 30112,
    12157 => 30113,
    12158 => 30114,
    12159 => 30115,
    12160 => 30117,
    12161 => 30118,
    12162 => 30119,
    12163 => 30120,
    12164 => 30122,
    12165 => 30123,
    12166 => 30124,
    12167 => 30125,
    12168 => 30126,
    12169 => 30128,
    12170 => 30129,
    12171 => 30130,
    12172 => 30131,
    12173 => 30133,
    12174 => 30134,
    12175 => 30135,
    12176 => 30136,
    12177 => 30138,
    12178 => 30139,
    12179 => 30140,
    12180 => 30141,
    12181 => 30143,
    12182 => 30144,
    12183 => 30145,
    12184 => 30146,
    12185 => 30147,
    12186 => 30149,
    12187 => 30150,
    12188 => 30151,
    12189 => 30152,
    12190 => 30154,
    12191 => 30155,
    12192 => 30156,
    12193 => 30157,
    12194 => 30159,
    12195 => 30160,
    12196 => 30161,
    12197 => 30162,
    12198 => 30163,
    12199 => 30165,
    12200 => 30166,
    12201 => 30167,
    12202 => 30168,
    12203 => 30170,
    12204 => 30171,
    12205 => 30172,
    12206 => 30173,
    12207 => 30174,
    12208 => 30176,
    12209 => 30177,
    12210 => 30178,
    12211 => 30179,
    12212 => 30181,
    12213 => 30182,
    12214 => 30183,
    12215 => 30184,
    12216 => 30185,
    12217 => 30187,
    12218 => 30188,
    12219 => 30189,
    12220 => 30190,
    12221 => 30192,
    12222 => 30193,
    12223 => 30194,
    12224 => 30195,
    12225 => 30196,
    12226 => 30198,
    12227 => 30199,
    12228 => 30200,
    12229 => 30201,
    12230 => 30203,
    12231 => 30204,
    12232 => 30205,
    12233 => 30206,
    12234 => 30207,
    12235 => 30209,
    12236 => 30210,
    12237 => 30211,
    12238 => 30212,
    12239 => 30214,
    12240 => 30215,
    12241 => 30216,
    12242 => 30217,
    12243 => 30218,
    12244 => 30220,
    12245 => 30221,
    12246 => 30222,
    12247 => 30223,
    12248 => 30224,
    12249 => 30226,
    12250 => 30227,
    12251 => 30228,
    12252 => 30229,
    12253 => 30231,
    12254 => 30232,
    12255 => 30233,
    12256 => 30234,
    12257 => 30235,
    12258 => 30237,
    12259 => 30238,
    12260 => 30239,
    12261 => 30240,
    12262 => 30241,
    12263 => 30243,
    12264 => 30244,
    12265 => 30245,
    12266 => 30246,
    12267 => 30247,
    12268 => 30249,
    12269 => 30250,
    12270 => 30251,
    12271 => 30252,
    12272 => 30253,
    12273 => 30255,
    12274 => 30256,
    12275 => 30257,
    12276 => 30258,
    12277 => 30260,
    12278 => 30261,
    12279 => 30262,
    12280 => 30263,
    12281 => 30264,
    12282 => 30266,
    12283 => 30267,
    12284 => 30268,
    12285 => 30269,
    12286 => 30270,
    12287 => 30272,
    12288 => 30273,
    12289 => 30274,
    12290 => 30275,
    12291 => 30276,
    12292 => 30278,
    12293 => 30279,
    12294 => 30280,
    12295 => 30281,
    12296 => 30282,
    12297 => 30284,
    12298 => 30285,
    12299 => 30286,
    12300 => 30287,
    12301 => 30288,
    12302 => 30290,
    12303 => 30291,
    12304 => 30292,
    12305 => 30293,
    12306 => 30294,
    12307 => 30296,
    12308 => 30297,
    12309 => 30298,
    12310 => 30299,
    12311 => 30300,
    12312 => 30302,
    12313 => 30303,
    12314 => 30304,
    12315 => 30305,
    12316 => 30306,
    12317 => 30308,
    12318 => 30309,
    12319 => 30310,
    12320 => 30311,
    12321 => 30312,
    12322 => 30313,
    12323 => 30315,
    12324 => 30316,
    12325 => 30317,
    12326 => 30318,
    12327 => 30319,
    12328 => 30321,
    12329 => 30322,
    12330 => 30323,
    12331 => 30324,
    12332 => 30325,
    12333 => 30327,
    12334 => 30328,
    12335 => 30329,
    12336 => 30330,
    12337 => 30331,
    12338 => 30333,
    12339 => 30334,
    12340 => 30335,
    12341 => 30336,
    12342 => 30337,
    12343 => 30338,
    12344 => 30340,
    12345 => 30341,
    12346 => 30342,
    12347 => 30343,
    12348 => 30344,
    12349 => 30346,
    12350 => 30347,
    12351 => 30348,
    12352 => 30349,
    12353 => 30350,
    12354 => 30351,
    12355 => 30353,
    12356 => 30354,
    12357 => 30355,
    12358 => 30356,
    12359 => 30357,
    12360 => 30359,
    12361 => 30360,
    12362 => 30361,
    12363 => 30362,
    12364 => 30363,
    12365 => 30365,
    12366 => 30366,
    12367 => 30367,
    12368 => 30368,
    12369 => 30369,
    12370 => 30370,
    12371 => 30372,
    12372 => 30373,
    12373 => 30374,
    12374 => 30375,
    12375 => 30376,
    12376 => 30377,
    12377 => 30379,
    12378 => 30380,
    12379 => 30381,
    12380 => 30382,
    12381 => 30383,
    12382 => 30385,
    12383 => 30386,
    12384 => 30387,
    12385 => 30388,
    12386 => 30389,
    12387 => 30390,
    12388 => 30392,
    12389 => 30393,
    12390 => 30394,
    12391 => 30395,
    12392 => 30396,
    12393 => 30397,
    12394 => 30399,
    12395 => 30400,
    12396 => 30401,
    12397 => 30402,
    12398 => 30403,
    12399 => 30404,
    12400 => 30406,
    12401 => 30407,
    12402 => 30408,
    12403 => 30409,
    12404 => 30410,
    12405 => 30412,
    12406 => 30413,
    12407 => 30414,
    12408 => 30415,
    12409 => 30416,
    12410 => 30417,
    12411 => 30419,
    12412 => 30420,
    12413 => 30421,
    12414 => 30422,
    12415 => 30423,
    12416 => 30424,
    12417 => 30426,
    12418 => 30427,
    12419 => 30428,
    12420 => 30429,
    12421 => 30430,
    12422 => 30431,
    12423 => 30433,
    12424 => 30434,
    12425 => 30435,
    12426 => 30436,
    12427 => 30437,
    12428 => 30438,
    12429 => 30439,
    12430 => 30441,
    12431 => 30442,
    12432 => 30443,
    12433 => 30444,
    12434 => 30445,
    12435 => 30446,
    12436 => 30448,
    12437 => 30449,
    12438 => 30450,
    12439 => 30451,
    12440 => 30452,
    12441 => 30453,
    12442 => 30455,
    12443 => 30456,
    12444 => 30457,
    12445 => 30458,
    12446 => 30459,
    12447 => 30460,
    12448 => 30462,
    12449 => 30463,
    12450 => 30464,
    12451 => 30465,
    12452 => 30466,
    12453 => 30467,
    12454 => 30468,
    12455 => 30470,
    12456 => 30471,
    12457 => 30472,
    12458 => 30473,
    12459 => 30474,
    12460 => 30475,
    12461 => 30477,
    12462 => 30478,
    12463 => 30479,
    12464 => 30480,
    12465 => 30481,
    12466 => 30482,
    12467 => 30483,
    12468 => 30485,
    12469 => 30486,
    12470 => 30487,
    12471 => 30488,
    12472 => 30489,
    12473 => 30490,
    12474 => 30492,
    12475 => 30493,
    12476 => 30494,
    12477 => 30495,
    12478 => 30496,
    12479 => 30497,
    12480 => 30498,
    12481 => 30500,
    12482 => 30501,
    12483 => 30502,
    12484 => 30503,
    12485 => 30504,
    12486 => 30505,
    12487 => 30506,
    12488 => 30508,
    12489 => 30509,
    12490 => 30510,
    12491 => 30511,
    12492 => 30512,
    12493 => 30513,
    12494 => 30514,
    12495 => 30516,
    12496 => 30517,
    12497 => 30518,
    12498 => 30519,
    12499 => 30520,
    12500 => 30521,
    12501 => 30522,
    12502 => 30524,
    12503 => 30525,
    12504 => 30526,
    12505 => 30527,
    12506 => 30528,
    12507 => 30529,
    12508 => 30530,
    12509 => 30532,
    12510 => 30533,
    12511 => 30534,
    12512 => 30535,
    12513 => 30536,
    12514 => 30537,
    12515 => 30538,
    12516 => 30540,
    12517 => 30541,
    12518 => 30542,
    12519 => 30543,
    12520 => 30544,
    12521 => 30545,
    12522 => 30546,
    12523 => 30548,
    12524 => 30549,
    12525 => 30550,
    12526 => 30551,
    12527 => 30552,
    12528 => 30553,
    12529 => 30554,
    12530 => 30556,
    12531 => 30557,
    12532 => 30558,
    12533 => 30559,
    12534 => 30560,
    12535 => 30561,
    12536 => 30562,
    12537 => 30563,
    12538 => 30565,
    12539 => 30566,
    12540 => 30567,
    12541 => 30568,
    12542 => 30569,
    12543 => 30570,
    12544 => 30571,
    12545 => 30573,
    12546 => 30574,
    12547 => 30575,
    12548 => 30576,
    12549 => 30577,
    12550 => 30578,
    12551 => 30579,
    12552 => 30580,
    12553 => 30582,
    12554 => 30583,
    12555 => 30584,
    12556 => 30585,
    12557 => 30586,
    12558 => 30587,
    12559 => 30588,
    12560 => 30589,
    12561 => 30591,
    12562 => 30592,
    12563 => 30593,
    12564 => 30594,
    12565 => 30595,
    12566 => 30596,
    12567 => 30597,
    12568 => 30598,
    12569 => 30600,
    12570 => 30601,
    12571 => 30602,
    12572 => 30603,
    12573 => 30604,
    12574 => 30605,
    12575 => 30606,
    12576 => 30607,
    12577 => 30609,
    12578 => 30610,
    12579 => 30611,
    12580 => 30612,
    12581 => 30613,
    12582 => 30614,
    12583 => 30615,
    12584 => 30616,
    12585 => 30617,
    12586 => 30619,
    12587 => 30620,
    12588 => 30621,
    12589 => 30622,
    12590 => 30623,
    12591 => 30624,
    12592 => 30625,
    12593 => 30626,
    12594 => 30628,
    12595 => 30629,
    12596 => 30630,
    12597 => 30631,
    12598 => 30632,
    12599 => 30633,
    12600 => 30634,
    12601 => 30635,
    12602 => 30636,
    12603 => 30638,
    12604 => 30639,
    12605 => 30640,
    12606 => 30641,
    12607 => 30642,
    12608 => 30643,
    12609 => 30644,
    12610 => 30645,
    12611 => 30646,
    12612 => 30648,
    12613 => 30649,
    12614 => 30650,
    12615 => 30651,
    12616 => 30652,
    12617 => 30653,
    12618 => 30654,
    12619 => 30655,
    12620 => 30656,
    12621 => 30658,
    12622 => 30659,
    12623 => 30660,
    12624 => 30661,
    12625 => 30662,
    12626 => 30663,
    12627 => 30664,
    12628 => 30665,
    12629 => 30666,
    12630 => 30668,
    12631 => 30669,
    12632 => 30670,
    12633 => 30671,
    12634 => 30672,
    12635 => 30673,
    12636 => 30674,
    12637 => 30675,
    12638 => 30676,
    12639 => 30678,
    12640 => 30679,
    12641 => 30680,
    12642 => 30681,
    12643 => 30682,
    12644 => 30683,
    12645 => 30684,
    12646 => 30685,
    12647 => 30686,
    12648 => 30687,
    12649 => 30689,
    12650 => 30690,
    12651 => 30691,
    12652 => 30692,
    12653 => 30693,
    12654 => 30694,
    12655 => 30695,
    12656 => 30696,
    12657 => 30697,
    12658 => 30698,
    12659 => 30700,
    12660 => 30701,
    12661 => 30702,
    12662 => 30703,
    12663 => 30704,
    12664 => 30705,
    12665 => 30706,
    12666 => 30707,
    12667 => 30708,
    12668 => 30709,
    12669 => 30711,
    12670 => 30712,
    12671 => 30713,
    12672 => 30714,
    12673 => 30715,
    12674 => 30716,
    12675 => 30717,
    12676 => 30718,
    12677 => 30719,
    12678 => 30720,
    12679 => 30721,
    12680 => 30723,
    12681 => 30724,
    12682 => 30725,
    12683 => 30726,
    12684 => 30727,
    12685 => 30728,
    12686 => 30729,
    12687 => 30730,
    12688 => 30731,
    12689 => 30732,
    12690 => 30733,
    12691 => 30735,
    12692 => 30736,
    12693 => 30737,
    12694 => 30738,
    12695 => 30739,
    12696 => 30740,
    12697 => 30741,
    12698 => 30742,
    12699 => 30743,
    12700 => 30744,
    12701 => 30745,
    12702 => 30746,
    12703 => 30748,
    12704 => 30749,
    12705 => 30750,
    12706 => 30751,
    12707 => 30752,
    12708 => 30753,
    12709 => 30754,
    12710 => 30755,
    12711 => 30756,
    12712 => 30757,
    12713 => 30758,
    12714 => 30760,
    12715 => 30761,
    12716 => 30762,
    12717 => 30763,
    12718 => 30764,
    12719 => 30765,
    12720 => 30766,
    12721 => 30767,
    12722 => 30768,
    12723 => 30769,
    12724 => 30770,
    12725 => 30771,
    12726 => 30772,
    12727 => 30774,
    12728 => 30775,
    12729 => 30776,
    12730 => 30777,
    12731 => 30778,
    12732 => 30779,
    12733 => 30780,
    12734 => 30781,
    12735 => 30782,
    12736 => 30783,
    12737 => 30784,
    12738 => 30785,
    12739 => 30786,
    12740 => 30788,
    12741 => 30789,
    12742 => 30790,
    12743 => 30791,
    12744 => 30792,
    12745 => 30793,
    12746 => 30794,
    12747 => 30795,
    12748 => 30796,
    12749 => 30797,
    12750 => 30798,
    12751 => 30799,
    12752 => 30800,
    12753 => 30802,
    12754 => 30803,
    12755 => 30804,
    12756 => 30805,
    12757 => 30806,
    12758 => 30807,
    12759 => 30808,
    12760 => 30809,
    12761 => 30810,
    12762 => 30811,
    12763 => 30812,
    12764 => 30813,
    12765 => 30814,
    12766 => 30815,
    12767 => 30816,
    12768 => 30818,
    12769 => 30819,
    12770 => 30820,
    12771 => 30821,
    12772 => 30822,
    12773 => 30823,
    12774 => 30824,
    12775 => 30825,
    12776 => 30826,
    12777 => 30827,
    12778 => 30828,
    12779 => 30829,
    12780 => 30830,
    12781 => 30831,
    12782 => 30832,
    12783 => 30834,
    12784 => 30835,
    12785 => 30836,
    12786 => 30837,
    12787 => 30838,
    12788 => 30839,
    12789 => 30840,
    12790 => 30841,
    12791 => 30842,
    12792 => 30843,
    12793 => 30844,
    12794 => 30845,
    12795 => 30846,
    12796 => 30847,
    12797 => 30848,
    12798 => 30849,
    12799 => 30851,
    12800 => 30852,
    12801 => 30853,
    12802 => 30854,
    12803 => 30855,
    12804 => 30856,
    12805 => 30857,
    12806 => 30858,
    12807 => 30859,
    12808 => 30860,
    12809 => 30861,
    12810 => 30862,
    12811 => 30863,
    12812 => 30864,
    12813 => 30865,
    12814 => 30866,
    12815 => 30867,
    12816 => 30868,
    12817 => 30870,
    12818 => 30871,
    12819 => 30872,
    12820 => 30873,
    12821 => 30874,
    12822 => 30875,
    12823 => 30876,
    12824 => 30877,
    12825 => 30878,
    12826 => 30879,
    12827 => 30880,
    12828 => 30881,
    12829 => 30882,
    12830 => 30883,
    12831 => 30884,
    12832 => 30885,
    12833 => 30886,
    12834 => 30887,
    12835 => 30888,
    12836 => 30889,
    12837 => 30891,
    12838 => 30892,
    12839 => 30893,
    12840 => 30894,
    12841 => 30895,
    12842 => 30896,
    12843 => 30897,
    12844 => 30898,
    12845 => 30899,
    12846 => 30900,
    12847 => 30901,
    12848 => 30902,
    12849 => 30903,
    12850 => 30904,
    12851 => 30905,
    12852 => 30906,
    12853 => 30907,
    12854 => 30908,
    12855 => 30909,
    12856 => 30910,
    12857 => 30911,
    12858 => 30912,
    12859 => 30914,
    12860 => 30915,
    12861 => 30916,
    12862 => 30917,
    12863 => 30918,
    12864 => 30919,
    12865 => 30920,
    12866 => 30921,
    12867 => 30922,
    12868 => 30923,
    12869 => 30924,
    12870 => 30925,
    12871 => 30926,
    12872 => 30927,
    12873 => 30928,
    12874 => 30929,
    12875 => 30930,
    12876 => 30931,
    12877 => 30932,
    12878 => 30933,
    12879 => 30934,
    12880 => 30935,
    12881 => 30936,
    12882 => 30937,
    12883 => 30938,
    12884 => 30939,
    12885 => 30941,
    12886 => 30942,
    12887 => 30943,
    12888 => 30944,
    12889 => 30945,
    12890 => 30946,
    12891 => 30947,
    12892 => 30948,
    12893 => 30949,
    12894 => 30950,
    12895 => 30951,
    12896 => 30952,
    12897 => 30953,
    12898 => 30954,
    12899 => 30955,
    12900 => 30956,
    12901 => 30957,
    12902 => 30958,
    12903 => 30959,
    12904 => 30960,
    12905 => 30961,
    12906 => 30962,
    12907 => 30963,
    12908 => 30964,
    12909 => 30965,
    12910 => 30966,
    12911 => 30967,
    12912 => 30968,
    12913 => 30969,
    12914 => 30970,
    12915 => 30971,
    12916 => 30972,
    12917 => 30973,
    12918 => 30974,
    12919 => 30976,
    12920 => 30977,
    12921 => 30978,
    12922 => 30979,
    12923 => 30980,
    12924 => 30981,
    12925 => 30982,
    12926 => 30983,
    12927 => 30984,
    12928 => 30985,
    12929 => 30986,
    12930 => 30987,
    12931 => 30988,
    12932 => 30989,
    12933 => 30990,
    12934 => 30991,
    12935 => 30992,
    12936 => 30993,
    12937 => 30994,
    12938 => 30995,
    12939 => 30996,
    12940 => 30997,
    12941 => 30998,
    12942 => 30999,
    12943 => 31000,
    12944 => 31001,
    12945 => 31002,
    12946 => 31003,
    12947 => 31004,
    12948 => 31005,
    12949 => 31006,
    12950 => 31007,
    12951 => 31008,
    12952 => 31009,
    12953 => 31010,
    12954 => 31011,
    12955 => 31012,
    12956 => 31013,
    12957 => 31014,
    12958 => 31015,
    12959 => 31016,
    12960 => 31017,
    12961 => 31018,
    12962 => 31019,
    12963 => 31020,
    12964 => 31021,
    12965 => 31022,
    12966 => 31023,
    12967 => 31024,
    12968 => 31025,
    12969 => 31026,
    12970 => 31027,
    12971 => 31028,
    12972 => 31029,
    12973 => 31030,
    12974 => 31031,
    12975 => 31032,
    12976 => 31033,
    12977 => 31034,
    12978 => 31035,
    12979 => 31036,
    12980 => 31037,
    12981 => 31038,
    12982 => 31039,
    12983 => 31040,
    12984 => 31041,
    12985 => 31043,
    12986 => 31044,
    12987 => 31045,
    12988 => 31046,
    12989 => 31047,
    12990 => 31048,
    12991 => 31049,
    12992 => 31050,
    12993 => 31051,
    12994 => 31052,
    12995 => 31053,
    12996 => 31054,
    12997 => 31055,
    12998 => 31056,
    12999 => 31057,
    13000 => 31058,
    13001 => 31059,
    13002 => 31060,
    13003 => 31061,
    13004 => 31062,
    13005 => 31063,
    13006 => 31064,
    13007 => 31065,
    13008 => 31066,
    13009 => 31067,
    13010 => 31068,
    13011 => 31069,
    13012 => 31070,
    13013 => 31071,
    13014 => 31072,
    13015 => 31073,
    13016 => 31074,
    13017 => 31075,
    13018 => 31076,
    13019 => 31077,
    13020 => 31078,
    13021 => 31079,
    13022 => 31080,
    13023 => 31081,
    13024 => 31082,
    13025 => 31083,
    13026 => 31083,
    13027 => 31084,
    13028 => 31085,
    13029 => 31086,
    13030 => 31087,
    13031 => 31088,
    13032 => 31089,
    13033 => 31090,
    13034 => 31091,
    13035 => 31092,
    13036 => 31093,
    13037 => 31094,
    13038 => 31095,
    13039 => 31096,
    13040 => 31097,
    13041 => 31098,
    13042 => 31099,
    13043 => 31100,
    13044 => 31101,
    13045 => 31102,
    13046 => 31103,
    13047 => 31104,
    13048 => 31105,
    13049 => 31106,
    13050 => 31107,
    13051 => 31108,
    13052 => 31109,
    13053 => 31110,
    13054 => 31111,
    13055 => 31112,
    13056 => 31113,
    13057 => 31114,
    13058 => 31115,
    13059 => 31116,
    13060 => 31117,
    13061 => 31118,
    13062 => 31119,
    13063 => 31120,
    13064 => 31121,
    13065 => 31122,
    13066 => 31123,
    13067 => 31124,
    13068 => 31125,
    13069 => 31126,
    13070 => 31127,
    13071 => 31128,
    13072 => 31129,
    13073 => 31130,
    13074 => 31131,
    13075 => 31132,
    13076 => 31133,
    13077 => 31134,
    13078 => 31135,
    13079 => 31136,
    13080 => 31137,
    13081 => 31138,
    13082 => 31139,
    13083 => 31140,
    13084 => 31141,
    13085 => 31142,
    13086 => 31143,
    13087 => 31144,
    13088 => 31145,
    13089 => 31146,
    13090 => 31147,
    13091 => 31148,
    13092 => 31148,
    13093 => 31149,
    13094 => 31150,
    13095 => 31151,
    13096 => 31152,
    13097 => 31153,
    13098 => 31154,
    13099 => 31155,
    13100 => 31156,
    13101 => 31157,
    13102 => 31158,
    13103 => 31159,
    13104 => 31160,
    13105 => 31161,
    13106 => 31162,
    13107 => 31163,
    13108 => 31164,
    13109 => 31165,
    13110 => 31166,
    13111 => 31167,
    13112 => 31168,
    13113 => 31169,
    13114 => 31170,
    13115 => 31171,
    13116 => 31172,
    13117 => 31173,
    13118 => 31174,
    13119 => 31175,
    13120 => 31176,
    13121 => 31177,
    13122 => 31178,
    13123 => 31179,
    13124 => 31180,
    13125 => 31181,
    13126 => 31181,
    13127 => 31182,
    13128 => 31183,
    13129 => 31184,
    13130 => 31185,
    13131 => 31186,
    13132 => 31187,
    13133 => 31188,
    13134 => 31189,
    13135 => 31190,
    13136 => 31191,
    13137 => 31192,
    13138 => 31193,
    13139 => 31194,
    13140 => 31195,
    13141 => 31196,
    13142 => 31197,
    13143 => 31198,
    13144 => 31199,
    13145 => 31200,
    13146 => 31201,
    13147 => 31202,
    13148 => 31203,
    13149 => 31204,
    13150 => 31205,
    13151 => 31206,
    13152 => 31206,
    13153 => 31207,
    13154 => 31208,
    13155 => 31209,
    13156 => 31210,
    13157 => 31211,
    13158 => 31212,
    13159 => 31213,
    13160 => 31214,
    13161 => 31215,
    13162 => 31216,
    13163 => 31217,
    13164 => 31218,
    13165 => 31219,
    13166 => 31220,
    13167 => 31221,
    13168 => 31222,
    13169 => 31223,
    13170 => 31224,
    13171 => 31225,
    13172 => 31226,
    13173 => 31227,
    13174 => 31227,
    13175 => 31228,
    13176 => 31229,
    13177 => 31230,
    13178 => 31231,
    13179 => 31232,
    13180 => 31233,
    13181 => 31234,
    13182 => 31235,
    13183 => 31236,
    13184 => 31237,
    13185 => 31238,
    13186 => 31239,
    13187 => 31240,
    13188 => 31241,
    13189 => 31242,
    13190 => 31243,
    13191 => 31244,
    13192 => 31245,
    13193 => 31246,
    13194 => 31246,
    13195 => 31247,
    13196 => 31248,
    13197 => 31249,
    13198 => 31250,
    13199 => 31251,
    13200 => 31252,
    13201 => 31253,
    13202 => 31254,
    13203 => 31255,
    13204 => 31256,
    13205 => 31257,
    13206 => 31258,
    13207 => 31259,
    13208 => 31260,
    13209 => 31261,
    13210 => 31262,
    13211 => 31262,
    13212 => 31263,
    13213 => 31264,
    13214 => 31265,
    13215 => 31266,
    13216 => 31267,
    13217 => 31268,
    13218 => 31269,
    13219 => 31270,
    13220 => 31271,
    13221 => 31272,
    13222 => 31273,
    13223 => 31274,
    13224 => 31275,
    13225 => 31276,
    13226 => 31277,
    13227 => 31278,
    13228 => 31278,
    13229 => 31279,
    13230 => 31280,
    13231 => 31281,
    13232 => 31282,
    13233 => 31283,
    13234 => 31284,
    13235 => 31285,
    13236 => 31286,
    13237 => 31287,
    13238 => 31288,
    13239 => 31289,
    13240 => 31290,
    13241 => 31291,
    13242 => 31292,
    13243 => 31292,
    13244 => 31293,
    13245 => 31294,
    13246 => 31295,
    13247 => 31296,
    13248 => 31297,
    13249 => 31298,
    13250 => 31299,
    13251 => 31300,
    13252 => 31301,
    13253 => 31302,
    13254 => 31303,
    13255 => 31304,
    13256 => 31305,
    13257 => 31305,
    13258 => 31306,
    13259 => 31307,
    13260 => 31308,
    13261 => 31309,
    13262 => 31310,
    13263 => 31311,
    13264 => 31312,
    13265 => 31313,
    13266 => 31314,
    13267 => 31315,
    13268 => 31316,
    13269 => 31317,
    13270 => 31318,
    13271 => 31318,
    13272 => 31319,
    13273 => 31320,
    13274 => 31321,
    13275 => 31322,
    13276 => 31323,
    13277 => 31324,
    13278 => 31325,
    13279 => 31326,
    13280 => 31327,
    13281 => 31328,
    13282 => 31329,
    13283 => 31329,
    13284 => 31330,
    13285 => 31331,
    13286 => 31332,
    13287 => 31333,
    13288 => 31334,
    13289 => 31335,
    13290 => 31336,
    13291 => 31337,
    13292 => 31338,
    13293 => 31339,
    13294 => 31340,
    13295 => 31341,
    13296 => 31341,
    13297 => 31342,
    13298 => 31343,
    13299 => 31344,
    13300 => 31345,
    13301 => 31346,
    13302 => 31347,
    13303 => 31348,
    13304 => 31349,
    13305 => 31350,
    13306 => 31351,
    13307 => 31352,
    13308 => 31352,
    13309 => 31353,
    13310 => 31354,
    13311 => 31355,
    13312 => 31356,
    13313 => 31357,
    13314 => 31358,
    13315 => 31359,
    13316 => 31360,
    13317 => 31361,
    13318 => 31362,
    13319 => 31362,
    13320 => 31363,
    13321 => 31364,
    13322 => 31365,
    13323 => 31366,
    13324 => 31367,
    13325 => 31368,
    13326 => 31369,
    13327 => 31370,
    13328 => 31371,
    13329 => 31372,
    13330 => 31372,
    13331 => 31373,
    13332 => 31374,
    13333 => 31375,
    13334 => 31376,
    13335 => 31377,
    13336 => 31378,
    13337 => 31379,
    13338 => 31380,
    13339 => 31381,
    13340 => 31381,
    13341 => 31382,
    13342 => 31383,
    13343 => 31384,
    13344 => 31385,
    13345 => 31386,
    13346 => 31387,
    13347 => 31388,
    13348 => 31389,
    13349 => 31390,
    13350 => 31391,
    13351 => 31391,
    13352 => 31392,
    13353 => 31393,
    13354 => 31394,
    13355 => 31395,
    13356 => 31396,
    13357 => 31397,
    13358 => 31398,
    13359 => 31399,
    13360 => 31400,
    13361 => 31400,
    13362 => 31401,
    13363 => 31402,
    13364 => 31403,
    13365 => 31404,
    13366 => 31405,
    13367 => 31406,
    13368 => 31407,
    13369 => 31408,
    13370 => 31408,
    13371 => 31409,
    13372 => 31410,
    13373 => 31411,
    13374 => 31412,
    13375 => 31413,
    13376 => 31414,
    13377 => 31415,
    13378 => 31416,
    13379 => 31417,
    13380 => 31417,
    13381 => 31418,
    13382 => 31419,
    13383 => 31420,
    13384 => 31421,
    13385 => 31422,
    13386 => 31423,
    13387 => 31424,
    13388 => 31425,
    13389 => 31425,
    13390 => 31426,
    13391 => 31427,
    13392 => 31428,
    13393 => 31429,
    13394 => 31430,
    13395 => 31431,
    13396 => 31432,
    13397 => 31433,
    13398 => 31433,
    13399 => 31434,
    13400 => 31435,
    13401 => 31436,
    13402 => 31437,
    13403 => 31438,
    13404 => 31439,
    13405 => 31440,
    13406 => 31441,
    13407 => 31441,
    13408 => 31442,
    13409 => 31443,
    13410 => 31444,
    13411 => 31445,
    13412 => 31446,
    13413 => 31447,
    13414 => 31448,
    13415 => 31448,
    13416 => 31449,
    13417 => 31450,
    13418 => 31451,
    13419 => 31452,
    13420 => 31453,
    13421 => 31454,
    13422 => 31455,
    13423 => 31456,
    13424 => 31456,
    13425 => 31457,
    13426 => 31458,
    13427 => 31459,
    13428 => 31460,
    13429 => 31461,
    13430 => 31462,
    13431 => 31463,
    13432 => 31463,
    13433 => 31464,
    13434 => 31465,
    13435 => 31466,
    13436 => 31467,
    13437 => 31468,
    13438 => 31469,
    13439 => 31470,
    13440 => 31470,
    13441 => 31471,
    13442 => 31472,
    13443 => 31473,
    13444 => 31474,
    13445 => 31475,
    13446 => 31476,
    13447 => 31477,
    13448 => 31477,
    13449 => 31478,
    13450 => 31479,
    13451 => 31480,
    13452 => 31481,
    13453 => 31482,
    13454 => 31483,
    13455 => 31484,
    13456 => 31484,
    13457 => 31485,
    13458 => 31486,
    13459 => 31487,
    13460 => 31488,
    13461 => 31489,
    13462 => 31490,
    13463 => 31490,
    13464 => 31491,
    13465 => 31492,
    13466 => 31493,
    13467 => 31494,
    13468 => 31495,
    13469 => 31496,
    13470 => 31497,
    13471 => 31497,
    13472 => 31498,
    13473 => 31499,
    13474 => 31500,
    13475 => 31501,
    13476 => 31502,
    13477 => 31503,
    13478 => 31503,
    13479 => 31504,
    13480 => 31505,
    13481 => 31506,
    13482 => 31507,
    13483 => 31508,
    13484 => 31509,
    13485 => 31510,
    13486 => 31510,
    13487 => 31511,
    13488 => 31512,
    13489 => 31513,
    13490 => 31514,
    13491 => 31515,
    13492 => 31516,
    13493 => 31516,
    13494 => 31517,
    13495 => 31518,
    13496 => 31519,
    13497 => 31520,
    13498 => 31521,
    13499 => 31522,
    13500 => 31522,
    13501 => 31523,
    13502 => 31524,
    13503 => 31525,
    13504 => 31526,
    13505 => 31527,
    13506 => 31528,
    13507 => 31528,
    13508 => 31529,
    13509 => 31530,
    13510 => 31531,
    13511 => 31532,
    13512 => 31533,
    13513 => 31534,
    13514 => 31534,
    13515 => 31535,
    13516 => 31536,
    13517 => 31537,
    13518 => 31538,
    13519 => 31539,
    13520 => 31539,
    13521 => 31540,
    13522 => 31541,
    13523 => 31542,
    13524 => 31543,
    13525 => 31544,
    13526 => 31545,
    13527 => 31545,
    13528 => 31546,
    13529 => 31547,
    13530 => 31548,
    13531 => 31549,
    13532 => 31550,
    13533 => 31551,
    13534 => 31551,
    13535 => 31552,
    13536 => 31553,
    13537 => 31554,
    13538 => 31555,
    13539 => 31556,
    13540 => 31556,
    13541 => 31557,
    13542 => 31558,
    13543 => 31559,
    13544 => 31560,
    13545 => 31561,
    13546 => 31562,
    13547 => 31562,
    13548 => 31563,
    13549 => 31564,
    13550 => 31565,
    13551 => 31566,
    13552 => 31567,
    13553 => 31567,
    13554 => 31568,
    13555 => 31569,
    13556 => 31570,
    13557 => 31571,
    13558 => 31572,
    13559 => 31572,
    13560 => 31573,
    13561 => 31574,
    13562 => 31575,
    13563 => 31576,
    13564 => 31577,
    13565 => 31578,
    13566 => 31578,
    13567 => 31579,
    13568 => 31580,
    13569 => 31581,
    13570 => 31582,
    13571 => 31583,
    13572 => 31583,
    13573 => 31584,
    13574 => 31585,
    13575 => 31586,
    13576 => 31587,
    13577 => 31588,
    13578 => 31588,
    13579 => 31589,
    13580 => 31590,
    13581 => 31591,
    13582 => 31592,
    13583 => 31593,
    13584 => 31593,
    13585 => 31594,
    13586 => 31595,
    13587 => 31596,
    13588 => 31597,
    13589 => 31598,
    13590 => 31598,
    13591 => 31599,
    13592 => 31600,
    13593 => 31601,
    13594 => 31602,
    13595 => 31603,
    13596 => 31603,
    13597 => 31604,
    13598 => 31605,
    13599 => 31606,
    13600 => 31607,
    13601 => 31608,
    13602 => 31608,
    13603 => 31609,
    13604 => 31610,
    13605 => 31611,
    13606 => 31612,
    13607 => 31613,
    13608 => 31613,
    13609 => 31614,
    13610 => 31615,
    13611 => 31616,
    13612 => 31617,
    13613 => 31617,
    13614 => 31618,
    13615 => 31619,
    13616 => 31620,
    13617 => 31621,
    13618 => 31622,
    13619 => 31622,
    13620 => 31623,
    13621 => 31624,
    13622 => 31625,
    13623 => 31626,
    13624 => 31627,
    13625 => 31627,
    13626 => 31628,
    13627 => 31629,
    13628 => 31630,
    13629 => 31631,
    13630 => 31631,
    13631 => 31632,
    13632 => 31633,
    13633 => 31634,
    13634 => 31635,
    13635 => 31636,
    13636 => 31636,
    13637 => 31637,
    13638 => 31638,
    13639 => 31639,
    13640 => 31640,
    13641 => 31640,
    13642 => 31641,
    13643 => 31642,
    13644 => 31643,
    13645 => 31644,
    13646 => 31645,
    13647 => 31645,
    13648 => 31646,
    13649 => 31647,
    13650 => 31648,
    13651 => 31649,
    13652 => 31649,
    13653 => 31650,
    13654 => 31651,
    13655 => 31652,
    13656 => 31653,
    13657 => 31653,
    13658 => 31654,
    13659 => 31655,
    13660 => 31656,
    13661 => 31657,
    13662 => 31658,
    13663 => 31658,
    13664 => 31659,
    13665 => 31660,
    13666 => 31661,
    13667 => 31662,
    13668 => 31662,
    13669 => 31663,
    13670 => 31664,
    13671 => 31665,
    13672 => 31666,
    13673 => 31666,
    13674 => 31667,
    13675 => 31668,
    13676 => 31669,
    13677 => 31670,
    13678 => 31670,
    13679 => 31671,
    13680 => 31672,
    13681 => 31673,
    13682 => 31674,
    13683 => 31674,
    13684 => 31675,
    13685 => 31676,
    13686 => 31677,
    13687 => 31678,
    13688 => 31679,
    13689 => 31679,
    13690 => 31680,
    13691 => 31681,
    13692 => 31682,
    13693 => 31683,
    13694 => 31683,
    13695 => 31684,
    13696 => 31685,
    13697 => 31686,
    13698 => 31687,
    13699 => 31687,
    13700 => 31688,
    13701 => 31689,
    13702 => 31690,
    13703 => 31691,
    13704 => 31691,
    13705 => 31692,
    13706 => 31693,
    13707 => 31694,
    13708 => 31695,
    13709 => 31695,
    13710 => 31696,
    13711 => 31697,
    13712 => 31698,
    13713 => 31698,
    13714 => 31699,
    13715 => 31700,
    13716 => 31701,
    13717 => 31702,
    13718 => 31702,
    13719 => 31703,
    13720 => 31704,
    13721 => 31705,
    13722 => 31706,
    13723 => 31706,
    13724 => 31707,
    13725 => 31708,
    13726 => 31709,
    13727 => 31710,
    13728 => 31710,
    13729 => 31711,
    13730 => 31712,
    13731 => 31713,
    13732 => 31714,
    13733 => 31714,
    13734 => 31715,
    13735 => 31716,
    13736 => 31717,
    13737 => 31718,
    13738 => 31718,
    13739 => 31719,
    13740 => 31720,
    13741 => 31721,
    13742 => 31721,
    13743 => 31722,
    13744 => 31723,
    13745 => 31724,
    13746 => 31725,
    13747 => 31725,
    13748 => 31726,
    13749 => 31727,
    13750 => 31728,
    13751 => 31729,
    13752 => 31729,
    13753 => 31730,
    13754 => 31731,
    13755 => 31732,
    13756 => 31732,
    13757 => 31733,
    13758 => 31734,
    13759 => 31735,
    13760 => 31736,
    13761 => 31736,
    13762 => 31737,
    13763 => 31738,
    13764 => 31739,
    13765 => 31739,
    13766 => 31740,
    13767 => 31741,
    13768 => 31742,
    13769 => 31743,
    13770 => 31743,
    13771 => 31744,
    13772 => 31745,
    13773 => 31746,
    13774 => 31746,
    13775 => 31747,
    13776 => 31748,
    13777 => 31749,
    13778 => 31750,
    13779 => 31750,
    13780 => 31751,
    13781 => 31752,
    13782 => 31753,
    13783 => 31753,
    13784 => 31754,
    13785 => 31755,
    13786 => 31756,
    13787 => 31757,
    13788 => 31757,
    13789 => 31758,
    13790 => 31759,
    13791 => 31760,
    13792 => 31760,
    13793 => 31761,
    13794 => 31762,
    13795 => 31763,
    13796 => 31764,
    13797 => 31764,
    13798 => 31765,
    13799 => 31766,
    13800 => 31767,
    13801 => 31767,
    13802 => 31768,
    13803 => 31769,
    13804 => 31770,
    13805 => 31770,
    13806 => 31771,
    13807 => 31772,
    13808 => 31773,
    13809 => 31774,
    13810 => 31774,
    13811 => 31775,
    13812 => 31776,
    13813 => 31777,
    13814 => 31777,
    13815 => 31778,
    13816 => 31779,
    13817 => 31780,
    13818 => 31780,
    13819 => 31781,
    13820 => 31782,
    13821 => 31783,
    13822 => 31783,
    13823 => 31784,
    13824 => 31785,
    13825 => 31786,
    13826 => 31787,
    13827 => 31787,
    13828 => 31788,
    13829 => 31789,
    13830 => 31790,
    13831 => 31790,
    13832 => 31791,
    13833 => 31792,
    13834 => 31793,
    13835 => 31793,
    13836 => 31794,
    13837 => 31795,
    13838 => 31796,
    13839 => 31796,
    13840 => 31797,
    13841 => 31798,
    13842 => 31799,
    13843 => 31799,
    13844 => 31800,
    13845 => 31801,
    13846 => 31802,
    13847 => 31802,
    13848 => 31803,
    13849 => 31804,
    13850 => 31805,
    13851 => 31806,
    13852 => 31806,
    13853 => 31807,
    13854 => 31808,
    13855 => 31809,
    13856 => 31809,
    13857 => 31810,
    13858 => 31811,
    13859 => 31812,
    13860 => 31812,
    13861 => 31813,
    13862 => 31814,
    13863 => 31815,
    13864 => 31815,
    13865 => 31816,
    13866 => 31817,
    13867 => 31818,
    13868 => 31818,
    13869 => 31819,
    13870 => 31820,
    13871 => 31821,
    13872 => 31821,
    13873 => 31822,
    13874 => 31823,
    13875 => 31824,
    13876 => 31824,
    13877 => 31825,
    13878 => 31826,
    13879 => 31827,
    13880 => 31827,
    13881 => 31828,
    13882 => 31829,
    13883 => 31830,
    13884 => 31830,
    13885 => 31831,
    13886 => 31832,
    13887 => 31833,
    13888 => 31833,
    13889 => 31834,
    13890 => 31835,
    13891 => 31836,
    13892 => 31836,
    13893 => 31837,
    13894 => 31838,
    13895 => 31838,
    13896 => 31839,
    13897 => 31840,
    13898 => 31841,
    13899 => 31841,
    13900 => 31842,
    13901 => 31843,
    13902 => 31844,
    13903 => 31844,
    13904 => 31845,
    13905 => 31846,
    13906 => 31847,
    13907 => 31847,
    13908 => 31848,
    13909 => 31849,
    13910 => 31850,
    13911 => 31850,
    13912 => 31851,
    13913 => 31852,
    13914 => 31853,
    13915 => 31853,
    13916 => 31854,
    13917 => 31855,
    13918 => 31855,
    13919 => 31856,
    13920 => 31857,
    13921 => 31858,
    13922 => 31858,
    13923 => 31859,
    13924 => 31860,
    13925 => 31861,
    13926 => 31861,
    13927 => 31862,
    13928 => 31863,
    13929 => 31864,
    13930 => 31864,
    13931 => 31865,
    13932 => 31866,
    13933 => 31866,
    13934 => 31867,
    13935 => 31868,
    13936 => 31869,
    13937 => 31869,
    13938 => 31870,
    13939 => 31871,
    13940 => 31872,
    13941 => 31872,
    13942 => 31873,
    13943 => 31874,
    13944 => 31875,
    13945 => 31875,
    13946 => 31876,
    13947 => 31877,
    13948 => 31877,
    13949 => 31878,
    13950 => 31879,
    13951 => 31880,
    13952 => 31880,
    13953 => 31881,
    13954 => 31882,
    13955 => 31882,
    13956 => 31883,
    13957 => 31884,
    13958 => 31885,
    13959 => 31885,
    13960 => 31886,
    13961 => 31887,
    13962 => 31888,
    13963 => 31888,
    13964 => 31889,
    13965 => 31890,
    13966 => 31890,
    13967 => 31891,
    13968 => 31892,
    13969 => 31893,
    13970 => 31893,
    13971 => 31894,
    13972 => 31895,
    13973 => 31896,
    13974 => 31896,
    13975 => 31897,
    13976 => 31898,
    13977 => 31898,
    13978 => 31899,
    13979 => 31900,
    13980 => 31901,
    13981 => 31901,
    13982 => 31902,
    13983 => 31903,
    13984 => 31903,
    13985 => 31904,
    13986 => 31905,
    13987 => 31906,
    13988 => 31906,
    13989 => 31907,
    13990 => 31908,
    13991 => 31908,
    13992 => 31909,
    13993 => 31910,
    13994 => 31911,
    13995 => 31911,
    13996 => 31912,
    13997 => 31913,
    13998 => 31913,
    13999 => 31914,
    14000 => 31915,
    14001 => 31916,
    14002 => 31916,
    14003 => 31917,
    14004 => 31918,
    14005 => 31918,
    14006 => 31919,
    14007 => 31920,
    14008 => 31921,
    14009 => 31921,
    14010 => 31922,
    14011 => 31923,
    14012 => 31923,
    14013 => 31924,
    14014 => 31925,
    14015 => 31925,
    14016 => 31926,
    14017 => 31927,
    14018 => 31928,
    14019 => 31928,
    14020 => 31929,
    14021 => 31930,
    14022 => 31930,
    14023 => 31931,
    14024 => 31932,
    14025 => 31933,
    14026 => 31933,
    14027 => 31934,
    14028 => 31935,
    14029 => 31935,
    14030 => 31936,
    14031 => 31937,
    14032 => 31937,
    14033 => 31938,
    14034 => 31939,
    14035 => 31940,
    14036 => 31940,
    14037 => 31941,
    14038 => 31942,
    14039 => 31942,
    14040 => 31943,
    14041 => 31944,
    14042 => 31944,
    14043 => 31945,
    14044 => 31946,
    14045 => 31947,
    14046 => 31947,
    14047 => 31948,
    14048 => 31949,
    14049 => 31949,
    14050 => 31950,
    14051 => 31951,
    14052 => 31951,
    14053 => 31952,
    14054 => 31953,
    14055 => 31954,
    14056 => 31954,
    14057 => 31955,
    14058 => 31956,
    14059 => 31956,
    14060 => 31957,
    14061 => 31958,
    14062 => 31958,
    14063 => 31959,
    14064 => 31960,
    14065 => 31960,
    14066 => 31961,
    14067 => 31962,
    14068 => 31963,
    14069 => 31963,
    14070 => 31964,
    14071 => 31965,
    14072 => 31965,
    14073 => 31966,
    14074 => 31967,
    14075 => 31967,
    14076 => 31968,
    14077 => 31969,
    14078 => 31969,
    14079 => 31970,
    14080 => 31971,
    14081 => 31972,
    14082 => 31972,
    14083 => 31973,
    14084 => 31974,
    14085 => 31974,
    14086 => 31975,
    14087 => 31976,
    14088 => 31976,
    14089 => 31977,
    14090 => 31978,
    14091 => 31978,
    14092 => 31979,
    14093 => 31980,
    14094 => 31980,
    14095 => 31981,
    14096 => 31982,
    14097 => 31982,
    14098 => 31983,
    14099 => 31984,
    14100 => 31985,
    14101 => 31985,
    14102 => 31986,
    14103 => 31987,
    14104 => 31987,
    14105 => 31988,
    14106 => 31989,
    14107 => 31989,
    14108 => 31990,
    14109 => 31991,
    14110 => 31991,
    14111 => 31992,
    14112 => 31993,
    14113 => 31993,
    14114 => 31994,
    14115 => 31995,
    14116 => 31995,
    14117 => 31996,
    14118 => 31997,
    14119 => 31997,
    14120 => 31998,
    14121 => 31999,
    14122 => 31999,
    14123 => 32000,
    14124 => 32001,
    14125 => 32002,
    14126 => 32002,
    14127 => 32003,
    14128 => 32004,
    14129 => 32004,
    14130 => 32005,
    14131 => 32006,
    14132 => 32006,
    14133 => 32007,
    14134 => 32008,
    14135 => 32008,
    14136 => 32009,
    14137 => 32010,
    14138 => 32010,
    14139 => 32011,
    14140 => 32012,
    14141 => 32012,
    14142 => 32013,
    14143 => 32014,
    14144 => 32014,
    14145 => 32015,
    14146 => 32016,
    14147 => 32016,
    14148 => 32017,
    14149 => 32018,
    14150 => 32018,
    14151 => 32019,
    14152 => 32020,
    14153 => 32020,
    14154 => 32021,
    14155 => 32022,
    14156 => 32022,
    14157 => 32023,
    14158 => 32024,
    14159 => 32024,
    14160 => 32025,
    14161 => 32026,
    14162 => 32026,
    14163 => 32027,
    14164 => 32028,
    14165 => 32028,
    14166 => 32029,
    14167 => 32030,
    14168 => 32030,
    14169 => 32031,
    14170 => 32032,
    14171 => 32032,
    14172 => 32033,
    14173 => 32034,
    14174 => 32034,
    14175 => 32035,
    14176 => 32036,
    14177 => 32036,
    14178 => 32037,
    14179 => 32038,
    14180 => 32038,
    14181 => 32039,
    14182 => 32040,
    14183 => 32040,
    14184 => 32041,
    14185 => 32041,
    14186 => 32042,
    14187 => 32043,
    14188 => 32043,
    14189 => 32044,
    14190 => 32045,
    14191 => 32045,
    14192 => 32046,
    14193 => 32047,
    14194 => 32047,
    14195 => 32048,
    14196 => 32049,
    14197 => 32049,
    14198 => 32050,
    14199 => 32051,
    14200 => 32051,
    14201 => 32052,
    14202 => 32053,
    14203 => 32053,
    14204 => 32054,
    14205 => 32055,
    14206 => 32055,
    14207 => 32056,
    14208 => 32057,
    14209 => 32057,
    14210 => 32058,
    14211 => 32058,
    14212 => 32059,
    14213 => 32060,
    14214 => 32060,
    14215 => 32061,
    14216 => 32062,
    14217 => 32062,
    14218 => 32063,
    14219 => 32064,
    14220 => 32064,
    14221 => 32065,
    14222 => 32066,
    14223 => 32066,
    14224 => 32067,
    14225 => 32068,
    14226 => 32068,
    14227 => 32069,
    14228 => 32069,
    14229 => 32070,
    14230 => 32071,
    14231 => 32071,
    14232 => 32072,
    14233 => 32073,
    14234 => 32073,
    14235 => 32074,
    14236 => 32075,
    14237 => 32075,
    14238 => 32076,
    14239 => 32077,
    14240 => 32077,
    14241 => 32078,
    14242 => 32078,
    14243 => 32079,
    14244 => 32080,
    14245 => 32080,
    14246 => 32081,
    14247 => 32082,
    14248 => 32082,
    14249 => 32083,
    14250 => 32084,
    14251 => 32084,
    14252 => 32085,
    14253 => 32086,
    14254 => 32086,
    14255 => 32087,
    14256 => 32087,
    14257 => 32088,
    14258 => 32089,
    14259 => 32089,
    14260 => 32090,
    14261 => 32091,
    14262 => 32091,
    14263 => 32092,
    14264 => 32092,
    14265 => 32093,
    14266 => 32094,
    14267 => 32094,
    14268 => 32095,
    14269 => 32096,
    14270 => 32096,
    14271 => 32097,
    14272 => 32098,
    14273 => 32098,
    14274 => 32099,
    14275 => 32099,
    14276 => 32100,
    14277 => 32101,
    14278 => 32101,
    14279 => 32102,
    14280 => 32103,
    14281 => 32103,
    14282 => 32104,
    14283 => 32104,
    14284 => 32105,
    14285 => 32106,
    14286 => 32106,
    14287 => 32107,
    14288 => 32108,
    14289 => 32108,
    14290 => 32109,
    14291 => 32110,
    14292 => 32110,
    14293 => 32111,
    14294 => 32111,
    14295 => 32112,
    14296 => 32113,
    14297 => 32113,
    14298 => 32114,
    14299 => 32115,
    14300 => 32115,
    14301 => 32116,
    14302 => 32116,
    14303 => 32117,
    14304 => 32118,
    14305 => 32118,
    14306 => 32119,
    14307 => 32119,
    14308 => 32120,
    14309 => 32121,
    14310 => 32121,
    14311 => 32122,
    14312 => 32123,
    14313 => 32123,
    14314 => 32124,
    14315 => 32124,
    14316 => 32125,
    14317 => 32126,
    14318 => 32126,
    14319 => 32127,
    14320 => 32128,
    14321 => 32128,
    14322 => 32129,
    14323 => 32129,
    14324 => 32130,
    14325 => 32131,
    14326 => 32131,
    14327 => 32132,
    14328 => 32132,
    14329 => 32133,
    14330 => 32134,
    14331 => 32134,
    14332 => 32135,
    14333 => 32136,
    14334 => 32136,
    14335 => 32137,
    14336 => 32137,
    14337 => 32138,
    14338 => 32139,
    14339 => 32139,
    14340 => 32140,
    14341 => 32140,
    14342 => 32141,
    14343 => 32142,
    14344 => 32142,
    14345 => 32143,
    14346 => 32144,
    14347 => 32144,
    14348 => 32145,
    14349 => 32145,
    14350 => 32146,
    14351 => 32147,
    14352 => 32147,
    14353 => 32148,
    14354 => 32148,
    14355 => 32149,
    14356 => 32150,
    14357 => 32150,
    14358 => 32151,
    14359 => 32151,
    14360 => 32152,
    14361 => 32153,
    14362 => 32153,
    14363 => 32154,
    14364 => 32154,
    14365 => 32155,
    14366 => 32156,
    14367 => 32156,
    14368 => 32157,
    14369 => 32157,
    14370 => 32158,
    14371 => 32159,
    14372 => 32159,
    14373 => 32160,
    14374 => 32160,
    14375 => 32161,
    14376 => 32162,
    14377 => 32162,
    14378 => 32163,
    14379 => 32163,
    14380 => 32164,
    14381 => 32165,
    14382 => 32165,
    14383 => 32166,
    14384 => 32166,
    14385 => 32167,
    14386 => 32168,
    14387 => 32168,
    14388 => 32169,
    14389 => 32169,
    14390 => 32170,
    14391 => 32171,
    14392 => 32171,
    14393 => 32172,
    14394 => 32172,
    14395 => 32173,
    14396 => 32174,
    14397 => 32174,
    14398 => 32175,
    14399 => 32175,
    14400 => 32176,
    14401 => 32177,
    14402 => 32177,
    14403 => 32178,
    14404 => 32178,
    14405 => 32179,
    14406 => 32180,
    14407 => 32180,
    14408 => 32181,
    14409 => 32181,
    14410 => 32182,
    14411 => 32183,
    14412 => 32183,
    14413 => 32184,
    14414 => 32184,
    14415 => 32185,
    14416 => 32185,
    14417 => 32186,
    14418 => 32187,
    14419 => 32187,
    14420 => 32188,
    14421 => 32188,
    14422 => 32189,
    14423 => 32190,
    14424 => 32190,
    14425 => 32191,
    14426 => 32191,
    14427 => 32192,
    14428 => 32193,
    14429 => 32193,
    14430 => 32194,
    14431 => 32194,
    14432 => 32195,
    14433 => 32195,
    14434 => 32196,
    14435 => 32197,
    14436 => 32197,
    14437 => 32198,
    14438 => 32198,
    14439 => 32199,
    14440 => 32200,
    14441 => 32200,
    14442 => 32201,
    14443 => 32201,
    14444 => 32202,
    14445 => 32202,
    14446 => 32203,
    14447 => 32204,
    14448 => 32204,
    14449 => 32205,
    14450 => 32205,
    14451 => 32206,
    14452 => 32206,
    14453 => 32207,
    14454 => 32208,
    14455 => 32208,
    14456 => 32209,
    14457 => 32209,
    14458 => 32210,
    14459 => 32211,
    14460 => 32211,
    14461 => 32212,
    14462 => 32212,
    14463 => 32213,
    14464 => 32213,
    14465 => 32214,
    14466 => 32215,
    14467 => 32215,
    14468 => 32216,
    14469 => 32216,
    14470 => 32217,
    14471 => 32217,
    14472 => 32218,
    14473 => 32219,
    14474 => 32219,
    14475 => 32220,
    14476 => 32220,
    14477 => 32221,
    14478 => 32221,
    14479 => 32222,
    14480 => 32223,
    14481 => 32223,
    14482 => 32224,
    14483 => 32224,
    14484 => 32225,
    14485 => 32225,
    14486 => 32226,
    14487 => 32227,
    14488 => 32227,
    14489 => 32228,
    14490 => 32228,
    14491 => 32229,
    14492 => 32229,
    14493 => 32230,
    14494 => 32231,
    14495 => 32231,
    14496 => 32232,
    14497 => 32232,
    14498 => 32233,
    14499 => 32233,
    14500 => 32234,
    14501 => 32234,
    14502 => 32235,
    14503 => 32236,
    14504 => 32236,
    14505 => 32237,
    14506 => 32237,
    14507 => 32238,
    14508 => 32238,
    14509 => 32239,
    14510 => 32240,
    14511 => 32240,
    14512 => 32241,
    14513 => 32241,
    14514 => 32242,
    14515 => 32242,
    14516 => 32243,
    14517 => 32243,
    14518 => 32244,
    14519 => 32245,
    14520 => 32245,
    14521 => 32246,
    14522 => 32246,
    14523 => 32247,
    14524 => 32247,
    14525 => 32248,
    14526 => 32248,
    14527 => 32249,
    14528 => 32250,
    14529 => 32250,
    14530 => 32251,
    14531 => 32251,
    14532 => 32252,
    14533 => 32252,
    14534 => 32253,
    14535 => 32253,
    14536 => 32254,
    14537 => 32255,
    14538 => 32255,
    14539 => 32256,
    14540 => 32256,
    14541 => 32257,
    14542 => 32257,
    14543 => 32258,
    14544 => 32258,
    14545 => 32259,
    14546 => 32260,
    14547 => 32260,
    14548 => 32261,
    14549 => 32261,
    14550 => 32262,
    14551 => 32262,
    14552 => 32263,
    14553 => 32263,
    14554 => 32264,
    14555 => 32265,
    14556 => 32265,
    14557 => 32266,
    14558 => 32266,
    14559 => 32267,
    14560 => 32267,
    14561 => 32268,
    14562 => 32268,
    14563 => 32269,
    14564 => 32269,
    14565 => 32270,
    14566 => 32271,
    14567 => 32271,
    14568 => 32272,
    14569 => 32272,
    14570 => 32273,
    14571 => 32273,
    14572 => 32274,
    14573 => 32274,
    14574 => 32275,
    14575 => 32275,
    14576 => 32276,
    14577 => 32277,
    14578 => 32277,
    14579 => 32278,
    14580 => 32278,
    14581 => 32279,
    14582 => 32279,
    14583 => 32280,
    14584 => 32280,
    14585 => 32281,
    14586 => 32281,
    14587 => 32282,
    14588 => 32282,
    14589 => 32283,
    14590 => 32284,
    14591 => 32284,
    14592 => 32285,
    14593 => 32285,
    14594 => 32286,
    14595 => 32286,
    14596 => 32287,
    14597 => 32287,
    14598 => 32288,
    14599 => 32288,
    14600 => 32289,
    14601 => 32289,
    14602 => 32290,
    14603 => 32290,
    14604 => 32291,
    14605 => 32292,
    14606 => 32292,
    14607 => 32293,
    14608 => 32293,
    14609 => 32294,
    14610 => 32294,
    14611 => 32295,
    14612 => 32295,
    14613 => 32296,
    14614 => 32296,
    14615 => 32297,
    14616 => 32297,
    14617 => 32298,
    14618 => 32298,
    14619 => 32299,
    14620 => 32300,
    14621 => 32300,
    14622 => 32301,
    14623 => 32301,
    14624 => 32302,
    14625 => 32302,
    14626 => 32303,
    14627 => 32303,
    14628 => 32304,
    14629 => 32304,
    14630 => 32305,
    14631 => 32305,
    14632 => 32306,
    14633 => 32306,
    14634 => 32307,
    14635 => 32307,
    14636 => 32308,
    14637 => 32308,
    14638 => 32309,
    14639 => 32310,
    14640 => 32310,
    14641 => 32311,
    14642 => 32311,
    14643 => 32312,
    14644 => 32312,
    14645 => 32313,
    14646 => 32313,
    14647 => 32314,
    14648 => 32314,
    14649 => 32315,
    14650 => 32315,
    14651 => 32316,
    14652 => 32316,
    14653 => 32317,
    14654 => 32317,
    14655 => 32318,
    14656 => 32318,
    14657 => 32319,
    14658 => 32319,
    14659 => 32320,
    14660 => 32320,
    14661 => 32321,
    14662 => 32321,
    14663 => 32322,
    14664 => 32322,
    14665 => 32323,
    14666 => 32324,
    14667 => 32324,
    14668 => 32325,
    14669 => 32325,
    14670 => 32326,
    14671 => 32326,
    14672 => 32327,
    14673 => 32327,
    14674 => 32328,
    14675 => 32328,
    14676 => 32329,
    14677 => 32329,
    14678 => 32330,
    14679 => 32330,
    14680 => 32331,
    14681 => 32331,
    14682 => 32332,
    14683 => 32332,
    14684 => 32333,
    14685 => 32333,
    14686 => 32334,
    14687 => 32334,
    14688 => 32335,
    14689 => 32335,
    14690 => 32336,
    14691 => 32336,
    14692 => 32337,
    14693 => 32337,
    14694 => 32338,
    14695 => 32338,
    14696 => 32339,
    14697 => 32339,
    14698 => 32340,
    14699 => 32340,
    14700 => 32341,
    14701 => 32341,
    14702 => 32342,
    14703 => 32342,
    14704 => 32343,
    14705 => 32343,
    14706 => 32344,
    14707 => 32344,
    14708 => 32345,
    14709 => 32345,
    14710 => 32346,
    14711 => 32346,
    14712 => 32347,
    14713 => 32347,
    14714 => 32348,
    14715 => 32348,
    14716 => 32349,
    14717 => 32349,
    14718 => 32350,
    14719 => 32350,
    14720 => 32351,
    14721 => 32351,
    14722 => 32352,
    14723 => 32352,
    14724 => 32353,
    14725 => 32353,
    14726 => 32354,
    14727 => 32354,
    14728 => 32355,
    14729 => 32355,
    14730 => 32356,
    14731 => 32356,
    14732 => 32357,
    14733 => 32357,
    14734 => 32358,
    14735 => 32358,
    14736 => 32359,
    14737 => 32359,
    14738 => 32360,
    14739 => 32360,
    14740 => 32361,
    14741 => 32361,
    14742 => 32362,
    14743 => 32362,
    14744 => 32363,
    14745 => 32363,
    14746 => 32364,
    14747 => 32364,
    14748 => 32365,
    14749 => 32365,
    14750 => 32366,
    14751 => 32366,
    14752 => 32367,
    14753 => 32367,
    14754 => 32368,
    14755 => 32368,
    14756 => 32369,
    14757 => 32369,
    14758 => 32370,
    14759 => 32370,
    14760 => 32371,
    14761 => 32371,
    14762 => 32372,
    14763 => 32372,
    14764 => 32373,
    14765 => 32373,
    14766 => 32374,
    14767 => 32374,
    14768 => 32375,
    14769 => 32375,
    14770 => 32375,
    14771 => 32376,
    14772 => 32376,
    14773 => 32377,
    14774 => 32377,
    14775 => 32378,
    14776 => 32378,
    14777 => 32379,
    14778 => 32379,
    14779 => 32380,
    14780 => 32380,
    14781 => 32381,
    14782 => 32381,
    14783 => 32382,
    14784 => 32382,
    14785 => 32383,
    14786 => 32383,
    14787 => 32384,
    14788 => 32384,
    14789 => 32385,
    14790 => 32385,
    14791 => 32386,
    14792 => 32386,
    14793 => 32387,
    14794 => 32387,
    14795 => 32387,
    14796 => 32388,
    14797 => 32388,
    14798 => 32389,
    14799 => 32389,
    14800 => 32390,
    14801 => 32390,
    14802 => 32391,
    14803 => 32391,
    14804 => 32392,
    14805 => 32392,
    14806 => 32393,
    14807 => 32393,
    14808 => 32394,
    14809 => 32394,
    14810 => 32395,
    14811 => 32395,
    14812 => 32396,
    14813 => 32396,
    14814 => 32397,
    14815 => 32397,
    14816 => 32397,
    14817 => 32398,
    14818 => 32398,
    14819 => 32399,
    14820 => 32399,
    14821 => 32400,
    14822 => 32400,
    14823 => 32401,
    14824 => 32401,
    14825 => 32402,
    14826 => 32402,
    14827 => 32403,
    14828 => 32403,
    14829 => 32404,
    14830 => 32404,
    14831 => 32404,
    14832 => 32405,
    14833 => 32405,
    14834 => 32406,
    14835 => 32406,
    14836 => 32407,
    14837 => 32407,
    14838 => 32408,
    14839 => 32408,
    14840 => 32409,
    14841 => 32409,
    14842 => 32410,
    14843 => 32410,
    14844 => 32411,
    14845 => 32411,
    14846 => 32411,
    14847 => 32412,
    14848 => 32412,
    14849 => 32413,
    14850 => 32413,
    14851 => 32414,
    14852 => 32414,
    14853 => 32415,
    14854 => 32415,
    14855 => 32416,
    14856 => 32416,
    14857 => 32416,
    14858 => 32417,
    14859 => 32417,
    14860 => 32418,
    14861 => 32418,
    14862 => 32419,
    14863 => 32419,
    14864 => 32420,
    14865 => 32420,
    14866 => 32421,
    14867 => 32421,
    14868 => 32422,
    14869 => 32422,
    14870 => 32422,
    14871 => 32423,
    14872 => 32423,
    14873 => 32424,
    14874 => 32424,
    14875 => 32425,
    14876 => 32425,
    14877 => 32426,
    14878 => 32426,
    14879 => 32426,
    14880 => 32427,
    14881 => 32427,
    14882 => 32428,
    14883 => 32428,
    14884 => 32429,
    14885 => 32429,
    14886 => 32430,
    14887 => 32430,
    14888 => 32431,
    14889 => 32431,
    14890 => 32431,
    14891 => 32432,
    14892 => 32432,
    14893 => 32433,
    14894 => 32433,
    14895 => 32434,
    14896 => 32434,
    14897 => 32435,
    14898 => 32435,
    14899 => 32435,
    14900 => 32436,
    14901 => 32436,
    14902 => 32437,
    14903 => 32437,
    14904 => 32438,
    14905 => 32438,
    14906 => 32439,
    14907 => 32439,
    14908 => 32439,
    14909 => 32440,
    14910 => 32440,
    14911 => 32441,
    14912 => 32441,
    14913 => 32442,
    14914 => 32442,
    14915 => 32443,
    14916 => 32443,
    14917 => 32443,
    14918 => 32444,
    14919 => 32444,
    14920 => 32445,
    14921 => 32445,
    14922 => 32446,
    14923 => 32446,
    14924 => 32447,
    14925 => 32447,
    14926 => 32447,
    14927 => 32448,
    14928 => 32448,
    14929 => 32449,
    14930 => 32449,
    14931 => 32450,
    14932 => 32450,
    14933 => 32450,
    14934 => 32451,
    14935 => 32451,
    14936 => 32452,
    14937 => 32452,
    14938 => 32453,
    14939 => 32453,
    14940 => 32453,
    14941 => 32454,
    14942 => 32454,
    14943 => 32455,
    14944 => 32455,
    14945 => 32456,
    14946 => 32456,
    14947 => 32457,
    14948 => 32457,
    14949 => 32457,
    14950 => 32458,
    14951 => 32458,
    14952 => 32459,
    14953 => 32459,
    14954 => 32460,
    14955 => 32460,
    14956 => 32460,
    14957 => 32461,
    14958 => 32461,
    14959 => 32462,
    14960 => 32462,
    14961 => 32463,
    14962 => 32463,
    14963 => 32463,
    14964 => 32464,
    14965 => 32464,
    14966 => 32465,
    14967 => 32465,
    14968 => 32466,
    14969 => 32466,
    14970 => 32466,
    14971 => 32467,
    14972 => 32467,
    14973 => 32468,
    14974 => 32468,
    14975 => 32468,
    14976 => 32469,
    14977 => 32469,
    14978 => 32470,
    14979 => 32470,
    14980 => 32471,
    14981 => 32471,
    14982 => 32471,
    14983 => 32472,
    14984 => 32472,
    14985 => 32473,
    14986 => 32473,
    14987 => 32474,
    14988 => 32474,
    14989 => 32474,
    14990 => 32475,
    14991 => 32475,
    14992 => 32476,
    14993 => 32476,
    14994 => 32476,
    14995 => 32477,
    14996 => 32477,
    14997 => 32478,
    14998 => 32478,
    14999 => 32479,
    15000 => 32479,
    15001 => 32479,
    15002 => 32480,
    15003 => 32480,
    15004 => 32481,
    15005 => 32481,
    15006 => 32481,
    15007 => 32482,
    15008 => 32482,
    15009 => 32483,
    15010 => 32483,
    15011 => 32484,
    15012 => 32484,
    15013 => 32484,
    15014 => 32485,
    15015 => 32485,
    15016 => 32486,
    15017 => 32486,
    15018 => 32486,
    15019 => 32487,
    15020 => 32487,
    15021 => 32488,
    15022 => 32488,
    15023 => 32488,
    15024 => 32489,
    15025 => 32489,
    15026 => 32490,
    15027 => 32490,
    15028 => 32490,
    15029 => 32491,
    15030 => 32491,
    15031 => 32492,
    15032 => 32492,
    15033 => 32493,
    15034 => 32493,
    15035 => 32493,
    15036 => 32494,
    15037 => 32494,
    15038 => 32495,
    15039 => 32495,
    15040 => 32495,
    15041 => 32496,
    15042 => 32496,
    15043 => 32497,
    15044 => 32497,
    15045 => 32497,
    15046 => 32498,
    15047 => 32498,
    15048 => 32499,
    15049 => 32499,
    15050 => 32499,
    15051 => 32500,
    15052 => 32500,
    15053 => 32501,
    15054 => 32501,
    15055 => 32501,
    15056 => 32502,
    15057 => 32502,
    15058 => 32503,
    15059 => 32503,
    15060 => 32503,
    15061 => 32504,
    15062 => 32504,
    15063 => 32505,
    15064 => 32505,
    15065 => 32505,
    15066 => 32506,
    15067 => 32506,
    15068 => 32507,
    15069 => 32507,
    15070 => 32507,
    15071 => 32508,
    15072 => 32508,
    15073 => 32509,
    15074 => 32509,
    15075 => 32509,
    15076 => 32510,
    15077 => 32510,
    15078 => 32510,
    15079 => 32511,
    15080 => 32511,
    15081 => 32512,
    15082 => 32512,
    15083 => 32512,
    15084 => 32513,
    15085 => 32513,
    15086 => 32514,
    15087 => 32514,
    15088 => 32514,
    15089 => 32515,
    15090 => 32515,
    15091 => 32516,
    15092 => 32516,
    15093 => 32516,
    15094 => 32517,
    15095 => 32517,
    15096 => 32517,
    15097 => 32518,
    15098 => 32518,
    15099 => 32519,
    15100 => 32519,
    15101 => 32519,
    15102 => 32520,
    15103 => 32520,
    15104 => 32521,
    15105 => 32521,
    15106 => 32521,
    15107 => 32522,
    15108 => 32522,
    15109 => 32522,
    15110 => 32523,
    15111 => 32523,
    15112 => 32524,
    15113 => 32524,
    15114 => 32524,
    15115 => 32525,
    15116 => 32525,
    15117 => 32526,
    15118 => 32526,
    15119 => 32526,
    15120 => 32527,
    15121 => 32527,
    15122 => 32527,
    15123 => 32528,
    15124 => 32528,
    15125 => 32529,
    15126 => 32529,
    15127 => 32529,
    15128 => 32530,
    15129 => 32530,
    15130 => 32530,
    15131 => 32531,
    15132 => 32531,
    15133 => 32532,
    15134 => 32532,
    15135 => 32532,
    15136 => 32533,
    15137 => 32533,
    15138 => 32533,
    15139 => 32534,
    15140 => 32534,
    15141 => 32535,
    15142 => 32535,
    15143 => 32535,
    15144 => 32536,
    15145 => 32536,
    15146 => 32536,
    15147 => 32537,
    15148 => 32537,
    15149 => 32538,
    15150 => 32538,
    15151 => 32538,
    15152 => 32539,
    15153 => 32539,
    15154 => 32539,
    15155 => 32540,
    15156 => 32540,
    15157 => 32541,
    15158 => 32541,
    15159 => 32541,
    15160 => 32542,
    15161 => 32542,
    15162 => 32542,
    15163 => 32543,
    15164 => 32543,
    15165 => 32543,
    15166 => 32544,
    15167 => 32544,
    15168 => 32545,
    15169 => 32545,
    15170 => 32545,
    15171 => 32546,
    15172 => 32546,
    15173 => 32546,
    15174 => 32547,
    15175 => 32547,
    15176 => 32547,
    15177 => 32548,
    15178 => 32548,
    15179 => 32549,
    15180 => 32549,
    15181 => 32549,
    15182 => 32550,
    15183 => 32550,
    15184 => 32550,
    15185 => 32551,
    15186 => 32551,
    15187 => 32551,
    15188 => 32552,
    15189 => 32552,
    15190 => 32553,
    15191 => 32553,
    15192 => 32553,
    15193 => 32554,
    15194 => 32554,
    15195 => 32554,
    15196 => 32555,
    15197 => 32555,
    15198 => 32555,
    15199 => 32556,
    15200 => 32556,
    15201 => 32556,
    15202 => 32557,
    15203 => 32557,
    15204 => 32558,
    15205 => 32558,
    15206 => 32558,
    15207 => 32559,
    15208 => 32559,
    15209 => 32559,
    15210 => 32560,
    15211 => 32560,
    15212 => 32560,
    15213 => 32561,
    15214 => 32561,
    15215 => 32561,
    15216 => 32562,
    15217 => 32562,
    15218 => 32562,
    15219 => 32563,
    15220 => 32563,
    15221 => 32564,
    15222 => 32564,
    15223 => 32564,
    15224 => 32565,
    15225 => 32565,
    15226 => 32565,
    15227 => 32566,
    15228 => 32566,
    15229 => 32566,
    15230 => 32567,
    15231 => 32567,
    15232 => 32567,
    15233 => 32568,
    15234 => 32568,
    15235 => 32568,
    15236 => 32569,
    15237 => 32569,
    15238 => 32569,
    15239 => 32570,
    15240 => 32570,
    15241 => 32570,
    15242 => 32571,
    15243 => 32571,
    15244 => 32571,
    15245 => 32572,
    15246 => 32572,
    15247 => 32573,
    15248 => 32573,
    15249 => 32573,
    15250 => 32574,
    15251 => 32574,
    15252 => 32574,
    15253 => 32575,
    15254 => 32575,
    15255 => 32575,
    15256 => 32576,
    15257 => 32576,
    15258 => 32576,
    15259 => 32577,
    15260 => 32577,
    15261 => 32577,
    15262 => 32578,
    15263 => 32578,
    15264 => 32578,
    15265 => 32579,
    15266 => 32579,
    15267 => 32579,
    15268 => 32580,
    15269 => 32580,
    15270 => 32580,
    15271 => 32581,
    15272 => 32581,
    15273 => 32581,
    15274 => 32582,
    15275 => 32582,
    15276 => 32582,
    15277 => 32583,
    15278 => 32583,
    15279 => 32583,
    15280 => 32584,
    15281 => 32584,
    15282 => 32584,
    15283 => 32585,
    15284 => 32585,
    15285 => 32585,
    15286 => 32586,
    15287 => 32586,
    15288 => 32586,
    15289 => 32587,
    15290 => 32587,
    15291 => 32587,
    15292 => 32588,
    15293 => 32588,
    15294 => 32588,
    15295 => 32589,
    15296 => 32589,
    15297 => 32589,
    15298 => 32590,
    15299 => 32590,
    15300 => 32590,
    15301 => 32591,
    15302 => 32591,
    15303 => 32591,
    15304 => 32592,
    15305 => 32592,
    15306 => 32592,
    15307 => 32592,
    15308 => 32593,
    15309 => 32593,
    15310 => 32593,
    15311 => 32594,
    15312 => 32594,
    15313 => 32594,
    15314 => 32595,
    15315 => 32595,
    15316 => 32595,
    15317 => 32596,
    15318 => 32596,
    15319 => 32596,
    15320 => 32597,
    15321 => 32597,
    15322 => 32597,
    15323 => 32598,
    15324 => 32598,
    15325 => 32598,
    15326 => 32599,
    15327 => 32599,
    15328 => 32599,
    15329 => 32600,
    15330 => 32600,
    15331 => 32600,
    15332 => 32600,
    15333 => 32601,
    15334 => 32601,
    15335 => 32601,
    15336 => 32602,
    15337 => 32602,
    15338 => 32602,
    15339 => 32603,
    15340 => 32603,
    15341 => 32603,
    15342 => 32604,
    15343 => 32604,
    15344 => 32604,
    15345 => 32605,
    15346 => 32605,
    15347 => 32605,
    15348 => 32606,
    15349 => 32606,
    15350 => 32606,
    15351 => 32606,
    15352 => 32607,
    15353 => 32607,
    15354 => 32607,
    15355 => 32608,
    15356 => 32608,
    15357 => 32608,
    15358 => 32609,
    15359 => 32609,
    15360 => 32609,
    15361 => 32610,
    15362 => 32610,
    15363 => 32610,
    15364 => 32610,
    15365 => 32611,
    15366 => 32611,
    15367 => 32611,
    15368 => 32612,
    15369 => 32612,
    15370 => 32612,
    15371 => 32613,
    15372 => 32613,
    15373 => 32613,
    15374 => 32613,
    15375 => 32614,
    15376 => 32614,
    15377 => 32614,
    15378 => 32615,
    15379 => 32615,
    15380 => 32615,
    15381 => 32616,
    15382 => 32616,
    15383 => 32616,
    15384 => 32617,
    15385 => 32617,
    15386 => 32617,
    15387 => 32617,
    15388 => 32618,
    15389 => 32618,
    15390 => 32618,
    15391 => 32619,
    15392 => 32619,
    15393 => 32619,
    15394 => 32620,
    15395 => 32620,
    15396 => 32620,
    15397 => 32620,
    15398 => 32621,
    15399 => 32621,
    15400 => 32621,
    15401 => 32622,
    15402 => 32622,
    15403 => 32622,
    15404 => 32622,
    15405 => 32623,
    15406 => 32623,
    15407 => 32623,
    15408 => 32624,
    15409 => 32624,
    15410 => 32624,
    15411 => 32625,
    15412 => 32625,
    15413 => 32625,
    15414 => 32625,
    15415 => 32626,
    15416 => 32626,
    15417 => 32626,
    15418 => 32627,
    15419 => 32627,
    15420 => 32627,
    15421 => 32627,
    15422 => 32628,
    15423 => 32628,
    15424 => 32628,
    15425 => 32629,
    15426 => 32629,
    15427 => 32629,
    15428 => 32629,
    15429 => 32630,
    15430 => 32630,
    15431 => 32630,
    15432 => 32631,
    15433 => 32631,
    15434 => 32631,
    15435 => 32631,
    15436 => 32632,
    15437 => 32632,
    15438 => 32632,
    15439 => 32633,
    15440 => 32633,
    15441 => 32633,
    15442 => 32633,
    15443 => 32634,
    15444 => 32634,
    15445 => 32634,
    15446 => 32635,
    15447 => 32635,
    15448 => 32635,
    15449 => 32635,
    15450 => 32636,
    15451 => 32636,
    15452 => 32636,
    15453 => 32637,
    15454 => 32637,
    15455 => 32637,
    15456 => 32637,
    15457 => 32638,
    15458 => 32638,
    15459 => 32638,
    15460 => 32639,
    15461 => 32639,
    15462 => 32639,
    15463 => 32639,
    15464 => 32640,
    15465 => 32640,
    15466 => 32640,
    15467 => 32640,
    15468 => 32641,
    15469 => 32641,
    15470 => 32641,
    15471 => 32642,
    15472 => 32642,
    15473 => 32642,
    15474 => 32642,
    15475 => 32643,
    15476 => 32643,
    15477 => 32643,
    15478 => 32643,
    15479 => 32644,
    15480 => 32644,
    15481 => 32644,
    15482 => 32645,
    15483 => 32645,
    15484 => 32645,
    15485 => 32645,
    15486 => 32646,
    15487 => 32646,
    15488 => 32646,
    15489 => 32646,
    15490 => 32647,
    15491 => 32647,
    15492 => 32647,
    15493 => 32648,
    15494 => 32648,
    15495 => 32648,
    15496 => 32648,
    15497 => 32649,
    15498 => 32649,
    15499 => 32649,
    15500 => 32649,
    15501 => 32650,
    15502 => 32650,
    15503 => 32650,
    15504 => 32650,
    15505 => 32651,
    15506 => 32651,
    15507 => 32651,
    15508 => 32652,
    15509 => 32652,
    15510 => 32652,
    15511 => 32652,
    15512 => 32653,
    15513 => 32653,
    15514 => 32653,
    15515 => 32653,
    15516 => 32654,
    15517 => 32654,
    15518 => 32654,
    15519 => 32654,
    15520 => 32655,
    15521 => 32655,
    15522 => 32655,
    15523 => 32655,
    15524 => 32656,
    15525 => 32656,
    15526 => 32656,
    15527 => 32656,
    15528 => 32657,
    15529 => 32657,
    15530 => 32657,
    15531 => 32657,
    15532 => 32658,
    15533 => 32658,
    15534 => 32658,
    15535 => 32659,
    15536 => 32659,
    15537 => 32659,
    15538 => 32659,
    15539 => 32660,
    15540 => 32660,
    15541 => 32660,
    15542 => 32660,
    15543 => 32661,
    15544 => 32661,
    15545 => 32661,
    15546 => 32661,
    15547 => 32662,
    15548 => 32662,
    15549 => 32662,
    15550 => 32662,
    15551 => 32663,
    15552 => 32663,
    15553 => 32663,
    15554 => 32663,
    15555 => 32664,
    15556 => 32664,
    15557 => 32664,
    15558 => 32664,
    15559 => 32665,
    15560 => 32665,
    15561 => 32665,
    15562 => 32665,
    15563 => 32666,
    15564 => 32666,
    15565 => 32666,
    15566 => 32666,
    15567 => 32667,
    15568 => 32667,
    15569 => 32667,
    15570 => 32667,
    15571 => 32668,
    15572 => 32668,
    15573 => 32668,
    15574 => 32668,
    15575 => 32668,
    15576 => 32669,
    15577 => 32669,
    15578 => 32669,
    15579 => 32669,
    15580 => 32670,
    15581 => 32670,
    15582 => 32670,
    15583 => 32670,
    15584 => 32671,
    15585 => 32671,
    15586 => 32671,
    15587 => 32671,
    15588 => 32672,
    15589 => 32672,
    15590 => 32672,
    15591 => 32672,
    15592 => 32673,
    15593 => 32673,
    15594 => 32673,
    15595 => 32673,
    15596 => 32674,
    15597 => 32674,
    15598 => 32674,
    15599 => 32674,
    15600 => 32674,
    15601 => 32675,
    15602 => 32675,
    15603 => 32675,
    15604 => 32675,
    15605 => 32676,
    15606 => 32676,
    15607 => 32676,
    15608 => 32676,
    15609 => 32677,
    15610 => 32677,
    15611 => 32677,
    15612 => 32677,
    15613 => 32678,
    15614 => 32678,
    15615 => 32678,
    15616 => 32678,
    15617 => 32678,
    15618 => 32679,
    15619 => 32679,
    15620 => 32679,
    15621 => 32679,
    15622 => 32680,
    15623 => 32680,
    15624 => 32680,
    15625 => 32680,
    15626 => 32681,
    15627 => 32681,
    15628 => 32681,
    15629 => 32681,
    15630 => 32681,
    15631 => 32682,
    15632 => 32682,
    15633 => 32682,
    15634 => 32682,
    15635 => 32683,
    15636 => 32683,
    15637 => 32683,
    15638 => 32683,
    15639 => 32683,
    15640 => 32684,
    15641 => 32684,
    15642 => 32684,
    15643 => 32684,
    15644 => 32685,
    15645 => 32685,
    15646 => 32685,
    15647 => 32685,
    15648 => 32685,
    15649 => 32686,
    15650 => 32686,
    15651 => 32686,
    15652 => 32686,
    15653 => 32687,
    15654 => 32687,
    15655 => 32687,
    15656 => 32687,
    15657 => 32687,
    15658 => 32688,
    15659 => 32688,
    15660 => 32688,
    15661 => 32688,
    15662 => 32689,
    15663 => 32689,
    15664 => 32689,
    15665 => 32689,
    15666 => 32689,
    15667 => 32690,
    15668 => 32690,
    15669 => 32690,
    15670 => 32690,
    15671 => 32690,
    15672 => 32691,
    15673 => 32691,
    15674 => 32691,
    15675 => 32691,
    15676 => 32692,
    15677 => 32692,
    15678 => 32692,
    15679 => 32692,
    15680 => 32692,
    15681 => 32693,
    15682 => 32693,
    15683 => 32693,
    15684 => 32693,
    15685 => 32693,
    15686 => 32694,
    15687 => 32694,
    15688 => 32694,
    15689 => 32694,
    15690 => 32694,
    15691 => 32695,
    15692 => 32695,
    15693 => 32695,
    15694 => 32695,
    15695 => 32696,
    15696 => 32696,
    15697 => 32696,
    15698 => 32696,
    15699 => 32696,
    15700 => 32697,
    15701 => 32697,
    15702 => 32697,
    15703 => 32697,
    15704 => 32697,
    15705 => 32698,
    15706 => 32698,
    15707 => 32698,
    15708 => 32698,
    15709 => 32698,
    15710 => 32699,
    15711 => 32699,
    15712 => 32699,
    15713 => 32699,
    15714 => 32699,
    15715 => 32700,
    15716 => 32700,
    15717 => 32700,
    15718 => 32700,
    15719 => 32700,
    15720 => 32701,
    15721 => 32701,
    15722 => 32701,
    15723 => 32701,
    15724 => 32701,
    15725 => 32702,
    15726 => 32702,
    15727 => 32702,
    15728 => 32702,
    15729 => 32702,
    15730 => 32703,
    15731 => 32703,
    15732 => 32703,
    15733 => 32703,
    15734 => 32703,
    15735 => 32704,
    15736 => 32704,
    15737 => 32704,
    15738 => 32704,
    15739 => 32704,
    15740 => 32705,
    15741 => 32705,
    15742 => 32705,
    15743 => 32705,
    15744 => 32705,
    15745 => 32706,
    15746 => 32706,
    15747 => 32706,
    15748 => 32706,
    15749 => 32706,
    15750 => 32706,
    15751 => 32707,
    15752 => 32707,
    15753 => 32707,
    15754 => 32707,
    15755 => 32707,
    15756 => 32708,
    15757 => 32708,
    15758 => 32708,
    15759 => 32708,
    15760 => 32708,
    15761 => 32709,
    15762 => 32709,
    15763 => 32709,
    15764 => 32709,
    15765 => 32709,
    15766 => 32710,
    15767 => 32710,
    15768 => 32710,
    15769 => 32710,
    15770 => 32710,
    15771 => 32710,
    15772 => 32711,
    15773 => 32711,
    15774 => 32711,
    15775 => 32711,
    15776 => 32711,
    15777 => 32712,
    15778 => 32712,
    15779 => 32712,
    15780 => 32712,
    15781 => 32712,
    15782 => 32712,
    15783 => 32713,
    15784 => 32713,
    15785 => 32713,
    15786 => 32713,
    15787 => 32713,
    15788 => 32714,
    15789 => 32714,
    15790 => 32714,
    15791 => 32714,
    15792 => 32714,
    15793 => 32714,
    15794 => 32715,
    15795 => 32715,
    15796 => 32715,
    15797 => 32715,
    15798 => 32715,
    15799 => 32715,
    15800 => 32716,
    15801 => 32716,
    15802 => 32716,
    15803 => 32716,
    15804 => 32716,
    15805 => 32717,
    15806 => 32717,
    15807 => 32717,
    15808 => 32717,
    15809 => 32717,
    15810 => 32717,
    15811 => 32718,
    15812 => 32718,
    15813 => 32718,
    15814 => 32718,
    15815 => 32718,
    15816 => 32718,
    15817 => 32719,
    15818 => 32719,
    15819 => 32719,
    15820 => 32719,
    15821 => 32719,
    15822 => 32719,
    15823 => 32720,
    15824 => 32720,
    15825 => 32720,
    15826 => 32720,
    15827 => 32720,
    15828 => 32720,
    15829 => 32721,
    15830 => 32721,
    15831 => 32721,
    15832 => 32721,
    15833 => 32721,
    15834 => 32721,
    15835 => 32722,
    15836 => 32722,
    15837 => 32722,
    15838 => 32722,
    15839 => 32722,
    15840 => 32722,
    15841 => 32723,
    15842 => 32723,
    15843 => 32723,
    15844 => 32723,
    15845 => 32723,
    15846 => 32723,
    15847 => 32724,
    15848 => 32724,
    15849 => 32724,
    15850 => 32724,
    15851 => 32724,
    15852 => 32724,
    15853 => 32725,
    15854 => 32725,
    15855 => 32725,
    15856 => 32725,
    15857 => 32725,
    15858 => 32725,
    15859 => 32726,
    15860 => 32726,
    15861 => 32726,
    15862 => 32726,
    15863 => 32726,
    15864 => 32726,
    15865 => 32726,
    15866 => 32727,
    15867 => 32727,
    15868 => 32727,
    15869 => 32727,
    15870 => 32727,
    15871 => 32727,
    15872 => 32728,
    15873 => 32728,
    15874 => 32728,
    15875 => 32728,
    15876 => 32728,
    15877 => 32728,
    15878 => 32728,
    15879 => 32729,
    15880 => 32729,
    15881 => 32729,
    15882 => 32729,
    15883 => 32729,
    15884 => 32729,
    15885 => 32730,
    15886 => 32730,
    15887 => 32730,
    15888 => 32730,
    15889 => 32730,
    15890 => 32730,
    15891 => 32730,
    15892 => 32731,
    15893 => 32731,
    15894 => 32731,
    15895 => 32731,
    15896 => 32731,
    15897 => 32731,
    15898 => 32731,
    15899 => 32732,
    15900 => 32732,
    15901 => 32732,
    15902 => 32732,
    15903 => 32732,
    15904 => 32732,
    15905 => 32732,
    15906 => 32733,
    15907 => 32733,
    15908 => 32733,
    15909 => 32733,
    15910 => 32733,
    15911 => 32733,
    15912 => 32733,
    15913 => 32734,
    15914 => 32734,
    15915 => 32734,
    15916 => 32734,
    15917 => 32734,
    15918 => 32734,
    15919 => 32734,
    15920 => 32735,
    15921 => 32735,
    15922 => 32735,
    15923 => 32735,
    15924 => 32735,
    15925 => 32735,
    15926 => 32735,
    15927 => 32736,
    15928 => 32736,
    15929 => 32736,
    15930 => 32736,
    15931 => 32736,
    15932 => 32736,
    15933 => 32736,
    15934 => 32737,
    15935 => 32737,
    15936 => 32737,
    15937 => 32737,
    15938 => 32737,
    15939 => 32737,
    15940 => 32737,
    15941 => 32737,
    15942 => 32738,
    15943 => 32738,
    15944 => 32738,
    15945 => 32738,
    15946 => 32738,
    15947 => 32738,
    15948 => 32738,
    15949 => 32739,
    15950 => 32739,
    15951 => 32739,
    15952 => 32739,
    15953 => 32739,
    15954 => 32739,
    15955 => 32739,
    15956 => 32739,
    15957 => 32740,
    15958 => 32740,
    15959 => 32740,
    15960 => 32740,
    15961 => 32740,
    15962 => 32740,
    15963 => 32740,
    15964 => 32740,
    15965 => 32741,
    15966 => 32741,
    15967 => 32741,
    15968 => 32741,
    15969 => 32741,
    15970 => 32741,
    15971 => 32741,
    15972 => 32741,
    15973 => 32742,
    15974 => 32742,
    15975 => 32742,
    15976 => 32742,
    15977 => 32742,
    15978 => 32742,
    15979 => 32742,
    15980 => 32742,
    15981 => 32743,
    15982 => 32743,
    15983 => 32743,
    15984 => 32743,
    15985 => 32743,
    15986 => 32743,
    15987 => 32743,
    15988 => 32743,
    15989 => 32744,
    15990 => 32744,
    15991 => 32744,
    15992 => 32744,
    15993 => 32744,
    15994 => 32744,
    15995 => 32744,
    15996 => 32744,
    15997 => 32744,
    15998 => 32745,
    15999 => 32745,
    16000 => 32745,
    16001 => 32745,
    16002 => 32745,
    16003 => 32745,
    16004 => 32745,
    16005 => 32745,
    16006 => 32745,
    16007 => 32746,
    16008 => 32746,
    16009 => 32746,
    16010 => 32746,
    16011 => 32746,
    16012 => 32746,
    16013 => 32746,
    16014 => 32746,
    16015 => 32746,
    16016 => 32747,
    16017 => 32747,
    16018 => 32747,
    16019 => 32747,
    16020 => 32747,
    16021 => 32747,
    16022 => 32747,
    16023 => 32747,
    16024 => 32747,
    16025 => 32748,
    16026 => 32748,
    16027 => 32748,
    16028 => 32748,
    16029 => 32748,
    16030 => 32748,
    16031 => 32748,
    16032 => 32748,
    16033 => 32748,
    16034 => 32749,
    16035 => 32749,
    16036 => 32749,
    16037 => 32749,
    16038 => 32749,
    16039 => 32749,
    16040 => 32749,
    16041 => 32749,
    16042 => 32749,
    16043 => 32749,
    16044 => 32750,
    16045 => 32750,
    16046 => 32750,
    16047 => 32750,
    16048 => 32750,
    16049 => 32750,
    16050 => 32750,
    16051 => 32750,
    16052 => 32750,
    16053 => 32751,
    16054 => 32751,
    16055 => 32751,
    16056 => 32751,
    16057 => 32751,
    16058 => 32751,
    16059 => 32751,
    16060 => 32751,
    16061 => 32751,
    16062 => 32751,
    16063 => 32751,
    16064 => 32752,
    16065 => 32752,
    16066 => 32752,
    16067 => 32752,
    16068 => 32752,
    16069 => 32752,
    16070 => 32752,
    16071 => 32752,
    16072 => 32752,
    16073 => 32752,
    16074 => 32753,
    16075 => 32753,
    16076 => 32753,
    16077 => 32753,
    16078 => 32753,
    16079 => 32753,
    16080 => 32753,
    16081 => 32753,
    16082 => 32753,
    16083 => 32753,
    16084 => 32753,
    16085 => 32754,
    16086 => 32754,
    16087 => 32754,
    16088 => 32754,
    16089 => 32754,
    16090 => 32754,
    16091 => 32754,
    16092 => 32754,
    16093 => 32754,
    16094 => 32754,
    16095 => 32754,
    16096 => 32755,
    16097 => 32755,
    16098 => 32755,
    16099 => 32755,
    16100 => 32755,
    16101 => 32755,
    16102 => 32755,
    16103 => 32755,
    16104 => 32755,
    16105 => 32755,
    16106 => 32755,
    16107 => 32755,
    16108 => 32756,
    16109 => 32756,
    16110 => 32756,
    16111 => 32756,
    16112 => 32756,
    16113 => 32756,
    16114 => 32756,
    16115 => 32756,
    16116 => 32756,
    16117 => 32756,
    16118 => 32756,
    16119 => 32756,
    16120 => 32757,
    16121 => 32757,
    16122 => 32757,
    16123 => 32757,
    16124 => 32757,
    16125 => 32757,
    16126 => 32757,
    16127 => 32757,
    16128 => 32757,
    16129 => 32757,
    16130 => 32757,
    16131 => 32757,
    16132 => 32757,
    16133 => 32758,
    16134 => 32758,
    16135 => 32758,
    16136 => 32758,
    16137 => 32758,
    16138 => 32758,
    16139 => 32758,
    16140 => 32758,
    16141 => 32758,
    16142 => 32758,
    16143 => 32758,
    16144 => 32758,
    16145 => 32758,
    16146 => 32758,
    16147 => 32759,
    16148 => 32759,
    16149 => 32759,
    16150 => 32759,
    16151 => 32759,
    16152 => 32759,
    16153 => 32759,
    16154 => 32759,
    16155 => 32759,
    16156 => 32759,
    16157 => 32759,
    16158 => 32759,
    16159 => 32759,
    16160 => 32759,
    16161 => 32760,
    16162 => 32760,
    16163 => 32760,
    16164 => 32760,
    16165 => 32760,
    16166 => 32760,
    16167 => 32760,
    16168 => 32760,
    16169 => 32760,
    16170 => 32760,
    16171 => 32760,
    16172 => 32760,
    16173 => 32760,
    16174 => 32760,
    16175 => 32760,
    16176 => 32760,
    16177 => 32761,
    16178 => 32761,
    16179 => 32761,
    16180 => 32761,
    16181 => 32761,
    16182 => 32761,
    16183 => 32761,
    16184 => 32761,
    16185 => 32761,
    16186 => 32761,
    16187 => 32761,
    16188 => 32761,
    16189 => 32761,
    16190 => 32761,
    16191 => 32761,
    16192 => 32761,
    16193 => 32762,
    16194 => 32762,
    16195 => 32762,
    16196 => 32762,
    16197 => 32762,
    16198 => 32762,
    16199 => 32762,
    16200 => 32762,
    16201 => 32762,
    16202 => 32762,
    16203 => 32762,
    16204 => 32762,
    16205 => 32762,
    16206 => 32762,
    16207 => 32762,
    16208 => 32762,
    16209 => 32762,
    16210 => 32762,
    16211 => 32762,
    16212 => 32763,
    16213 => 32763,
    16214 => 32763,
    16215 => 32763,
    16216 => 32763,
    16217 => 32763,
    16218 => 32763,
    16219 => 32763,
    16220 => 32763,
    16221 => 32763,
    16222 => 32763,
    16223 => 32763,
    16224 => 32763,
    16225 => 32763,
    16226 => 32763,
    16227 => 32763,
    16228 => 32763,
    16229 => 32763,
    16230 => 32763,
    16231 => 32763,
    16232 => 32764,
    16233 => 32764,
    16234 => 32764,
    16235 => 32764,
    16236 => 32764,
    16237 => 32764,
    16238 => 32764,
    16239 => 32764,
    16240 => 32764,
    16241 => 32764,
    16242 => 32764,
    16243 => 32764,
    16244 => 32764,
    16245 => 32764,
    16246 => 32764,
    16247 => 32764,
    16248 => 32764,
    16249 => 32764,
    16250 => 32764,
    16251 => 32764,
    16252 => 32764,
    16253 => 32764,
    16254 => 32764,
    16255 => 32764,
    16256 => 32765,
    16257 => 32765,
    16258 => 32765,
    16259 => 32765,
    16260 => 32765,
    16261 => 32765,
    16262 => 32765,
    16263 => 32765,
    16264 => 32765,
    16265 => 32765,
    16266 => 32765,
    16267 => 32765,
    16268 => 32765,
    16269 => 32765,
    16270 => 32765,
    16271 => 32765,
    16272 => 32765,
    16273 => 32765,
    16274 => 32765,
    16275 => 32765,
    16276 => 32765,
    16277 => 32765,
    16278 => 32765,
    16279 => 32765,
    16280 => 32765,
    16281 => 32765,
    16282 => 32765,
    16283 => 32765,
    16284 => 32765,
    16285 => 32766,
    16286 => 32766,
    16287 => 32766,
    16288 => 32766,
    16289 => 32766,
    16290 => 32766,
    16291 => 32766,
    16292 => 32766,
    16293 => 32766,
    16294 => 32766,
    16295 => 32766,
    16296 => 32766,
    16297 => 32766,
    16298 => 32766,
    16299 => 32766,
    16300 => 32766,
    16301 => 32766,
    16302 => 32766,
    16303 => 32766,
    16304 => 32766,
    16305 => 32766,
    16306 => 32766,
    16307 => 32766,
    16308 => 32766,
    16309 => 32766,
    16310 => 32766,
    16311 => 32766,
    16312 => 32766,
    16313 => 32766,
    16314 => 32766,
    16315 => 32766,
    16316 => 32766,
    16317 => 32766,
    16318 => 32766,
    16319 => 32766,
    16320 => 32766,
    16321 => 32766,
    16322 => 32766,
    16323 => 32766,
    16324 => 32766,
    16325 => 32766,
    16326 => 32766,
    16327 => 32767,
    16328 => 32767,
    16329 => 32767,
    16330 => 32767,
    16331 => 32767,
    16332 => 32767,
    16333 => 32767,
    16334 => 32767,
    16335 => 32767,
    16336 => 32767,
    16337 => 32767,
    16338 => 32767,
    16339 => 32767,
    16340 => 32767,
    16341 => 32767,
    16342 => 32767,
    16343 => 32767,
    16344 => 32767,
    16345 => 32767,
    16346 => 32767,
    16347 => 32767,
    16348 => 32767,
    16349 => 32767,
    16350 => 32767,
    16351 => 32767,
    16352 => 32767,
    16353 => 32767,
    16354 => 32767,
    16355 => 32767,
    16356 => 32767,
    16357 => 32767,
    16358 => 32767,
    16359 => 32767,
    16360 => 32767,
    16361 => 32767,
    16362 => 32767,
    16363 => 32767,
    16364 => 32767,
    16365 => 32767,
    16366 => 32767,
    16367 => 32767,
    16368 => 32767,
    16369 => 32767,
    16370 => 32767,
    16371 => 32767,
    16372 => 32767,
    16373 => 32767,
    16374 => 32767,
    16375 => 32767,
    16376 => 32767,
    16377 => 32767,
    16378 => 32767,
    16379 => 32767,
    16380 => 32767,
    16381 => 32767,
    16382 => 32767,
    16383 => 32767,
    16384 => 32767,
    16385 => 32767,
    16386 => 32767,
    16387 => 32767,
    16388 => 32767,
    16389 => 32767,
    16390 => 32767,
    16391 => 32767,
    16392 => 32767,
    16393 => 32767,
    16394 => 32767,
    16395 => 32767,
    16396 => 32767,
    16397 => 32767,
    16398 => 32767,
    16399 => 32767,
    16400 => 32767,
    16401 => 32767,
    16402 => 32767,
    16403 => 32767,
    16404 => 32767,
    16405 => 32767,
    16406 => 32767,
    16407 => 32767,
    16408 => 32767,
    16409 => 32767,
    16410 => 32767,
    16411 => 32767,
    16412 => 32767,
    16413 => 32767,
    16414 => 32767,
    16415 => 32767,
    16416 => 32767,
    16417 => 32767,
    16418 => 32767,
    16419 => 32767,
    16420 => 32767,
    16421 => 32767,
    16422 => 32767,
    16423 => 32767,
    16424 => 32767,
    16425 => 32767,
    16426 => 32767,
    16427 => 32767,
    16428 => 32767,
    16429 => 32767,
    16430 => 32767,
    16431 => 32767,
    16432 => 32767,
    16433 => 32767,
    16434 => 32767,
    16435 => 32767,
    16436 => 32767,
    16437 => 32767,
    16438 => 32767,
    16439 => 32767,
    16440 => 32767,
    16441 => 32767,
    16442 => 32766,
    16443 => 32766,
    16444 => 32766,
    16445 => 32766,
    16446 => 32766,
    16447 => 32766,
    16448 => 32766,
    16449 => 32766,
    16450 => 32766,
    16451 => 32766,
    16452 => 32766,
    16453 => 32766,
    16454 => 32766,
    16455 => 32766,
    16456 => 32766,
    16457 => 32766,
    16458 => 32766,
    16459 => 32766,
    16460 => 32766,
    16461 => 32766,
    16462 => 32766,
    16463 => 32766,
    16464 => 32766,
    16465 => 32766,
    16466 => 32766,
    16467 => 32766,
    16468 => 32766,
    16469 => 32766,
    16470 => 32766,
    16471 => 32766,
    16472 => 32766,
    16473 => 32766,
    16474 => 32766,
    16475 => 32766,
    16476 => 32766,
    16477 => 32766,
    16478 => 32766,
    16479 => 32766,
    16480 => 32766,
    16481 => 32766,
    16482 => 32766,
    16483 => 32766,
    16484 => 32765,
    16485 => 32765,
    16486 => 32765,
    16487 => 32765,
    16488 => 32765,
    16489 => 32765,
    16490 => 32765,
    16491 => 32765,
    16492 => 32765,
    16493 => 32765,
    16494 => 32765,
    16495 => 32765,
    16496 => 32765,
    16497 => 32765,
    16498 => 32765,
    16499 => 32765,
    16500 => 32765,
    16501 => 32765,
    16502 => 32765,
    16503 => 32765,
    16504 => 32765,
    16505 => 32765,
    16506 => 32765,
    16507 => 32765,
    16508 => 32765,
    16509 => 32765,
    16510 => 32765,
    16511 => 32765,
    16512 => 32765,
    16513 => 32764,
    16514 => 32764,
    16515 => 32764,
    16516 => 32764,
    16517 => 32764,
    16518 => 32764,
    16519 => 32764,
    16520 => 32764,
    16521 => 32764,
    16522 => 32764,
    16523 => 32764,
    16524 => 32764,
    16525 => 32764,
    16526 => 32764,
    16527 => 32764,
    16528 => 32764,
    16529 => 32764,
    16530 => 32764,
    16531 => 32764,
    16532 => 32764,
    16533 => 32764,
    16534 => 32764,
    16535 => 32764,
    16536 => 32764,
    16537 => 32763,
    16538 => 32763,
    16539 => 32763,
    16540 => 32763,
    16541 => 32763,
    16542 => 32763,
    16543 => 32763,
    16544 => 32763,
    16545 => 32763,
    16546 => 32763,
    16547 => 32763,
    16548 => 32763,
    16549 => 32763,
    16550 => 32763,
    16551 => 32763,
    16552 => 32763,
    16553 => 32763,
    16554 => 32763,
    16555 => 32763,
    16556 => 32763,
    16557 => 32762,
    16558 => 32762,
    16559 => 32762,
    16560 => 32762,
    16561 => 32762,
    16562 => 32762,
    16563 => 32762,
    16564 => 32762,
    16565 => 32762,
    16566 => 32762,
    16567 => 32762,
    16568 => 32762,
    16569 => 32762,
    16570 => 32762,
    16571 => 32762,
    16572 => 32762,
    16573 => 32762,
    16574 => 32762,
    16575 => 32762,
    16576 => 32761,
    16577 => 32761,
    16578 => 32761,
    16579 => 32761,
    16580 => 32761,
    16581 => 32761,
    16582 => 32761,
    16583 => 32761,
    16584 => 32761,
    16585 => 32761,
    16586 => 32761,
    16587 => 32761,
    16588 => 32761,
    16589 => 32761,
    16590 => 32761,
    16591 => 32761,
    16592 => 32760,
    16593 => 32760,
    16594 => 32760,
    16595 => 32760,
    16596 => 32760,
    16597 => 32760,
    16598 => 32760,
    16599 => 32760,
    16600 => 32760,
    16601 => 32760,
    16602 => 32760,
    16603 => 32760,
    16604 => 32760,
    16605 => 32760,
    16606 => 32760,
    16607 => 32760,
    16608 => 32759,
    16609 => 32759,
    16610 => 32759,
    16611 => 32759,
    16612 => 32759,
    16613 => 32759,
    16614 => 32759,
    16615 => 32759,
    16616 => 32759,
    16617 => 32759,
    16618 => 32759,
    16619 => 32759,
    16620 => 32759,
    16621 => 32759,
    16622 => 32758,
    16623 => 32758,
    16624 => 32758,
    16625 => 32758,
    16626 => 32758,
    16627 => 32758,
    16628 => 32758,
    16629 => 32758,
    16630 => 32758,
    16631 => 32758,
    16632 => 32758,
    16633 => 32758,
    16634 => 32758,
    16635 => 32758,
    16636 => 32757,
    16637 => 32757,
    16638 => 32757,
    16639 => 32757,
    16640 => 32757,
    16641 => 32757,
    16642 => 32757,
    16643 => 32757,
    16644 => 32757,
    16645 => 32757,
    16646 => 32757,
    16647 => 32757,
    16648 => 32757,
    16649 => 32756,
    16650 => 32756,
    16651 => 32756,
    16652 => 32756,
    16653 => 32756,
    16654 => 32756,
    16655 => 32756,
    16656 => 32756,
    16657 => 32756,
    16658 => 32756,
    16659 => 32756,
    16660 => 32756,
    16661 => 32755,
    16662 => 32755,
    16663 => 32755,
    16664 => 32755,
    16665 => 32755,
    16666 => 32755,
    16667 => 32755,
    16668 => 32755,
    16669 => 32755,
    16670 => 32755,
    16671 => 32755,
    16672 => 32755,
    16673 => 32754,
    16674 => 32754,
    16675 => 32754,
    16676 => 32754,
    16677 => 32754,
    16678 => 32754,
    16679 => 32754,
    16680 => 32754,
    16681 => 32754,
    16682 => 32754,
    16683 => 32754,
    16684 => 32753,
    16685 => 32753,
    16686 => 32753,
    16687 => 32753,
    16688 => 32753,
    16689 => 32753,
    16690 => 32753,
    16691 => 32753,
    16692 => 32753,
    16693 => 32753,
    16694 => 32753,
    16695 => 32752,
    16696 => 32752,
    16697 => 32752,
    16698 => 32752,
    16699 => 32752,
    16700 => 32752,
    16701 => 32752,
    16702 => 32752,
    16703 => 32752,
    16704 => 32752,
    16705 => 32751,
    16706 => 32751,
    16707 => 32751,
    16708 => 32751,
    16709 => 32751,
    16710 => 32751,
    16711 => 32751,
    16712 => 32751,
    16713 => 32751,
    16714 => 32751,
    16715 => 32751,
    16716 => 32750,
    16717 => 32750,
    16718 => 32750,
    16719 => 32750,
    16720 => 32750,
    16721 => 32750,
    16722 => 32750,
    16723 => 32750,
    16724 => 32750,
    16725 => 32749,
    16726 => 32749,
    16727 => 32749,
    16728 => 32749,
    16729 => 32749,
    16730 => 32749,
    16731 => 32749,
    16732 => 32749,
    16733 => 32749,
    16734 => 32749,
    16735 => 32748,
    16736 => 32748,
    16737 => 32748,
    16738 => 32748,
    16739 => 32748,
    16740 => 32748,
    16741 => 32748,
    16742 => 32748,
    16743 => 32748,
    16744 => 32747,
    16745 => 32747,
    16746 => 32747,
    16747 => 32747,
    16748 => 32747,
    16749 => 32747,
    16750 => 32747,
    16751 => 32747,
    16752 => 32747,
    16753 => 32746,
    16754 => 32746,
    16755 => 32746,
    16756 => 32746,
    16757 => 32746,
    16758 => 32746,
    16759 => 32746,
    16760 => 32746,
    16761 => 32746,
    16762 => 32745,
    16763 => 32745,
    16764 => 32745,
    16765 => 32745,
    16766 => 32745,
    16767 => 32745,
    16768 => 32745,
    16769 => 32745,
    16770 => 32745,
    16771 => 32744,
    16772 => 32744,
    16773 => 32744,
    16774 => 32744,
    16775 => 32744,
    16776 => 32744,
    16777 => 32744,
    16778 => 32744,
    16779 => 32744,
    16780 => 32743,
    16781 => 32743,
    16782 => 32743,
    16783 => 32743,
    16784 => 32743,
    16785 => 32743,
    16786 => 32743,
    16787 => 32743,
    16788 => 32742,
    16789 => 32742,
    16790 => 32742,
    16791 => 32742,
    16792 => 32742,
    16793 => 32742,
    16794 => 32742,
    16795 => 32742,
    16796 => 32741,
    16797 => 32741,
    16798 => 32741,
    16799 => 32741,
    16800 => 32741,
    16801 => 32741,
    16802 => 32741,
    16803 => 32741,
    16804 => 32740,
    16805 => 32740,
    16806 => 32740,
    16807 => 32740,
    16808 => 32740,
    16809 => 32740,
    16810 => 32740,
    16811 => 32740,
    16812 => 32739,
    16813 => 32739,
    16814 => 32739,
    16815 => 32739,
    16816 => 32739,
    16817 => 32739,
    16818 => 32739,
    16819 => 32739,
    16820 => 32738,
    16821 => 32738,
    16822 => 32738,
    16823 => 32738,
    16824 => 32738,
    16825 => 32738,
    16826 => 32738,
    16827 => 32737,
    16828 => 32737,
    16829 => 32737,
    16830 => 32737,
    16831 => 32737,
    16832 => 32737,
    16833 => 32737,
    16834 => 32737,
    16835 => 32736,
    16836 => 32736,
    16837 => 32736,
    16838 => 32736,
    16839 => 32736,
    16840 => 32736,
    16841 => 32736,
    16842 => 32735,
    16843 => 32735,
    16844 => 32735,
    16845 => 32735,
    16846 => 32735,
    16847 => 32735,
    16848 => 32735,
    16849 => 32734,
    16850 => 32734,
    16851 => 32734,
    16852 => 32734,
    16853 => 32734,
    16854 => 32734,
    16855 => 32734,
    16856 => 32733,
    16857 => 32733,
    16858 => 32733,
    16859 => 32733,
    16860 => 32733,
    16861 => 32733,
    16862 => 32733,
    16863 => 32732,
    16864 => 32732,
    16865 => 32732,
    16866 => 32732,
    16867 => 32732,
    16868 => 32732,
    16869 => 32732,
    16870 => 32731,
    16871 => 32731,
    16872 => 32731,
    16873 => 32731,
    16874 => 32731,
    16875 => 32731,
    16876 => 32731,
    16877 => 32730,
    16878 => 32730,
    16879 => 32730,
    16880 => 32730,
    16881 => 32730,
    16882 => 32730,
    16883 => 32730,
    16884 => 32729,
    16885 => 32729,
    16886 => 32729,
    16887 => 32729,
    16888 => 32729,
    16889 => 32729,
    16890 => 32728,
    16891 => 32728,
    16892 => 32728,
    16893 => 32728,
    16894 => 32728,
    16895 => 32728,
    16896 => 32728,
    16897 => 32727,
    16898 => 32727,
    16899 => 32727,
    16900 => 32727,
    16901 => 32727,
    16902 => 32727,
    16903 => 32726,
    16904 => 32726,
    16905 => 32726,
    16906 => 32726,
    16907 => 32726,
    16908 => 32726,
    16909 => 32726,
    16910 => 32725,
    16911 => 32725,
    16912 => 32725,
    16913 => 32725,
    16914 => 32725,
    16915 => 32725,
    16916 => 32724,
    16917 => 32724,
    16918 => 32724,
    16919 => 32724,
    16920 => 32724,
    16921 => 32724,
    16922 => 32723,
    16923 => 32723,
    16924 => 32723,
    16925 => 32723,
    16926 => 32723,
    16927 => 32723,
    16928 => 32722,
    16929 => 32722,
    16930 => 32722,
    16931 => 32722,
    16932 => 32722,
    16933 => 32722,
    16934 => 32721,
    16935 => 32721,
    16936 => 32721,
    16937 => 32721,
    16938 => 32721,
    16939 => 32721,
    16940 => 32720,
    16941 => 32720,
    16942 => 32720,
    16943 => 32720,
    16944 => 32720,
    16945 => 32720,
    16946 => 32719,
    16947 => 32719,
    16948 => 32719,
    16949 => 32719,
    16950 => 32719,
    16951 => 32719,
    16952 => 32718,
    16953 => 32718,
    16954 => 32718,
    16955 => 32718,
    16956 => 32718,
    16957 => 32718,
    16958 => 32717,
    16959 => 32717,
    16960 => 32717,
    16961 => 32717,
    16962 => 32717,
    16963 => 32717,
    16964 => 32716,
    16965 => 32716,
    16966 => 32716,
    16967 => 32716,
    16968 => 32716,
    16969 => 32715,
    16970 => 32715,
    16971 => 32715,
    16972 => 32715,
    16973 => 32715,
    16974 => 32715,
    16975 => 32714,
    16976 => 32714,
    16977 => 32714,
    16978 => 32714,
    16979 => 32714,
    16980 => 32714,
    16981 => 32713,
    16982 => 32713,
    16983 => 32713,
    16984 => 32713,
    16985 => 32713,
    16986 => 32712,
    16987 => 32712,
    16988 => 32712,
    16989 => 32712,
    16990 => 32712,
    16991 => 32712,
    16992 => 32711,
    16993 => 32711,
    16994 => 32711,
    16995 => 32711,
    16996 => 32711,
    16997 => 32710,
    16998 => 32710,
    16999 => 32710,
    17000 => 32710,
    17001 => 32710,
    17002 => 32710,
    17003 => 32709,
    17004 => 32709,
    17005 => 32709,
    17006 => 32709,
    17007 => 32709,
    17008 => 32708,
    17009 => 32708,
    17010 => 32708,
    17011 => 32708,
    17012 => 32708,
    17013 => 32707,
    17014 => 32707,
    17015 => 32707,
    17016 => 32707,
    17017 => 32707,
    17018 => 32706,
    17019 => 32706,
    17020 => 32706,
    17021 => 32706,
    17022 => 32706,
    17023 => 32706,
    17024 => 32705,
    17025 => 32705,
    17026 => 32705,
    17027 => 32705,
    17028 => 32705,
    17029 => 32704,
    17030 => 32704,
    17031 => 32704,
    17032 => 32704,
    17033 => 32704,
    17034 => 32703,
    17035 => 32703,
    17036 => 32703,
    17037 => 32703,
    17038 => 32703,
    17039 => 32702,
    17040 => 32702,
    17041 => 32702,
    17042 => 32702,
    17043 => 32702,
    17044 => 32701,
    17045 => 32701,
    17046 => 32701,
    17047 => 32701,
    17048 => 32701,
    17049 => 32700,
    17050 => 32700,
    17051 => 32700,
    17052 => 32700,
    17053 => 32700,
    17054 => 32699,
    17055 => 32699,
    17056 => 32699,
    17057 => 32699,
    17058 => 32699,
    17059 => 32698,
    17060 => 32698,
    17061 => 32698,
    17062 => 32698,
    17063 => 32698,
    17064 => 32697,
    17065 => 32697,
    17066 => 32697,
    17067 => 32697,
    17068 => 32697,
    17069 => 32696,
    17070 => 32696,
    17071 => 32696,
    17072 => 32696,
    17073 => 32696,
    17074 => 32695,
    17075 => 32695,
    17076 => 32695,
    17077 => 32695,
    17078 => 32694,
    17079 => 32694,
    17080 => 32694,
    17081 => 32694,
    17082 => 32694,
    17083 => 32693,
    17084 => 32693,
    17085 => 32693,
    17086 => 32693,
    17087 => 32693,
    17088 => 32692,
    17089 => 32692,
    17090 => 32692,
    17091 => 32692,
    17092 => 32692,
    17093 => 32691,
    17094 => 32691,
    17095 => 32691,
    17096 => 32691,
    17097 => 32690,
    17098 => 32690,
    17099 => 32690,
    17100 => 32690,
    17101 => 32690,
    17102 => 32689,
    17103 => 32689,
    17104 => 32689,
    17105 => 32689,
    17106 => 32689,
    17107 => 32688,
    17108 => 32688,
    17109 => 32688,
    17110 => 32688,
    17111 => 32687,
    17112 => 32687,
    17113 => 32687,
    17114 => 32687,
    17115 => 32687,
    17116 => 32686,
    17117 => 32686,
    17118 => 32686,
    17119 => 32686,
    17120 => 32685,
    17121 => 32685,
    17122 => 32685,
    17123 => 32685,
    17124 => 32685,
    17125 => 32684,
    17126 => 32684,
    17127 => 32684,
    17128 => 32684,
    17129 => 32683,
    17130 => 32683,
    17131 => 32683,
    17132 => 32683,
    17133 => 32683,
    17134 => 32682,
    17135 => 32682,
    17136 => 32682,
    17137 => 32682,
    17138 => 32681,
    17139 => 32681,
    17140 => 32681,
    17141 => 32681,
    17142 => 32681,
    17143 => 32680,
    17144 => 32680,
    17145 => 32680,
    17146 => 32680,
    17147 => 32679,
    17148 => 32679,
    17149 => 32679,
    17150 => 32679,
    17151 => 32678,
    17152 => 32678,
    17153 => 32678,
    17154 => 32678,
    17155 => 32678,
    17156 => 32677,
    17157 => 32677,
    17158 => 32677,
    17159 => 32677,
    17160 => 32676,
    17161 => 32676,
    17162 => 32676,
    17163 => 32676,
    17164 => 32675,
    17165 => 32675,
    17166 => 32675,
    17167 => 32675,
    17168 => 32674,
    17169 => 32674,
    17170 => 32674,
    17171 => 32674,
    17172 => 32674,
    17173 => 32673,
    17174 => 32673,
    17175 => 32673,
    17176 => 32673,
    17177 => 32672,
    17178 => 32672,
    17179 => 32672,
    17180 => 32672,
    17181 => 32671,
    17182 => 32671,
    17183 => 32671,
    17184 => 32671,
    17185 => 32670,
    17186 => 32670,
    17187 => 32670,
    17188 => 32670,
    17189 => 32669,
    17190 => 32669,
    17191 => 32669,
    17192 => 32669,
    17193 => 32668,
    17194 => 32668,
    17195 => 32668,
    17196 => 32668,
    17197 => 32668,
    17198 => 32667,
    17199 => 32667,
    17200 => 32667,
    17201 => 32667,
    17202 => 32666,
    17203 => 32666,
    17204 => 32666,
    17205 => 32666,
    17206 => 32665,
    17207 => 32665,
    17208 => 32665,
    17209 => 32665,
    17210 => 32664,
    17211 => 32664,
    17212 => 32664,
    17213 => 32664,
    17214 => 32663,
    17215 => 32663,
    17216 => 32663,
    17217 => 32663,
    17218 => 32662,
    17219 => 32662,
    17220 => 32662,
    17221 => 32662,
    17222 => 32661,
    17223 => 32661,
    17224 => 32661,
    17225 => 32661,
    17226 => 32660,
    17227 => 32660,
    17228 => 32660,
    17229 => 32660,
    17230 => 32659,
    17231 => 32659,
    17232 => 32659,
    17233 => 32659,
    17234 => 32658,
    17235 => 32658,
    17236 => 32658,
    17237 => 32657,
    17238 => 32657,
    17239 => 32657,
    17240 => 32657,
    17241 => 32656,
    17242 => 32656,
    17243 => 32656,
    17244 => 32656,
    17245 => 32655,
    17246 => 32655,
    17247 => 32655,
    17248 => 32655,
    17249 => 32654,
    17250 => 32654,
    17251 => 32654,
    17252 => 32654,
    17253 => 32653,
    17254 => 32653,
    17255 => 32653,
    17256 => 32653,
    17257 => 32652,
    17258 => 32652,
    17259 => 32652,
    17260 => 32652,
    17261 => 32651,
    17262 => 32651,
    17263 => 32651,
    17264 => 32650,
    17265 => 32650,
    17266 => 32650,
    17267 => 32650,
    17268 => 32649,
    17269 => 32649,
    17270 => 32649,
    17271 => 32649,
    17272 => 32648,
    17273 => 32648,
    17274 => 32648,
    17275 => 32648,
    17276 => 32647,
    17277 => 32647,
    17278 => 32647,
    17279 => 32646,
    17280 => 32646,
    17281 => 32646,
    17282 => 32646,
    17283 => 32645,
    17284 => 32645,
    17285 => 32645,
    17286 => 32645,
    17287 => 32644,
    17288 => 32644,
    17289 => 32644,
    17290 => 32643,
    17291 => 32643,
    17292 => 32643,
    17293 => 32643,
    17294 => 32642,
    17295 => 32642,
    17296 => 32642,
    17297 => 32642,
    17298 => 32641,
    17299 => 32641,
    17300 => 32641,
    17301 => 32640,
    17302 => 32640,
    17303 => 32640,
    17304 => 32640,
    17305 => 32639,
    17306 => 32639,
    17307 => 32639,
    17308 => 32639,
    17309 => 32638,
    17310 => 32638,
    17311 => 32638,
    17312 => 32637,
    17313 => 32637,
    17314 => 32637,
    17315 => 32637,
    17316 => 32636,
    17317 => 32636,
    17318 => 32636,
    17319 => 32635,
    17320 => 32635,
    17321 => 32635,
    17322 => 32635,
    17323 => 32634,
    17324 => 32634,
    17325 => 32634,
    17326 => 32633,
    17327 => 32633,
    17328 => 32633,
    17329 => 32633,
    17330 => 32632,
    17331 => 32632,
    17332 => 32632,
    17333 => 32631,
    17334 => 32631,
    17335 => 32631,
    17336 => 32631,
    17337 => 32630,
    17338 => 32630,
    17339 => 32630,
    17340 => 32629,
    17341 => 32629,
    17342 => 32629,
    17343 => 32629,
    17344 => 32628,
    17345 => 32628,
    17346 => 32628,
    17347 => 32627,
    17348 => 32627,
    17349 => 32627,
    17350 => 32627,
    17351 => 32626,
    17352 => 32626,
    17353 => 32626,
    17354 => 32625,
    17355 => 32625,
    17356 => 32625,
    17357 => 32625,
    17358 => 32624,
    17359 => 32624,
    17360 => 32624,
    17361 => 32623,
    17362 => 32623,
    17363 => 32623,
    17364 => 32622,
    17365 => 32622,
    17366 => 32622,
    17367 => 32622,
    17368 => 32621,
    17369 => 32621,
    17370 => 32621,
    17371 => 32620,
    17372 => 32620,
    17373 => 32620,
    17374 => 32620,
    17375 => 32619,
    17376 => 32619,
    17377 => 32619,
    17378 => 32618,
    17379 => 32618,
    17380 => 32618,
    17381 => 32617,
    17382 => 32617,
    17383 => 32617,
    17384 => 32617,
    17385 => 32616,
    17386 => 32616,
    17387 => 32616,
    17388 => 32615,
    17389 => 32615,
    17390 => 32615,
    17391 => 32614,
    17392 => 32614,
    17393 => 32614,
    17394 => 32613,
    17395 => 32613,
    17396 => 32613,
    17397 => 32613,
    17398 => 32612,
    17399 => 32612,
    17400 => 32612,
    17401 => 32611,
    17402 => 32611,
    17403 => 32611,
    17404 => 32610,
    17405 => 32610,
    17406 => 32610,
    17407 => 32610,
    17408 => 32609,
    17409 => 32609,
    17410 => 32609,
    17411 => 32608,
    17412 => 32608,
    17413 => 32608,
    17414 => 32607,
    17415 => 32607,
    17416 => 32607,
    17417 => 32606,
    17418 => 32606,
    17419 => 32606,
    17420 => 32606,
    17421 => 32605,
    17422 => 32605,
    17423 => 32605,
    17424 => 32604,
    17425 => 32604,
    17426 => 32604,
    17427 => 32603,
    17428 => 32603,
    17429 => 32603,
    17430 => 32602,
    17431 => 32602,
    17432 => 32602,
    17433 => 32601,
    17434 => 32601,
    17435 => 32601,
    17436 => 32600,
    17437 => 32600,
    17438 => 32600,
    17439 => 32600,
    17440 => 32599,
    17441 => 32599,
    17442 => 32599,
    17443 => 32598,
    17444 => 32598,
    17445 => 32598,
    17446 => 32597,
    17447 => 32597,
    17448 => 32597,
    17449 => 32596,
    17450 => 32596,
    17451 => 32596,
    17452 => 32595,
    17453 => 32595,
    17454 => 32595,
    17455 => 32594,
    17456 => 32594,
    17457 => 32594,
    17458 => 32593,
    17459 => 32593,
    17460 => 32593,
    17461 => 32592,
    17462 => 32592,
    17463 => 32592,
    17464 => 32592,
    17465 => 32591,
    17466 => 32591,
    17467 => 32591,
    17468 => 32590,
    17469 => 32590,
    17470 => 32590,
    17471 => 32589,
    17472 => 32589,
    17473 => 32589,
    17474 => 32588,
    17475 => 32588,
    17476 => 32588,
    17477 => 32587,
    17478 => 32587,
    17479 => 32587,
    17480 => 32586,
    17481 => 32586,
    17482 => 32586,
    17483 => 32585,
    17484 => 32585,
    17485 => 32585,
    17486 => 32584,
    17487 => 32584,
    17488 => 32584,
    17489 => 32583,
    17490 => 32583,
    17491 => 32583,
    17492 => 32582,
    17493 => 32582,
    17494 => 32582,
    17495 => 32581,
    17496 => 32581,
    17497 => 32581,
    17498 => 32580,
    17499 => 32580,
    17500 => 32580,
    17501 => 32579,
    17502 => 32579,
    17503 => 32579,
    17504 => 32578,
    17505 => 32578,
    17506 => 32578,
    17507 => 32577,
    17508 => 32577,
    17509 => 32577,
    17510 => 32576,
    17511 => 32576,
    17512 => 32576,
    17513 => 32575,
    17514 => 32575,
    17515 => 32575,
    17516 => 32574,
    17517 => 32574,
    17518 => 32574,
    17519 => 32573,
    17520 => 32573,
    17521 => 32573,
    17522 => 32572,
    17523 => 32572,
    17524 => 32571,
    17525 => 32571,
    17526 => 32571,
    17527 => 32570,
    17528 => 32570,
    17529 => 32570,
    17530 => 32569,
    17531 => 32569,
    17532 => 32569,
    17533 => 32568,
    17534 => 32568,
    17535 => 32568,
    17536 => 32567,
    17537 => 32567,
    17538 => 32567,
    17539 => 32566,
    17540 => 32566,
    17541 => 32566,
    17542 => 32565,
    17543 => 32565,
    17544 => 32565,
    17545 => 32564,
    17546 => 32564,
    17547 => 32564,
    17548 => 32563,
    17549 => 32563,
    17550 => 32562,
    17551 => 32562,
    17552 => 32562,
    17553 => 32561,
    17554 => 32561,
    17555 => 32561,
    17556 => 32560,
    17557 => 32560,
    17558 => 32560,
    17559 => 32559,
    17560 => 32559,
    17561 => 32559,
    17562 => 32558,
    17563 => 32558,
    17564 => 32558,
    17565 => 32557,
    17566 => 32557,
    17567 => 32556,
    17568 => 32556,
    17569 => 32556,
    17570 => 32555,
    17571 => 32555,
    17572 => 32555,
    17573 => 32554,
    17574 => 32554,
    17575 => 32554,
    17576 => 32553,
    17577 => 32553,
    17578 => 32553,
    17579 => 32552,
    17580 => 32552,
    17581 => 32551,
    17582 => 32551,
    17583 => 32551,
    17584 => 32550,
    17585 => 32550,
    17586 => 32550,
    17587 => 32549,
    17588 => 32549,
    17589 => 32549,
    17590 => 32548,
    17591 => 32548,
    17592 => 32547,
    17593 => 32547,
    17594 => 32547,
    17595 => 32546,
    17596 => 32546,
    17597 => 32546,
    17598 => 32545,
    17599 => 32545,
    17600 => 32545,
    17601 => 32544,
    17602 => 32544,
    17603 => 32543,
    17604 => 32543,
    17605 => 32543,
    17606 => 32542,
    17607 => 32542,
    17608 => 32542,
    17609 => 32541,
    17610 => 32541,
    17611 => 32541,
    17612 => 32540,
    17613 => 32540,
    17614 => 32539,
    17615 => 32539,
    17616 => 32539,
    17617 => 32538,
    17618 => 32538,
    17619 => 32538,
    17620 => 32537,
    17621 => 32537,
    17622 => 32536,
    17623 => 32536,
    17624 => 32536,
    17625 => 32535,
    17626 => 32535,
    17627 => 32535,
    17628 => 32534,
    17629 => 32534,
    17630 => 32533,
    17631 => 32533,
    17632 => 32533,
    17633 => 32532,
    17634 => 32532,
    17635 => 32532,
    17636 => 32531,
    17637 => 32531,
    17638 => 32530,
    17639 => 32530,
    17640 => 32530,
    17641 => 32529,
    17642 => 32529,
    17643 => 32529,
    17644 => 32528,
    17645 => 32528,
    17646 => 32527,
    17647 => 32527,
    17648 => 32527,
    17649 => 32526,
    17650 => 32526,
    17651 => 32526,
    17652 => 32525,
    17653 => 32525,
    17654 => 32524,
    17655 => 32524,
    17656 => 32524,
    17657 => 32523,
    17658 => 32523,
    17659 => 32522,
    17660 => 32522,
    17661 => 32522,
    17662 => 32521,
    17663 => 32521,
    17664 => 32521,
    17665 => 32520,
    17666 => 32520,
    17667 => 32519,
    17668 => 32519,
    17669 => 32519,
    17670 => 32518,
    17671 => 32518,
    17672 => 32517,
    17673 => 32517,
    17674 => 32517,
    17675 => 32516,
    17676 => 32516,
    17677 => 32516,
    17678 => 32515,
    17679 => 32515,
    17680 => 32514,
    17681 => 32514,
    17682 => 32514,
    17683 => 32513,
    17684 => 32513,
    17685 => 32512,
    17686 => 32512,
    17687 => 32512,
    17688 => 32511,
    17689 => 32511,
    17690 => 32510,
    17691 => 32510,
    17692 => 32510,
    17693 => 32509,
    17694 => 32509,
    17695 => 32509,
    17696 => 32508,
    17697 => 32508,
    17698 => 32507,
    17699 => 32507,
    17700 => 32507,
    17701 => 32506,
    17702 => 32506,
    17703 => 32505,
    17704 => 32505,
    17705 => 32505,
    17706 => 32504,
    17707 => 32504,
    17708 => 32503,
    17709 => 32503,
    17710 => 32503,
    17711 => 32502,
    17712 => 32502,
    17713 => 32501,
    17714 => 32501,
    17715 => 32501,
    17716 => 32500,
    17717 => 32500,
    17718 => 32499,
    17719 => 32499,
    17720 => 32499,
    17721 => 32498,
    17722 => 32498,
    17723 => 32497,
    17724 => 32497,
    17725 => 32497,
    17726 => 32496,
    17727 => 32496,
    17728 => 32495,
    17729 => 32495,
    17730 => 32495,
    17731 => 32494,
    17732 => 32494,
    17733 => 32493,
    17734 => 32493,
    17735 => 32493,
    17736 => 32492,
    17737 => 32492,
    17738 => 32491,
    17739 => 32491,
    17740 => 32490,
    17741 => 32490,
    17742 => 32490,
    17743 => 32489,
    17744 => 32489,
    17745 => 32488,
    17746 => 32488,
    17747 => 32488,
    17748 => 32487,
    17749 => 32487,
    17750 => 32486,
    17751 => 32486,
    17752 => 32486,
    17753 => 32485,
    17754 => 32485,
    17755 => 32484,
    17756 => 32484,
    17757 => 32484,
    17758 => 32483,
    17759 => 32483,
    17760 => 32482,
    17761 => 32482,
    17762 => 32481,
    17763 => 32481,
    17764 => 32481,
    17765 => 32480,
    17766 => 32480,
    17767 => 32479,
    17768 => 32479,
    17769 => 32479,
    17770 => 32478,
    17771 => 32478,
    17772 => 32477,
    17773 => 32477,
    17774 => 32476,
    17775 => 32476,
    17776 => 32476,
    17777 => 32475,
    17778 => 32475,
    17779 => 32474,
    17780 => 32474,
    17781 => 32474,
    17782 => 32473,
    17783 => 32473,
    17784 => 32472,
    17785 => 32472,
    17786 => 32471,
    17787 => 32471,
    17788 => 32471,
    17789 => 32470,
    17790 => 32470,
    17791 => 32469,
    17792 => 32469,
    17793 => 32468,
    17794 => 32468,
    17795 => 32468,
    17796 => 32467,
    17797 => 32467,
    17798 => 32466,
    17799 => 32466,
    17800 => 32466,
    17801 => 32465,
    17802 => 32465,
    17803 => 32464,
    17804 => 32464,
    17805 => 32463,
    17806 => 32463,
    17807 => 32463,
    17808 => 32462,
    17809 => 32462,
    17810 => 32461,
    17811 => 32461,
    17812 => 32460,
    17813 => 32460,
    17814 => 32460,
    17815 => 32459,
    17816 => 32459,
    17817 => 32458,
    17818 => 32458,
    17819 => 32457,
    17820 => 32457,
    17821 => 32457,
    17822 => 32456,
    17823 => 32456,
    17824 => 32455,
    17825 => 32455,
    17826 => 32454,
    17827 => 32454,
    17828 => 32453,
    17829 => 32453,
    17830 => 32453,
    17831 => 32452,
    17832 => 32452,
    17833 => 32451,
    17834 => 32451,
    17835 => 32450,
    17836 => 32450,
    17837 => 32450,
    17838 => 32449,
    17839 => 32449,
    17840 => 32448,
    17841 => 32448,
    17842 => 32447,
    17843 => 32447,
    17844 => 32447,
    17845 => 32446,
    17846 => 32446,
    17847 => 32445,
    17848 => 32445,
    17849 => 32444,
    17850 => 32444,
    17851 => 32443,
    17852 => 32443,
    17853 => 32443,
    17854 => 32442,
    17855 => 32442,
    17856 => 32441,
    17857 => 32441,
    17858 => 32440,
    17859 => 32440,
    17860 => 32439,
    17861 => 32439,
    17862 => 32439,
    17863 => 32438,
    17864 => 32438,
    17865 => 32437,
    17866 => 32437,
    17867 => 32436,
    17868 => 32436,
    17869 => 32435,
    17870 => 32435,
    17871 => 32435,
    17872 => 32434,
    17873 => 32434,
    17874 => 32433,
    17875 => 32433,
    17876 => 32432,
    17877 => 32432,
    17878 => 32431,
    17879 => 32431,
    17880 => 32431,
    17881 => 32430,
    17882 => 32430,
    17883 => 32429,
    17884 => 32429,
    17885 => 32428,
    17886 => 32428,
    17887 => 32427,
    17888 => 32427,
    17889 => 32426,
    17890 => 32426,
    17891 => 32426,
    17892 => 32425,
    17893 => 32425,
    17894 => 32424,
    17895 => 32424,
    17896 => 32423,
    17897 => 32423,
    17898 => 32422,
    17899 => 32422,
    17900 => 32422,
    17901 => 32421,
    17902 => 32421,
    17903 => 32420,
    17904 => 32420,
    17905 => 32419,
    17906 => 32419,
    17907 => 32418,
    17908 => 32418,
    17909 => 32417,
    17910 => 32417,
    17911 => 32416,
    17912 => 32416,
    17913 => 32416,
    17914 => 32415,
    17915 => 32415,
    17916 => 32414,
    17917 => 32414,
    17918 => 32413,
    17919 => 32413,
    17920 => 32412,
    17921 => 32412,
    17922 => 32411,
    17923 => 32411,
    17924 => 32411,
    17925 => 32410,
    17926 => 32410,
    17927 => 32409,
    17928 => 32409,
    17929 => 32408,
    17930 => 32408,
    17931 => 32407,
    17932 => 32407,
    17933 => 32406,
    17934 => 32406,
    17935 => 32405,
    17936 => 32405,
    17937 => 32404,
    17938 => 32404,
    17939 => 32404,
    17940 => 32403,
    17941 => 32403,
    17942 => 32402,
    17943 => 32402,
    17944 => 32401,
    17945 => 32401,
    17946 => 32400,
    17947 => 32400,
    17948 => 32399,
    17949 => 32399,
    17950 => 32398,
    17951 => 32398,
    17952 => 32397,
    17953 => 32397,
    17954 => 32397,
    17955 => 32396,
    17956 => 32396,
    17957 => 32395,
    17958 => 32395,
    17959 => 32394,
    17960 => 32394,
    17961 => 32393,
    17962 => 32393,
    17963 => 32392,
    17964 => 32392,
    17965 => 32391,
    17966 => 32391,
    17967 => 32390,
    17968 => 32390,
    17969 => 32389,
    17970 => 32389,
    17971 => 32388,
    17972 => 32388,
    17973 => 32387,
    17974 => 32387,
    17975 => 32387,
    17976 => 32386,
    17977 => 32386,
    17978 => 32385,
    17979 => 32385,
    17980 => 32384,
    17981 => 32384,
    17982 => 32383,
    17983 => 32383,
    17984 => 32382,
    17985 => 32382,
    17986 => 32381,
    17987 => 32381,
    17988 => 32380,
    17989 => 32380,
    17990 => 32379,
    17991 => 32379,
    17992 => 32378,
    17993 => 32378,
    17994 => 32377,
    17995 => 32377,
    17996 => 32376,
    17997 => 32376,
    17998 => 32375,
    17999 => 32375,
    18000 => 32375,
    18001 => 32374,
    18002 => 32374,
    18003 => 32373,
    18004 => 32373,
    18005 => 32372,
    18006 => 32372,
    18007 => 32371,
    18008 => 32371,
    18009 => 32370,
    18010 => 32370,
    18011 => 32369,
    18012 => 32369,
    18013 => 32368,
    18014 => 32368,
    18015 => 32367,
    18016 => 32367,
    18017 => 32366,
    18018 => 32366,
    18019 => 32365,
    18020 => 32365,
    18021 => 32364,
    18022 => 32364,
    18023 => 32363,
    18024 => 32363,
    18025 => 32362,
    18026 => 32362,
    18027 => 32361,
    18028 => 32361,
    18029 => 32360,
    18030 => 32360,
    18031 => 32359,
    18032 => 32359,
    18033 => 32358,
    18034 => 32358,
    18035 => 32357,
    18036 => 32357,
    18037 => 32356,
    18038 => 32356,
    18039 => 32355,
    18040 => 32355,
    18041 => 32354,
    18042 => 32354,
    18043 => 32353,
    18044 => 32353,
    18045 => 32352,
    18046 => 32352,
    18047 => 32351,
    18048 => 32351,
    18049 => 32350,
    18050 => 32350,
    18051 => 32349,
    18052 => 32349,
    18053 => 32348,
    18054 => 32348,
    18055 => 32347,
    18056 => 32347,
    18057 => 32346,
    18058 => 32346,
    18059 => 32345,
    18060 => 32345,
    18061 => 32344,
    18062 => 32344,
    18063 => 32343,
    18064 => 32343,
    18065 => 32342,
    18066 => 32342,
    18067 => 32341,
    18068 => 32341,
    18069 => 32340,
    18070 => 32340,
    18071 => 32339,
    18072 => 32339,
    18073 => 32338,
    18074 => 32338,
    18075 => 32337,
    18076 => 32337,
    18077 => 32336,
    18078 => 32336,
    18079 => 32335,
    18080 => 32335,
    18081 => 32334,
    18082 => 32334,
    18083 => 32333,
    18084 => 32333,
    18085 => 32332,
    18086 => 32332,
    18087 => 32331,
    18088 => 32331,
    18089 => 32330,
    18090 => 32330,
    18091 => 32329,
    18092 => 32329,
    18093 => 32328,
    18094 => 32328,
    18095 => 32327,
    18096 => 32327,
    18097 => 32326,
    18098 => 32326,
    18099 => 32325,
    18100 => 32325,
    18101 => 32324,
    18102 => 32324,
    18103 => 32323,
    18104 => 32322,
    18105 => 32322,
    18106 => 32321,
    18107 => 32321,
    18108 => 32320,
    18109 => 32320,
    18110 => 32319,
    18111 => 32319,
    18112 => 32318,
    18113 => 32318,
    18114 => 32317,
    18115 => 32317,
    18116 => 32316,
    18117 => 32316,
    18118 => 32315,
    18119 => 32315,
    18120 => 32314,
    18121 => 32314,
    18122 => 32313,
    18123 => 32313,
    18124 => 32312,
    18125 => 32312,
    18126 => 32311,
    18127 => 32311,
    18128 => 32310,
    18129 => 32310,
    18130 => 32309,
    18131 => 32308,
    18132 => 32308,
    18133 => 32307,
    18134 => 32307,
    18135 => 32306,
    18136 => 32306,
    18137 => 32305,
    18138 => 32305,
    18139 => 32304,
    18140 => 32304,
    18141 => 32303,
    18142 => 32303,
    18143 => 32302,
    18144 => 32302,
    18145 => 32301,
    18146 => 32301,
    18147 => 32300,
    18148 => 32300,
    18149 => 32299,
    18150 => 32298,
    18151 => 32298,
    18152 => 32297,
    18153 => 32297,
    18154 => 32296,
    18155 => 32296,
    18156 => 32295,
    18157 => 32295,
    18158 => 32294,
    18159 => 32294,
    18160 => 32293,
    18161 => 32293,
    18162 => 32292,
    18163 => 32292,
    18164 => 32291,
    18165 => 32290,
    18166 => 32290,
    18167 => 32289,
    18168 => 32289,
    18169 => 32288,
    18170 => 32288,
    18171 => 32287,
    18172 => 32287,
    18173 => 32286,
    18174 => 32286,
    18175 => 32285,
    18176 => 32285,
    18177 => 32284,
    18178 => 32284,
    18179 => 32283,
    18180 => 32282,
    18181 => 32282,
    18182 => 32281,
    18183 => 32281,
    18184 => 32280,
    18185 => 32280,
    18186 => 32279,
    18187 => 32279,
    18188 => 32278,
    18189 => 32278,
    18190 => 32277,
    18191 => 32277,
    18192 => 32276,
    18193 => 32275,
    18194 => 32275,
    18195 => 32274,
    18196 => 32274,
    18197 => 32273,
    18198 => 32273,
    18199 => 32272,
    18200 => 32272,
    18201 => 32271,
    18202 => 32271,
    18203 => 32270,
    18204 => 32269,
    18205 => 32269,
    18206 => 32268,
    18207 => 32268,
    18208 => 32267,
    18209 => 32267,
    18210 => 32266,
    18211 => 32266,
    18212 => 32265,
    18213 => 32265,
    18214 => 32264,
    18215 => 32263,
    18216 => 32263,
    18217 => 32262,
    18218 => 32262,
    18219 => 32261,
    18220 => 32261,
    18221 => 32260,
    18222 => 32260,
    18223 => 32259,
    18224 => 32258,
    18225 => 32258,
    18226 => 32257,
    18227 => 32257,
    18228 => 32256,
    18229 => 32256,
    18230 => 32255,
    18231 => 32255,
    18232 => 32254,
    18233 => 32253,
    18234 => 32253,
    18235 => 32252,
    18236 => 32252,
    18237 => 32251,
    18238 => 32251,
    18239 => 32250,
    18240 => 32250,
    18241 => 32249,
    18242 => 32248,
    18243 => 32248,
    18244 => 32247,
    18245 => 32247,
    18246 => 32246,
    18247 => 32246,
    18248 => 32245,
    18249 => 32245,
    18250 => 32244,
    18251 => 32243,
    18252 => 32243,
    18253 => 32242,
    18254 => 32242,
    18255 => 32241,
    18256 => 32241,
    18257 => 32240,
    18258 => 32240,
    18259 => 32239,
    18260 => 32238,
    18261 => 32238,
    18262 => 32237,
    18263 => 32237,
    18264 => 32236,
    18265 => 32236,
    18266 => 32235,
    18267 => 32234,
    18268 => 32234,
    18269 => 32233,
    18270 => 32233,
    18271 => 32232,
    18272 => 32232,
    18273 => 32231,
    18274 => 32231,
    18275 => 32230,
    18276 => 32229,
    18277 => 32229,
    18278 => 32228,
    18279 => 32228,
    18280 => 32227,
    18281 => 32227,
    18282 => 32226,
    18283 => 32225,
    18284 => 32225,
    18285 => 32224,
    18286 => 32224,
    18287 => 32223,
    18288 => 32223,
    18289 => 32222,
    18290 => 32221,
    18291 => 32221,
    18292 => 32220,
    18293 => 32220,
    18294 => 32219,
    18295 => 32219,
    18296 => 32218,
    18297 => 32217,
    18298 => 32217,
    18299 => 32216,
    18300 => 32216,
    18301 => 32215,
    18302 => 32215,
    18303 => 32214,
    18304 => 32213,
    18305 => 32213,
    18306 => 32212,
    18307 => 32212,
    18308 => 32211,
    18309 => 32211,
    18310 => 32210,
    18311 => 32209,
    18312 => 32209,
    18313 => 32208,
    18314 => 32208,
    18315 => 32207,
    18316 => 32206,
    18317 => 32206,
    18318 => 32205,
    18319 => 32205,
    18320 => 32204,
    18321 => 32204,
    18322 => 32203,
    18323 => 32202,
    18324 => 32202,
    18325 => 32201,
    18326 => 32201,
    18327 => 32200,
    18328 => 32200,
    18329 => 32199,
    18330 => 32198,
    18331 => 32198,
    18332 => 32197,
    18333 => 32197,
    18334 => 32196,
    18335 => 32195,
    18336 => 32195,
    18337 => 32194,
    18338 => 32194,
    18339 => 32193,
    18340 => 32193,
    18341 => 32192,
    18342 => 32191,
    18343 => 32191,
    18344 => 32190,
    18345 => 32190,
    18346 => 32189,
    18347 => 32188,
    18348 => 32188,
    18349 => 32187,
    18350 => 32187,
    18351 => 32186,
    18352 => 32185,
    18353 => 32185,
    18354 => 32184,
    18355 => 32184,
    18356 => 32183,
    18357 => 32183,
    18358 => 32182,
    18359 => 32181,
    18360 => 32181,
    18361 => 32180,
    18362 => 32180,
    18363 => 32179,
    18364 => 32178,
    18365 => 32178,
    18366 => 32177,
    18367 => 32177,
    18368 => 32176,
    18369 => 32175,
    18370 => 32175,
    18371 => 32174,
    18372 => 32174,
    18373 => 32173,
    18374 => 32172,
    18375 => 32172,
    18376 => 32171,
    18377 => 32171,
    18378 => 32170,
    18379 => 32169,
    18380 => 32169,
    18381 => 32168,
    18382 => 32168,
    18383 => 32167,
    18384 => 32166,
    18385 => 32166,
    18386 => 32165,
    18387 => 32165,
    18388 => 32164,
    18389 => 32163,
    18390 => 32163,
    18391 => 32162,
    18392 => 32162,
    18393 => 32161,
    18394 => 32160,
    18395 => 32160,
    18396 => 32159,
    18397 => 32159,
    18398 => 32158,
    18399 => 32157,
    18400 => 32157,
    18401 => 32156,
    18402 => 32156,
    18403 => 32155,
    18404 => 32154,
    18405 => 32154,
    18406 => 32153,
    18407 => 32153,
    18408 => 32152,
    18409 => 32151,
    18410 => 32151,
    18411 => 32150,
    18412 => 32150,
    18413 => 32149,
    18414 => 32148,
    18415 => 32148,
    18416 => 32147,
    18417 => 32147,
    18418 => 32146,
    18419 => 32145,
    18420 => 32145,
    18421 => 32144,
    18422 => 32144,
    18423 => 32143,
    18424 => 32142,
    18425 => 32142,
    18426 => 32141,
    18427 => 32140,
    18428 => 32140,
    18429 => 32139,
    18430 => 32139,
    18431 => 32138,
    18432 => 32137,
    18433 => 32137,
    18434 => 32136,
    18435 => 32136,
    18436 => 32135,
    18437 => 32134,
    18438 => 32134,
    18439 => 32133,
    18440 => 32132,
    18441 => 32132,
    18442 => 32131,
    18443 => 32131,
    18444 => 32130,
    18445 => 32129,
    18446 => 32129,
    18447 => 32128,
    18448 => 32128,
    18449 => 32127,
    18450 => 32126,
    18451 => 32126,
    18452 => 32125,
    18453 => 32124,
    18454 => 32124,
    18455 => 32123,
    18456 => 32123,
    18457 => 32122,
    18458 => 32121,
    18459 => 32121,
    18460 => 32120,
    18461 => 32119,
    18462 => 32119,
    18463 => 32118,
    18464 => 32118,
    18465 => 32117,
    18466 => 32116,
    18467 => 32116,
    18468 => 32115,
    18469 => 32115,
    18470 => 32114,
    18471 => 32113,
    18472 => 32113,
    18473 => 32112,
    18474 => 32111,
    18475 => 32111,
    18476 => 32110,
    18477 => 32110,
    18478 => 32109,
    18479 => 32108,
    18480 => 32108,
    18481 => 32107,
    18482 => 32106,
    18483 => 32106,
    18484 => 32105,
    18485 => 32104,
    18486 => 32104,
    18487 => 32103,
    18488 => 32103,
    18489 => 32102,
    18490 => 32101,
    18491 => 32101,
    18492 => 32100,
    18493 => 32099,
    18494 => 32099,
    18495 => 32098,
    18496 => 32098,
    18497 => 32097,
    18498 => 32096,
    18499 => 32096,
    18500 => 32095,
    18501 => 32094,
    18502 => 32094,
    18503 => 32093,
    18504 => 32092,
    18505 => 32092,
    18506 => 32091,
    18507 => 32091,
    18508 => 32090,
    18509 => 32089,
    18510 => 32089,
    18511 => 32088,
    18512 => 32087,
    18513 => 32087,
    18514 => 32086,
    18515 => 32086,
    18516 => 32085,
    18517 => 32084,
    18518 => 32084,
    18519 => 32083,
    18520 => 32082,
    18521 => 32082,
    18522 => 32081,
    18523 => 32080,
    18524 => 32080,
    18525 => 32079,
    18526 => 32078,
    18527 => 32078,
    18528 => 32077,
    18529 => 32077,
    18530 => 32076,
    18531 => 32075,
    18532 => 32075,
    18533 => 32074,
    18534 => 32073,
    18535 => 32073,
    18536 => 32072,
    18537 => 32071,
    18538 => 32071,
    18539 => 32070,
    18540 => 32069,
    18541 => 32069,
    18542 => 32068,
    18543 => 32068,
    18544 => 32067,
    18545 => 32066,
    18546 => 32066,
    18547 => 32065,
    18548 => 32064,
    18549 => 32064,
    18550 => 32063,
    18551 => 32062,
    18552 => 32062,
    18553 => 32061,
    18554 => 32060,
    18555 => 32060,
    18556 => 32059,
    18557 => 32058,
    18558 => 32058,
    18559 => 32057,
    18560 => 32057,
    18561 => 32056,
    18562 => 32055,
    18563 => 32055,
    18564 => 32054,
    18565 => 32053,
    18566 => 32053,
    18567 => 32052,
    18568 => 32051,
    18569 => 32051,
    18570 => 32050,
    18571 => 32049,
    18572 => 32049,
    18573 => 32048,
    18574 => 32047,
    18575 => 32047,
    18576 => 32046,
    18577 => 32045,
    18578 => 32045,
    18579 => 32044,
    18580 => 32043,
    18581 => 32043,
    18582 => 32042,
    18583 => 32041,
    18584 => 32041,
    18585 => 32040,
    18586 => 32040,
    18587 => 32039,
    18588 => 32038,
    18589 => 32038,
    18590 => 32037,
    18591 => 32036,
    18592 => 32036,
    18593 => 32035,
    18594 => 32034,
    18595 => 32034,
    18596 => 32033,
    18597 => 32032,
    18598 => 32032,
    18599 => 32031,
    18600 => 32030,
    18601 => 32030,
    18602 => 32029,
    18603 => 32028,
    18604 => 32028,
    18605 => 32027,
    18606 => 32026,
    18607 => 32026,
    18608 => 32025,
    18609 => 32024,
    18610 => 32024,
    18611 => 32023,
    18612 => 32022,
    18613 => 32022,
    18614 => 32021,
    18615 => 32020,
    18616 => 32020,
    18617 => 32019,
    18618 => 32018,
    18619 => 32018,
    18620 => 32017,
    18621 => 32016,
    18622 => 32016,
    18623 => 32015,
    18624 => 32014,
    18625 => 32014,
    18626 => 32013,
    18627 => 32012,
    18628 => 32012,
    18629 => 32011,
    18630 => 32010,
    18631 => 32010,
    18632 => 32009,
    18633 => 32008,
    18634 => 32008,
    18635 => 32007,
    18636 => 32006,
    18637 => 32006,
    18638 => 32005,
    18639 => 32004,
    18640 => 32004,
    18641 => 32003,
    18642 => 32002,
    18643 => 32002,
    18644 => 32001,
    18645 => 32000,
    18646 => 31999,
    18647 => 31999,
    18648 => 31998,
    18649 => 31997,
    18650 => 31997,
    18651 => 31996,
    18652 => 31995,
    18653 => 31995,
    18654 => 31994,
    18655 => 31993,
    18656 => 31993,
    18657 => 31992,
    18658 => 31991,
    18659 => 31991,
    18660 => 31990,
    18661 => 31989,
    18662 => 31989,
    18663 => 31988,
    18664 => 31987,
    18665 => 31987,
    18666 => 31986,
    18667 => 31985,
    18668 => 31985,
    18669 => 31984,
    18670 => 31983,
    18671 => 31982,
    18672 => 31982,
    18673 => 31981,
    18674 => 31980,
    18675 => 31980,
    18676 => 31979,
    18677 => 31978,
    18678 => 31978,
    18679 => 31977,
    18680 => 31976,
    18681 => 31976,
    18682 => 31975,
    18683 => 31974,
    18684 => 31974,
    18685 => 31973,
    18686 => 31972,
    18687 => 31972,
    18688 => 31971,
    18689 => 31970,
    18690 => 31969,
    18691 => 31969,
    18692 => 31968,
    18693 => 31967,
    18694 => 31967,
    18695 => 31966,
    18696 => 31965,
    18697 => 31965,
    18698 => 31964,
    18699 => 31963,
    18700 => 31963,
    18701 => 31962,
    18702 => 31961,
    18703 => 31960,
    18704 => 31960,
    18705 => 31959,
    18706 => 31958,
    18707 => 31958,
    18708 => 31957,
    18709 => 31956,
    18710 => 31956,
    18711 => 31955,
    18712 => 31954,
    18713 => 31954,
    18714 => 31953,
    18715 => 31952,
    18716 => 31951,
    18717 => 31951,
    18718 => 31950,
    18719 => 31949,
    18720 => 31949,
    18721 => 31948,
    18722 => 31947,
    18723 => 31947,
    18724 => 31946,
    18725 => 31945,
    18726 => 31944,
    18727 => 31944,
    18728 => 31943,
    18729 => 31942,
    18730 => 31942,
    18731 => 31941,
    18732 => 31940,
    18733 => 31940,
    18734 => 31939,
    18735 => 31938,
    18736 => 31937,
    18737 => 31937,
    18738 => 31936,
    18739 => 31935,
    18740 => 31935,
    18741 => 31934,
    18742 => 31933,
    18743 => 31933,
    18744 => 31932,
    18745 => 31931,
    18746 => 31930,
    18747 => 31930,
    18748 => 31929,
    18749 => 31928,
    18750 => 31928,
    18751 => 31927,
    18752 => 31926,
    18753 => 31925,
    18754 => 31925,
    18755 => 31924,
    18756 => 31923,
    18757 => 31923,
    18758 => 31922,
    18759 => 31921,
    18760 => 31921,
    18761 => 31920,
    18762 => 31919,
    18763 => 31918,
    18764 => 31918,
    18765 => 31917,
    18766 => 31916,
    18767 => 31916,
    18768 => 31915,
    18769 => 31914,
    18770 => 31913,
    18771 => 31913,
    18772 => 31912,
    18773 => 31911,
    18774 => 31911,
    18775 => 31910,
    18776 => 31909,
    18777 => 31908,
    18778 => 31908,
    18779 => 31907,
    18780 => 31906,
    18781 => 31906,
    18782 => 31905,
    18783 => 31904,
    18784 => 31903,
    18785 => 31903,
    18786 => 31902,
    18787 => 31901,
    18788 => 31901,
    18789 => 31900,
    18790 => 31899,
    18791 => 31898,
    18792 => 31898,
    18793 => 31897,
    18794 => 31896,
    18795 => 31896,
    18796 => 31895,
    18797 => 31894,
    18798 => 31893,
    18799 => 31893,
    18800 => 31892,
    18801 => 31891,
    18802 => 31890,
    18803 => 31890,
    18804 => 31889,
    18805 => 31888,
    18806 => 31888,
    18807 => 31887,
    18808 => 31886,
    18809 => 31885,
    18810 => 31885,
    18811 => 31884,
    18812 => 31883,
    18813 => 31882,
    18814 => 31882,
    18815 => 31881,
    18816 => 31880,
    18817 => 31880,
    18818 => 31879,
    18819 => 31878,
    18820 => 31877,
    18821 => 31877,
    18822 => 31876,
    18823 => 31875,
    18824 => 31875,
    18825 => 31874,
    18826 => 31873,
    18827 => 31872,
    18828 => 31872,
    18829 => 31871,
    18830 => 31870,
    18831 => 31869,
    18832 => 31869,
    18833 => 31868,
    18834 => 31867,
    18835 => 31866,
    18836 => 31866,
    18837 => 31865,
    18838 => 31864,
    18839 => 31864,
    18840 => 31863,
    18841 => 31862,
    18842 => 31861,
    18843 => 31861,
    18844 => 31860,
    18845 => 31859,
    18846 => 31858,
    18847 => 31858,
    18848 => 31857,
    18849 => 31856,
    18850 => 31855,
    18851 => 31855,
    18852 => 31854,
    18853 => 31853,
    18854 => 31853,
    18855 => 31852,
    18856 => 31851,
    18857 => 31850,
    18858 => 31850,
    18859 => 31849,
    18860 => 31848,
    18861 => 31847,
    18862 => 31847,
    18863 => 31846,
    18864 => 31845,
    18865 => 31844,
    18866 => 31844,
    18867 => 31843,
    18868 => 31842,
    18869 => 31841,
    18870 => 31841,
    18871 => 31840,
    18872 => 31839,
    18873 => 31838,
    18874 => 31838,
    18875 => 31837,
    18876 => 31836,
    18877 => 31836,
    18878 => 31835,
    18879 => 31834,
    18880 => 31833,
    18881 => 31833,
    18882 => 31832,
    18883 => 31831,
    18884 => 31830,
    18885 => 31830,
    18886 => 31829,
    18887 => 31828,
    18888 => 31827,
    18889 => 31827,
    18890 => 31826,
    18891 => 31825,
    18892 => 31824,
    18893 => 31824,
    18894 => 31823,
    18895 => 31822,
    18896 => 31821,
    18897 => 31821,
    18898 => 31820,
    18899 => 31819,
    18900 => 31818,
    18901 => 31818,
    18902 => 31817,
    18903 => 31816,
    18904 => 31815,
    18905 => 31815,
    18906 => 31814,
    18907 => 31813,
    18908 => 31812,
    18909 => 31812,
    18910 => 31811,
    18911 => 31810,
    18912 => 31809,
    18913 => 31809,
    18914 => 31808,
    18915 => 31807,
    18916 => 31806,
    18917 => 31806,
    18918 => 31805,
    18919 => 31804,
    18920 => 31803,
    18921 => 31802,
    18922 => 31802,
    18923 => 31801,
    18924 => 31800,
    18925 => 31799,
    18926 => 31799,
    18927 => 31798,
    18928 => 31797,
    18929 => 31796,
    18930 => 31796,
    18931 => 31795,
    18932 => 31794,
    18933 => 31793,
    18934 => 31793,
    18935 => 31792,
    18936 => 31791,
    18937 => 31790,
    18938 => 31790,
    18939 => 31789,
    18940 => 31788,
    18941 => 31787,
    18942 => 31787,
    18943 => 31786,
    18944 => 31785,
    18945 => 31784,
    18946 => 31783,
    18947 => 31783,
    18948 => 31782,
    18949 => 31781,
    18950 => 31780,
    18951 => 31780,
    18952 => 31779,
    18953 => 31778,
    18954 => 31777,
    18955 => 31777,
    18956 => 31776,
    18957 => 31775,
    18958 => 31774,
    18959 => 31774,
    18960 => 31773,
    18961 => 31772,
    18962 => 31771,
    18963 => 31770,
    18964 => 31770,
    18965 => 31769,
    18966 => 31768,
    18967 => 31767,
    18968 => 31767,
    18969 => 31766,
    18970 => 31765,
    18971 => 31764,
    18972 => 31764,
    18973 => 31763,
    18974 => 31762,
    18975 => 31761,
    18976 => 31760,
    18977 => 31760,
    18978 => 31759,
    18979 => 31758,
    18980 => 31757,
    18981 => 31757,
    18982 => 31756,
    18983 => 31755,
    18984 => 31754,
    18985 => 31753,
    18986 => 31753,
    18987 => 31752,
    18988 => 31751,
    18989 => 31750,
    18990 => 31750,
    18991 => 31749,
    18992 => 31748,
    18993 => 31747,
    18994 => 31746,
    18995 => 31746,
    18996 => 31745,
    18997 => 31744,
    18998 => 31743,
    18999 => 31743,
    19000 => 31742,
    19001 => 31741,
    19002 => 31740,
    19003 => 31739,
    19004 => 31739,
    19005 => 31738,
    19006 => 31737,
    19007 => 31736,
    19008 => 31736,
    19009 => 31735,
    19010 => 31734,
    19011 => 31733,
    19012 => 31732,
    19013 => 31732,
    19014 => 31731,
    19015 => 31730,
    19016 => 31729,
    19017 => 31729,
    19018 => 31728,
    19019 => 31727,
    19020 => 31726,
    19021 => 31725,
    19022 => 31725,
    19023 => 31724,
    19024 => 31723,
    19025 => 31722,
    19026 => 31721,
    19027 => 31721,
    19028 => 31720,
    19029 => 31719,
    19030 => 31718,
    19031 => 31718,
    19032 => 31717,
    19033 => 31716,
    19034 => 31715,
    19035 => 31714,
    19036 => 31714,
    19037 => 31713,
    19038 => 31712,
    19039 => 31711,
    19040 => 31710,
    19041 => 31710,
    19042 => 31709,
    19043 => 31708,
    19044 => 31707,
    19045 => 31706,
    19046 => 31706,
    19047 => 31705,
    19048 => 31704,
    19049 => 31703,
    19050 => 31702,
    19051 => 31702,
    19052 => 31701,
    19053 => 31700,
    19054 => 31699,
    19055 => 31698,
    19056 => 31698,
    19057 => 31697,
    19058 => 31696,
    19059 => 31695,
    19060 => 31695,
    19061 => 31694,
    19062 => 31693,
    19063 => 31692,
    19064 => 31691,
    19065 => 31691,
    19066 => 31690,
    19067 => 31689,
    19068 => 31688,
    19069 => 31687,
    19070 => 31687,
    19071 => 31686,
    19072 => 31685,
    19073 => 31684,
    19074 => 31683,
    19075 => 31683,
    19076 => 31682,
    19077 => 31681,
    19078 => 31680,
    19079 => 31679,
    19080 => 31679,
    19081 => 31678,
    19082 => 31677,
    19083 => 31676,
    19084 => 31675,
    19085 => 31674,
    19086 => 31674,
    19087 => 31673,
    19088 => 31672,
    19089 => 31671,
    19090 => 31670,
    19091 => 31670,
    19092 => 31669,
    19093 => 31668,
    19094 => 31667,
    19095 => 31666,
    19096 => 31666,
    19097 => 31665,
    19098 => 31664,
    19099 => 31663,
    19100 => 31662,
    19101 => 31662,
    19102 => 31661,
    19103 => 31660,
    19104 => 31659,
    19105 => 31658,
    19106 => 31658,
    19107 => 31657,
    19108 => 31656,
    19109 => 31655,
    19110 => 31654,
    19111 => 31653,
    19112 => 31653,
    19113 => 31652,
    19114 => 31651,
    19115 => 31650,
    19116 => 31649,
    19117 => 31649,
    19118 => 31648,
    19119 => 31647,
    19120 => 31646,
    19121 => 31645,
    19122 => 31645,
    19123 => 31644,
    19124 => 31643,
    19125 => 31642,
    19126 => 31641,
    19127 => 31640,
    19128 => 31640,
    19129 => 31639,
    19130 => 31638,
    19131 => 31637,
    19132 => 31636,
    19133 => 31636,
    19134 => 31635,
    19135 => 31634,
    19136 => 31633,
    19137 => 31632,
    19138 => 31631,
    19139 => 31631,
    19140 => 31630,
    19141 => 31629,
    19142 => 31628,
    19143 => 31627,
    19144 => 31627,
    19145 => 31626,
    19146 => 31625,
    19147 => 31624,
    19148 => 31623,
    19149 => 31622,
    19150 => 31622,
    19151 => 31621,
    19152 => 31620,
    19153 => 31619,
    19154 => 31618,
    19155 => 31617,
    19156 => 31617,
    19157 => 31616,
    19158 => 31615,
    19159 => 31614,
    19160 => 31613,
    19161 => 31613,
    19162 => 31612,
    19163 => 31611,
    19164 => 31610,
    19165 => 31609,
    19166 => 31608,
    19167 => 31608,
    19168 => 31607,
    19169 => 31606,
    19170 => 31605,
    19171 => 31604,
    19172 => 31603,
    19173 => 31603,
    19174 => 31602,
    19175 => 31601,
    19176 => 31600,
    19177 => 31599,
    19178 => 31598,
    19179 => 31598,
    19180 => 31597,
    19181 => 31596,
    19182 => 31595,
    19183 => 31594,
    19184 => 31593,
    19185 => 31593,
    19186 => 31592,
    19187 => 31591,
    19188 => 31590,
    19189 => 31589,
    19190 => 31588,
    19191 => 31588,
    19192 => 31587,
    19193 => 31586,
    19194 => 31585,
    19195 => 31584,
    19196 => 31583,
    19197 => 31583,
    19198 => 31582,
    19199 => 31581,
    19200 => 31580,
    19201 => 31579,
    19202 => 31578,
    19203 => 31578,
    19204 => 31577,
    19205 => 31576,
    19206 => 31575,
    19207 => 31574,
    19208 => 31573,
    19209 => 31572,
    19210 => 31572,
    19211 => 31571,
    19212 => 31570,
    19213 => 31569,
    19214 => 31568,
    19215 => 31567,
    19216 => 31567,
    19217 => 31566,
    19218 => 31565,
    19219 => 31564,
    19220 => 31563,
    19221 => 31562,
    19222 => 31562,
    19223 => 31561,
    19224 => 31560,
    19225 => 31559,
    19226 => 31558,
    19227 => 31557,
    19228 => 31556,
    19229 => 31556,
    19230 => 31555,
    19231 => 31554,
    19232 => 31553,
    19233 => 31552,
    19234 => 31551,
    19235 => 31551,
    19236 => 31550,
    19237 => 31549,
    19238 => 31548,
    19239 => 31547,
    19240 => 31546,
    19241 => 31545,
    19242 => 31545,
    19243 => 31544,
    19244 => 31543,
    19245 => 31542,
    19246 => 31541,
    19247 => 31540,
    19248 => 31539,
    19249 => 31539,
    19250 => 31538,
    19251 => 31537,
    19252 => 31536,
    19253 => 31535,
    19254 => 31534,
    19255 => 31534,
    19256 => 31533,
    19257 => 31532,
    19258 => 31531,
    19259 => 31530,
    19260 => 31529,
    19261 => 31528,
    19262 => 31528,
    19263 => 31527,
    19264 => 31526,
    19265 => 31525,
    19266 => 31524,
    19267 => 31523,
    19268 => 31522,
    19269 => 31522,
    19270 => 31521,
    19271 => 31520,
    19272 => 31519,
    19273 => 31518,
    19274 => 31517,
    19275 => 31516,
    19276 => 31516,
    19277 => 31515,
    19278 => 31514,
    19279 => 31513,
    19280 => 31512,
    19281 => 31511,
    19282 => 31510,
    19283 => 31510,
    19284 => 31509,
    19285 => 31508,
    19286 => 31507,
    19287 => 31506,
    19288 => 31505,
    19289 => 31504,
    19290 => 31503,
    19291 => 31503,
    19292 => 31502,
    19293 => 31501,
    19294 => 31500,
    19295 => 31499,
    19296 => 31498,
    19297 => 31497,
    19298 => 31497,
    19299 => 31496,
    19300 => 31495,
    19301 => 31494,
    19302 => 31493,
    19303 => 31492,
    19304 => 31491,
    19305 => 31490,
    19306 => 31490,
    19307 => 31489,
    19308 => 31488,
    19309 => 31487,
    19310 => 31486,
    19311 => 31485,
    19312 => 31484,
    19313 => 31484,
    19314 => 31483,
    19315 => 31482,
    19316 => 31481,
    19317 => 31480,
    19318 => 31479,
    19319 => 31478,
    19320 => 31477,
    19321 => 31477,
    19322 => 31476,
    19323 => 31475,
    19324 => 31474,
    19325 => 31473,
    19326 => 31472,
    19327 => 31471,
    19328 => 31470,
    19329 => 31470,
    19330 => 31469,
    19331 => 31468,
    19332 => 31467,
    19333 => 31466,
    19334 => 31465,
    19335 => 31464,
    19336 => 31463,
    19337 => 31463,
    19338 => 31462,
    19339 => 31461,
    19340 => 31460,
    19341 => 31459,
    19342 => 31458,
    19343 => 31457,
    19344 => 31456,
    19345 => 31456,
    19346 => 31455,
    19347 => 31454,
    19348 => 31453,
    19349 => 31452,
    19350 => 31451,
    19351 => 31450,
    19352 => 31449,
    19353 => 31448,
    19354 => 31448,
    19355 => 31447,
    19356 => 31446,
    19357 => 31445,
    19358 => 31444,
    19359 => 31443,
    19360 => 31442,
    19361 => 31441,
    19362 => 31441,
    19363 => 31440,
    19364 => 31439,
    19365 => 31438,
    19366 => 31437,
    19367 => 31436,
    19368 => 31435,
    19369 => 31434,
    19370 => 31433,
    19371 => 31433,
    19372 => 31432,
    19373 => 31431,
    19374 => 31430,
    19375 => 31429,
    19376 => 31428,
    19377 => 31427,
    19378 => 31426,
    19379 => 31425,
    19380 => 31425,
    19381 => 31424,
    19382 => 31423,
    19383 => 31422,
    19384 => 31421,
    19385 => 31420,
    19386 => 31419,
    19387 => 31418,
    19388 => 31417,
    19389 => 31417,
    19390 => 31416,
    19391 => 31415,
    19392 => 31414,
    19393 => 31413,
    19394 => 31412,
    19395 => 31411,
    19396 => 31410,
    19397 => 31409,
    19398 => 31408,
    19399 => 31408,
    19400 => 31407,
    19401 => 31406,
    19402 => 31405,
    19403 => 31404,
    19404 => 31403,
    19405 => 31402,
    19406 => 31401,
    19407 => 31400,
    19408 => 31400,
    19409 => 31399,
    19410 => 31398,
    19411 => 31397,
    19412 => 31396,
    19413 => 31395,
    19414 => 31394,
    19415 => 31393,
    19416 => 31392,
    19417 => 31391,
    19418 => 31391,
    19419 => 31390,
    19420 => 31389,
    19421 => 31388,
    19422 => 31387,
    19423 => 31386,
    19424 => 31385,
    19425 => 31384,
    19426 => 31383,
    19427 => 31382,
    19428 => 31381,
    19429 => 31381,
    19430 => 31380,
    19431 => 31379,
    19432 => 31378,
    19433 => 31377,
    19434 => 31376,
    19435 => 31375,
    19436 => 31374,
    19437 => 31373,
    19438 => 31372,
    19439 => 31372,
    19440 => 31371,
    19441 => 31370,
    19442 => 31369,
    19443 => 31368,
    19444 => 31367,
    19445 => 31366,
    19446 => 31365,
    19447 => 31364,
    19448 => 31363,
    19449 => 31362,
    19450 => 31362,
    19451 => 31361,
    19452 => 31360,
    19453 => 31359,
    19454 => 31358,
    19455 => 31357,
    19456 => 31356,
    19457 => 31355,
    19458 => 31354,
    19459 => 31353,
    19460 => 31352,
    19461 => 31352,
    19462 => 31351,
    19463 => 31350,
    19464 => 31349,
    19465 => 31348,
    19466 => 31347,
    19467 => 31346,
    19468 => 31345,
    19469 => 31344,
    19470 => 31343,
    19471 => 31342,
    19472 => 31341,
    19473 => 31341,
    19474 => 31340,
    19475 => 31339,
    19476 => 31338,
    19477 => 31337,
    19478 => 31336,
    19479 => 31335,
    19480 => 31334,
    19481 => 31333,
    19482 => 31332,
    19483 => 31331,
    19484 => 31330,
    19485 => 31329,
    19486 => 31329,
    19487 => 31328,
    19488 => 31327,
    19489 => 31326,
    19490 => 31325,
    19491 => 31324,
    19492 => 31323,
    19493 => 31322,
    19494 => 31321,
    19495 => 31320,
    19496 => 31319,
    19497 => 31318,
    19498 => 31318,
    19499 => 31317,
    19500 => 31316,
    19501 => 31315,
    19502 => 31314,
    19503 => 31313,
    19504 => 31312,
    19505 => 31311,
    19506 => 31310,
    19507 => 31309,
    19508 => 31308,
    19509 => 31307,
    19510 => 31306,
    19511 => 31305,
    19512 => 31305,
    19513 => 31304,
    19514 => 31303,
    19515 => 31302,
    19516 => 31301,
    19517 => 31300,
    19518 => 31299,
    19519 => 31298,
    19520 => 31297,
    19521 => 31296,
    19522 => 31295,
    19523 => 31294,
    19524 => 31293,
    19525 => 31292,
    19526 => 31292,
    19527 => 31291,
    19528 => 31290,
    19529 => 31289,
    19530 => 31288,
    19531 => 31287,
    19532 => 31286,
    19533 => 31285,
    19534 => 31284,
    19535 => 31283,
    19536 => 31282,
    19537 => 31281,
    19538 => 31280,
    19539 => 31279,
    19540 => 31278,
    19541 => 31278,
    19542 => 31277,
    19543 => 31276,
    19544 => 31275,
    19545 => 31274,
    19546 => 31273,
    19547 => 31272,
    19548 => 31271,
    19549 => 31270,
    19550 => 31269,
    19551 => 31268,
    19552 => 31267,
    19553 => 31266,
    19554 => 31265,
    19555 => 31264,
    19556 => 31263,
    19557 => 31262,
    19558 => 31262,
    19559 => 31261,
    19560 => 31260,
    19561 => 31259,
    19562 => 31258,
    19563 => 31257,
    19564 => 31256,
    19565 => 31255,
    19566 => 31254,
    19567 => 31253,
    19568 => 31252,
    19569 => 31251,
    19570 => 31250,
    19571 => 31249,
    19572 => 31248,
    19573 => 31247,
    19574 => 31246,
    19575 => 31246,
    19576 => 31245,
    19577 => 31244,
    19578 => 31243,
    19579 => 31242,
    19580 => 31241,
    19581 => 31240,
    19582 => 31239,
    19583 => 31238,
    19584 => 31237,
    19585 => 31236,
    19586 => 31235,
    19587 => 31234,
    19588 => 31233,
    19589 => 31232,
    19590 => 31231,
    19591 => 31230,
    19592 => 31229,
    19593 => 31228,
    19594 => 31227,
    19595 => 31227,
    19596 => 31226,
    19597 => 31225,
    19598 => 31224,
    19599 => 31223,
    19600 => 31222,
    19601 => 31221,
    19602 => 31220,
    19603 => 31219,
    19604 => 31218,
    19605 => 31217,
    19606 => 31216,
    19607 => 31215,
    19608 => 31214,
    19609 => 31213,
    19610 => 31212,
    19611 => 31211,
    19612 => 31210,
    19613 => 31209,
    19614 => 31208,
    19615 => 31207,
    19616 => 31206,
    19617 => 31206,
    19618 => 31205,
    19619 => 31204,
    19620 => 31203,
    19621 => 31202,
    19622 => 31201,
    19623 => 31200,
    19624 => 31199,
    19625 => 31198,
    19626 => 31197,
    19627 => 31196,
    19628 => 31195,
    19629 => 31194,
    19630 => 31193,
    19631 => 31192,
    19632 => 31191,
    19633 => 31190,
    19634 => 31189,
    19635 => 31188,
    19636 => 31187,
    19637 => 31186,
    19638 => 31185,
    19639 => 31184,
    19640 => 31183,
    19641 => 31182,
    19642 => 31181,
    19643 => 31181,
    19644 => 31180,
    19645 => 31179,
    19646 => 31178,
    19647 => 31177,
    19648 => 31176,
    19649 => 31175,
    19650 => 31174,
    19651 => 31173,
    19652 => 31172,
    19653 => 31171,
    19654 => 31170,
    19655 => 31169,
    19656 => 31168,
    19657 => 31167,
    19658 => 31166,
    19659 => 31165,
    19660 => 31164,
    19661 => 31163,
    19662 => 31162,
    19663 => 31161,
    19664 => 31160,
    19665 => 31159,
    19666 => 31158,
    19667 => 31157,
    19668 => 31156,
    19669 => 31155,
    19670 => 31154,
    19671 => 31153,
    19672 => 31152,
    19673 => 31151,
    19674 => 31150,
    19675 => 31149,
    19676 => 31148,
    19677 => 31148,
    19678 => 31147,
    19679 => 31146,
    19680 => 31145,
    19681 => 31144,
    19682 => 31143,
    19683 => 31142,
    19684 => 31141,
    19685 => 31140,
    19686 => 31139,
    19687 => 31138,
    19688 => 31137,
    19689 => 31136,
    19690 => 31135,
    19691 => 31134,
    19692 => 31133,
    19693 => 31132,
    19694 => 31131,
    19695 => 31130,
    19696 => 31129,
    19697 => 31128,
    19698 => 31127,
    19699 => 31126,
    19700 => 31125,
    19701 => 31124,
    19702 => 31123,
    19703 => 31122,
    19704 => 31121,
    19705 => 31120,
    19706 => 31119,
    19707 => 31118,
    19708 => 31117,
    19709 => 31116,
    19710 => 31115,
    19711 => 31114,
    19712 => 31113,
    19713 => 31112,
    19714 => 31111,
    19715 => 31110,
    19716 => 31109,
    19717 => 31108,
    19718 => 31107,
    19719 => 31106,
    19720 => 31105,
    19721 => 31104,
    19722 => 31103,
    19723 => 31102,
    19724 => 31101,
    19725 => 31100,
    19726 => 31099,
    19727 => 31098,
    19728 => 31097,
    19729 => 31096,
    19730 => 31095,
    19731 => 31094,
    19732 => 31093,
    19733 => 31092,
    19734 => 31091,
    19735 => 31090,
    19736 => 31089,
    19737 => 31088,
    19738 => 31087,
    19739 => 31086,
    19740 => 31085,
    19741 => 31084,
    19742 => 31083,
    19743 => 31083,
    19744 => 31082,
    19745 => 31081,
    19746 => 31080,
    19747 => 31079,
    19748 => 31078,
    19749 => 31077,
    19750 => 31076,
    19751 => 31075,
    19752 => 31074,
    19753 => 31073,
    19754 => 31072,
    19755 => 31071,
    19756 => 31070,
    19757 => 31069,
    19758 => 31068,
    19759 => 31067,
    19760 => 31066,
    19761 => 31065,
    19762 => 31064,
    19763 => 31063,
    19764 => 31062,
    19765 => 31061,
    19766 => 31060,
    19767 => 31059,
    19768 => 31058,
    19769 => 31057,
    19770 => 31056,
    19771 => 31055,
    19772 => 31054,
    19773 => 31053,
    19774 => 31052,
    19775 => 31051,
    19776 => 31050,
    19777 => 31049,
    19778 => 31048,
    19779 => 31047,
    19780 => 31046,
    19781 => 31045,
    19782 => 31044,
    19783 => 31043,
    19784 => 31041,
    19785 => 31040,
    19786 => 31039,
    19787 => 31038,
    19788 => 31037,
    19789 => 31036,
    19790 => 31035,
    19791 => 31034,
    19792 => 31033,
    19793 => 31032,
    19794 => 31031,
    19795 => 31030,
    19796 => 31029,
    19797 => 31028,
    19798 => 31027,
    19799 => 31026,
    19800 => 31025,
    19801 => 31024,
    19802 => 31023,
    19803 => 31022,
    19804 => 31021,
    19805 => 31020,
    19806 => 31019,
    19807 => 31018,
    19808 => 31017,
    19809 => 31016,
    19810 => 31015,
    19811 => 31014,
    19812 => 31013,
    19813 => 31012,
    19814 => 31011,
    19815 => 31010,
    19816 => 31009,
    19817 => 31008,
    19818 => 31007,
    19819 => 31006,
    19820 => 31005,
    19821 => 31004,
    19822 => 31003,
    19823 => 31002,
    19824 => 31001,
    19825 => 31000,
    19826 => 30999,
    19827 => 30998,
    19828 => 30997,
    19829 => 30996,
    19830 => 30995,
    19831 => 30994,
    19832 => 30993,
    19833 => 30992,
    19834 => 30991,
    19835 => 30990,
    19836 => 30989,
    19837 => 30988,
    19838 => 30987,
    19839 => 30986,
    19840 => 30985,
    19841 => 30984,
    19842 => 30983,
    19843 => 30982,
    19844 => 30981,
    19845 => 30980,
    19846 => 30979,
    19847 => 30978,
    19848 => 30977,
    19849 => 30976,
    19850 => 30974,
    19851 => 30973,
    19852 => 30972,
    19853 => 30971,
    19854 => 30970,
    19855 => 30969,
    19856 => 30968,
    19857 => 30967,
    19858 => 30966,
    19859 => 30965,
    19860 => 30964,
    19861 => 30963,
    19862 => 30962,
    19863 => 30961,
    19864 => 30960,
    19865 => 30959,
    19866 => 30958,
    19867 => 30957,
    19868 => 30956,
    19869 => 30955,
    19870 => 30954,
    19871 => 30953,
    19872 => 30952,
    19873 => 30951,
    19874 => 30950,
    19875 => 30949,
    19876 => 30948,
    19877 => 30947,
    19878 => 30946,
    19879 => 30945,
    19880 => 30944,
    19881 => 30943,
    19882 => 30942,
    19883 => 30941,
    19884 => 30939,
    19885 => 30938,
    19886 => 30937,
    19887 => 30936,
    19888 => 30935,
    19889 => 30934,
    19890 => 30933,
    19891 => 30932,
    19892 => 30931,
    19893 => 30930,
    19894 => 30929,
    19895 => 30928,
    19896 => 30927,
    19897 => 30926,
    19898 => 30925,
    19899 => 30924,
    19900 => 30923,
    19901 => 30922,
    19902 => 30921,
    19903 => 30920,
    19904 => 30919,
    19905 => 30918,
    19906 => 30917,
    19907 => 30916,
    19908 => 30915,
    19909 => 30914,
    19910 => 30912,
    19911 => 30911,
    19912 => 30910,
    19913 => 30909,
    19914 => 30908,
    19915 => 30907,
    19916 => 30906,
    19917 => 30905,
    19918 => 30904,
    19919 => 30903,
    19920 => 30902,
    19921 => 30901,
    19922 => 30900,
    19923 => 30899,
    19924 => 30898,
    19925 => 30897,
    19926 => 30896,
    19927 => 30895,
    19928 => 30894,
    19929 => 30893,
    19930 => 30892,
    19931 => 30891,
    19932 => 30889,
    19933 => 30888,
    19934 => 30887,
    19935 => 30886,
    19936 => 30885,
    19937 => 30884,
    19938 => 30883,
    19939 => 30882,
    19940 => 30881,
    19941 => 30880,
    19942 => 30879,
    19943 => 30878,
    19944 => 30877,
    19945 => 30876,
    19946 => 30875,
    19947 => 30874,
    19948 => 30873,
    19949 => 30872,
    19950 => 30871,
    19951 => 30870,
    19952 => 30868,
    19953 => 30867,
    19954 => 30866,
    19955 => 30865,
    19956 => 30864,
    19957 => 30863,
    19958 => 30862,
    19959 => 30861,
    19960 => 30860,
    19961 => 30859,
    19962 => 30858,
    19963 => 30857,
    19964 => 30856,
    19965 => 30855,
    19966 => 30854,
    19967 => 30853,
    19968 => 30852,
    19969 => 30851,
    19970 => 30849,
    19971 => 30848,
    19972 => 30847,
    19973 => 30846,
    19974 => 30845,
    19975 => 30844,
    19976 => 30843,
    19977 => 30842,
    19978 => 30841,
    19979 => 30840,
    19980 => 30839,
    19981 => 30838,
    19982 => 30837,
    19983 => 30836,
    19984 => 30835,
    19985 => 30834,
    19986 => 30832,
    19987 => 30831,
    19988 => 30830,
    19989 => 30829,
    19990 => 30828,
    19991 => 30827,
    19992 => 30826,
    19993 => 30825,
    19994 => 30824,
    19995 => 30823,
    19996 => 30822,
    19997 => 30821,
    19998 => 30820,
    19999 => 30819,
    20000 => 30818,
    20001 => 30816,
    20002 => 30815,
    20003 => 30814,
    20004 => 30813,
    20005 => 30812,
    20006 => 30811,
    20007 => 30810,
    20008 => 30809,
    20009 => 30808,
    20010 => 30807,
    20011 => 30806,
    20012 => 30805,
    20013 => 30804,
    20014 => 30803,
    20015 => 30802,
    20016 => 30800,
    20017 => 30799,
    20018 => 30798,
    20019 => 30797,
    20020 => 30796,
    20021 => 30795,
    20022 => 30794,
    20023 => 30793,
    20024 => 30792,
    20025 => 30791,
    20026 => 30790,
    20027 => 30789,
    20028 => 30788,
    20029 => 30786,
    20030 => 30785,
    20031 => 30784,
    20032 => 30783,
    20033 => 30782,
    20034 => 30781,
    20035 => 30780,
    20036 => 30779,
    20037 => 30778,
    20038 => 30777,
    20039 => 30776,
    20040 => 30775,
    20041 => 30774,
    20042 => 30772,
    20043 => 30771,
    20044 => 30770,
    20045 => 30769,
    20046 => 30768,
    20047 => 30767,
    20048 => 30766,
    20049 => 30765,
    20050 => 30764,
    20051 => 30763,
    20052 => 30762,
    20053 => 30761,
    20054 => 30760,
    20055 => 30758,
    20056 => 30757,
    20057 => 30756,
    20058 => 30755,
    20059 => 30754,
    20060 => 30753,
    20061 => 30752,
    20062 => 30751,
    20063 => 30750,
    20064 => 30749,
    20065 => 30748,
    20066 => 30746,
    20067 => 30745,
    20068 => 30744,
    20069 => 30743,
    20070 => 30742,
    20071 => 30741,
    20072 => 30740,
    20073 => 30739,
    20074 => 30738,
    20075 => 30737,
    20076 => 30736,
    20077 => 30735,
    20078 => 30733,
    20079 => 30732,
    20080 => 30731,
    20081 => 30730,
    20082 => 30729,
    20083 => 30728,
    20084 => 30727,
    20085 => 30726,
    20086 => 30725,
    20087 => 30724,
    20088 => 30723,
    20089 => 30721,
    20090 => 30720,
    20091 => 30719,
    20092 => 30718,
    20093 => 30717,
    20094 => 30716,
    20095 => 30715,
    20096 => 30714,
    20097 => 30713,
    20098 => 30712,
    20099 => 30711,
    20100 => 30709,
    20101 => 30708,
    20102 => 30707,
    20103 => 30706,
    20104 => 30705,
    20105 => 30704,
    20106 => 30703,
    20107 => 30702,
    20108 => 30701,
    20109 => 30700,
    20110 => 30698,
    20111 => 30697,
    20112 => 30696,
    20113 => 30695,
    20114 => 30694,
    20115 => 30693,
    20116 => 30692,
    20117 => 30691,
    20118 => 30690,
    20119 => 30689,
    20120 => 30687,
    20121 => 30686,
    20122 => 30685,
    20123 => 30684,
    20124 => 30683,
    20125 => 30682,
    20126 => 30681,
    20127 => 30680,
    20128 => 30679,
    20129 => 30678,
    20130 => 30676,
    20131 => 30675,
    20132 => 30674,
    20133 => 30673,
    20134 => 30672,
    20135 => 30671,
    20136 => 30670,
    20137 => 30669,
    20138 => 30668,
    20139 => 30666,
    20140 => 30665,
    20141 => 30664,
    20142 => 30663,
    20143 => 30662,
    20144 => 30661,
    20145 => 30660,
    20146 => 30659,
    20147 => 30658,
    20148 => 30656,
    20149 => 30655,
    20150 => 30654,
    20151 => 30653,
    20152 => 30652,
    20153 => 30651,
    20154 => 30650,
    20155 => 30649,
    20156 => 30648,
    20157 => 30646,
    20158 => 30645,
    20159 => 30644,
    20160 => 30643,
    20161 => 30642,
    20162 => 30641,
    20163 => 30640,
    20164 => 30639,
    20165 => 30638,
    20166 => 30636,
    20167 => 30635,
    20168 => 30634,
    20169 => 30633,
    20170 => 30632,
    20171 => 30631,
    20172 => 30630,
    20173 => 30629,
    20174 => 30628,
    20175 => 30626,
    20176 => 30625,
    20177 => 30624,
    20178 => 30623,
    20179 => 30622,
    20180 => 30621,
    20181 => 30620,
    20182 => 30619,
    20183 => 30617,
    20184 => 30616,
    20185 => 30615,
    20186 => 30614,
    20187 => 30613,
    20188 => 30612,
    20189 => 30611,
    20190 => 30610,
    20191 => 30609,
    20192 => 30607,
    20193 => 30606,
    20194 => 30605,
    20195 => 30604,
    20196 => 30603,
    20197 => 30602,
    20198 => 30601,
    20199 => 30600,
    20200 => 30598,
    20201 => 30597,
    20202 => 30596,
    20203 => 30595,
    20204 => 30594,
    20205 => 30593,
    20206 => 30592,
    20207 => 30591,
    20208 => 30589,
    20209 => 30588,
    20210 => 30587,
    20211 => 30586,
    20212 => 30585,
    20213 => 30584,
    20214 => 30583,
    20215 => 30582,
    20216 => 30580,
    20217 => 30579,
    20218 => 30578,
    20219 => 30577,
    20220 => 30576,
    20221 => 30575,
    20222 => 30574,
    20223 => 30573,
    20224 => 30571,
    20225 => 30570,
    20226 => 30569,
    20227 => 30568,
    20228 => 30567,
    20229 => 30566,
    20230 => 30565,
    20231 => 30563,
    20232 => 30562,
    20233 => 30561,
    20234 => 30560,
    20235 => 30559,
    20236 => 30558,
    20237 => 30557,
    20238 => 30556,
    20239 => 30554,
    20240 => 30553,
    20241 => 30552,
    20242 => 30551,
    20243 => 30550,
    20244 => 30549,
    20245 => 30548,
    20246 => 30546,
    20247 => 30545,
    20248 => 30544,
    20249 => 30543,
    20250 => 30542,
    20251 => 30541,
    20252 => 30540,
    20253 => 30538,
    20254 => 30537,
    20255 => 30536,
    20256 => 30535,
    20257 => 30534,
    20258 => 30533,
    20259 => 30532,
    20260 => 30530,
    20261 => 30529,
    20262 => 30528,
    20263 => 30527,
    20264 => 30526,
    20265 => 30525,
    20266 => 30524,
    20267 => 30522,
    20268 => 30521,
    20269 => 30520,
    20270 => 30519,
    20271 => 30518,
    20272 => 30517,
    20273 => 30516,
    20274 => 30514,
    20275 => 30513,
    20276 => 30512,
    20277 => 30511,
    20278 => 30510,
    20279 => 30509,
    20280 => 30508,
    20281 => 30506,
    20282 => 30505,
    20283 => 30504,
    20284 => 30503,
    20285 => 30502,
    20286 => 30501,
    20287 => 30500,
    20288 => 30498,
    20289 => 30497,
    20290 => 30496,
    20291 => 30495,
    20292 => 30494,
    20293 => 30493,
    20294 => 30492,
    20295 => 30490,
    20296 => 30489,
    20297 => 30488,
    20298 => 30487,
    20299 => 30486,
    20300 => 30485,
    20301 => 30483,
    20302 => 30482,
    20303 => 30481,
    20304 => 30480,
    20305 => 30479,
    20306 => 30478,
    20307 => 30477,
    20308 => 30475,
    20309 => 30474,
    20310 => 30473,
    20311 => 30472,
    20312 => 30471,
    20313 => 30470,
    20314 => 30468,
    20315 => 30467,
    20316 => 30466,
    20317 => 30465,
    20318 => 30464,
    20319 => 30463,
    20320 => 30462,
    20321 => 30460,
    20322 => 30459,
    20323 => 30458,
    20324 => 30457,
    20325 => 30456,
    20326 => 30455,
    20327 => 30453,
    20328 => 30452,
    20329 => 30451,
    20330 => 30450,
    20331 => 30449,
    20332 => 30448,
    20333 => 30446,
    20334 => 30445,
    20335 => 30444,
    20336 => 30443,
    20337 => 30442,
    20338 => 30441,
    20339 => 30439,
    20340 => 30438,
    20341 => 30437,
    20342 => 30436,
    20343 => 30435,
    20344 => 30434,
    20345 => 30433,
    20346 => 30431,
    20347 => 30430,
    20348 => 30429,
    20349 => 30428,
    20350 => 30427,
    20351 => 30426,
    20352 => 30424,
    20353 => 30423,
    20354 => 30422,
    20355 => 30421,
    20356 => 30420,
    20357 => 30419,
    20358 => 30417,
    20359 => 30416,
    20360 => 30415,
    20361 => 30414,
    20362 => 30413,
    20363 => 30412,
    20364 => 30410,
    20365 => 30409,
    20366 => 30408,
    20367 => 30407,
    20368 => 30406,
    20369 => 30404,
    20370 => 30403,
    20371 => 30402,
    20372 => 30401,
    20373 => 30400,
    20374 => 30399,
    20375 => 30397,
    20376 => 30396,
    20377 => 30395,
    20378 => 30394,
    20379 => 30393,
    20380 => 30392,
    20381 => 30390,
    20382 => 30389,
    20383 => 30388,
    20384 => 30387,
    20385 => 30386,
    20386 => 30385,
    20387 => 30383,
    20388 => 30382,
    20389 => 30381,
    20390 => 30380,
    20391 => 30379,
    20392 => 30377,
    20393 => 30376,
    20394 => 30375,
    20395 => 30374,
    20396 => 30373,
    20397 => 30372,
    20398 => 30370,
    20399 => 30369,
    20400 => 30368,
    20401 => 30367,
    20402 => 30366,
    20403 => 30365,
    20404 => 30363,
    20405 => 30362,
    20406 => 30361,
    20407 => 30360,
    20408 => 30359,
    20409 => 30357,
    20410 => 30356,
    20411 => 30355,
    20412 => 30354,
    20413 => 30353,
    20414 => 30351,
    20415 => 30350,
    20416 => 30349,
    20417 => 30348,
    20418 => 30347,
    20419 => 30346,
    20420 => 30344,
    20421 => 30343,
    20422 => 30342,
    20423 => 30341,
    20424 => 30340,
    20425 => 30338,
    20426 => 30337,
    20427 => 30336,
    20428 => 30335,
    20429 => 30334,
    20430 => 30333,
    20431 => 30331,
    20432 => 30330,
    20433 => 30329,
    20434 => 30328,
    20435 => 30327,
    20436 => 30325,
    20437 => 30324,
    20438 => 30323,
    20439 => 30322,
    20440 => 30321,
    20441 => 30319,
    20442 => 30318,
    20443 => 30317,
    20444 => 30316,
    20445 => 30315,
    20446 => 30313,
    20447 => 30312,
    20448 => 30311,
    20449 => 30310,
    20450 => 30309,
    20451 => 30308,
    20452 => 30306,
    20453 => 30305,
    20454 => 30304,
    20455 => 30303,
    20456 => 30302,
    20457 => 30300,
    20458 => 30299,
    20459 => 30298,
    20460 => 30297,
    20461 => 30296,
    20462 => 30294,
    20463 => 30293,
    20464 => 30292,
    20465 => 30291,
    20466 => 30290,
    20467 => 30288,
    20468 => 30287,
    20469 => 30286,
    20470 => 30285,
    20471 => 30284,
    20472 => 30282,
    20473 => 30281,
    20474 => 30280,
    20475 => 30279,
    20476 => 30278,
    20477 => 30276,
    20478 => 30275,
    20479 => 30274,
    20480 => 30273,
    20481 => 30272,
    20482 => 30270,
    20483 => 30269,
    20484 => 30268,
    20485 => 30267,
    20486 => 30266,
    20487 => 30264,
    20488 => 30263,
    20489 => 30262,
    20490 => 30261,
    20491 => 30260,
    20492 => 30258,
    20493 => 30257,
    20494 => 30256,
    20495 => 30255,
    20496 => 30253,
    20497 => 30252,
    20498 => 30251,
    20499 => 30250,
    20500 => 30249,
    20501 => 30247,
    20502 => 30246,
    20503 => 30245,
    20504 => 30244,
    20505 => 30243,
    20506 => 30241,
    20507 => 30240,
    20508 => 30239,
    20509 => 30238,
    20510 => 30237,
    20511 => 30235,
    20512 => 30234,
    20513 => 30233,
    20514 => 30232,
    20515 => 30231,
    20516 => 30229,
    20517 => 30228,
    20518 => 30227,
    20519 => 30226,
    20520 => 30224,
    20521 => 30223,
    20522 => 30222,
    20523 => 30221,
    20524 => 30220,
    20525 => 30218,
    20526 => 30217,
    20527 => 30216,
    20528 => 30215,
    20529 => 30214,
    20530 => 30212,
    20531 => 30211,
    20532 => 30210,
    20533 => 30209,
    20534 => 30207,
    20535 => 30206,
    20536 => 30205,
    20537 => 30204,
    20538 => 30203,
    20539 => 30201,
    20540 => 30200,
    20541 => 30199,
    20542 => 30198,
    20543 => 30196,
    20544 => 30195,
    20545 => 30194,
    20546 => 30193,
    20547 => 30192,
    20548 => 30190,
    20549 => 30189,
    20550 => 30188,
    20551 => 30187,
    20552 => 30185,
    20553 => 30184,
    20554 => 30183,
    20555 => 30182,
    20556 => 30181,
    20557 => 30179,
    20558 => 30178,
    20559 => 30177,
    20560 => 30176,
    20561 => 30174,
    20562 => 30173,
    20563 => 30172,
    20564 => 30171,
    20565 => 30170,
    20566 => 30168,
    20567 => 30167,
    20568 => 30166,
    20569 => 30165,
    20570 => 30163,
    20571 => 30162,
    20572 => 30161,
    20573 => 30160,
    20574 => 30159,
    20575 => 30157,
    20576 => 30156,
    20577 => 30155,
    20578 => 30154,
    20579 => 30152,
    20580 => 30151,
    20581 => 30150,
    20582 => 30149,
    20583 => 30147,
    20584 => 30146,
    20585 => 30145,
    20586 => 30144,
    20587 => 30143,
    20588 => 30141,
    20589 => 30140,
    20590 => 30139,
    20591 => 30138,
    20592 => 30136,
    20593 => 30135,
    20594 => 30134,
    20595 => 30133,
    20596 => 30131,
    20597 => 30130,
    20598 => 30129,
    20599 => 30128,
    20600 => 30126,
    20601 => 30125,
    20602 => 30124,
    20603 => 30123,
    20604 => 30122,
    20605 => 30120,
    20606 => 30119,
    20607 => 30118,
    20608 => 30117,
    20609 => 30115,
    20610 => 30114,
    20611 => 30113,
    20612 => 30112,
    20613 => 30110,
    20614 => 30109,
    20615 => 30108,
    20616 => 30107,
    20617 => 30105,
    20618 => 30104,
    20619 => 30103,
    20620 => 30102,
    20621 => 30100,
    20622 => 30099,
    20623 => 30098,
    20624 => 30097,
    20625 => 30096,
    20626 => 30094,
    20627 => 30093,
    20628 => 30092,
    20629 => 30091,
    20630 => 30089,
    20631 => 30088,
    20632 => 30087,
    20633 => 30086,
    20634 => 30084,
    20635 => 30083,
    20636 => 30082,
    20637 => 30081,
    20638 => 30079,
    20639 => 30078,
    20640 => 30077,
    20641 => 30076,
    20642 => 30074,
    20643 => 30073,
    20644 => 30072,
    20645 => 30071,
    20646 => 30069,
    20647 => 30068,
    20648 => 30067,
    20649 => 30066,
    20650 => 30064,
    20651 => 30063,
    20652 => 30062,
    20653 => 30061,
    20654 => 30059,
    20655 => 30058,
    20656 => 30057,
    20657 => 30056,
    20658 => 30054,
    20659 => 30053,
    20660 => 30052,
    20661 => 30051,
    20662 => 30049,
    20663 => 30048,
    20664 => 30047,
    20665 => 30046,
    20666 => 30044,
    20667 => 30043,
    20668 => 30042,
    20669 => 30041,
    20670 => 30039,
    20671 => 30038,
    20672 => 30037,
    20673 => 30036,
    20674 => 30034,
    20675 => 30033,
    20676 => 30032,
    20677 => 30031,
    20678 => 30029,
    20679 => 30028,
    20680 => 30027,
    20681 => 30026,
    20682 => 30024,
    20683 => 30023,
    20684 => 30022,
    20685 => 30020,
    20686 => 30019,
    20687 => 30018,
    20688 => 30017,
    20689 => 30015,
    20690 => 30014,
    20691 => 30013,
    20692 => 30012,
    20693 => 30010,
    20694 => 30009,
    20695 => 30008,
    20696 => 30007,
    20697 => 30005,
    20698 => 30004,
    20699 => 30003,
    20700 => 30002,
    20701 => 30000,
    20702 => 29999,
    20703 => 29998,
    20704 => 29997,
    20705 => 29995,
    20706 => 29994,
    20707 => 29993,
    20708 => 29991,
    20709 => 29990,
    20710 => 29989,
    20711 => 29988,
    20712 => 29986,
    20713 => 29985,
    20714 => 29984,
    20715 => 29983,
    20716 => 29981,
    20717 => 29980,
    20718 => 29979,
    20719 => 29978,
    20720 => 29976,
    20721 => 29975,
    20722 => 29974,
    20723 => 29972,
    20724 => 29971,
    20725 => 29970,
    20726 => 29969,
    20727 => 29967,
    20728 => 29966,
    20729 => 29965,
    20730 => 29964,
    20731 => 29962,
    20732 => 29961,
    20733 => 29960,
    20734 => 29958,
    20735 => 29957,
    20736 => 29956,
    20737 => 29955,
    20738 => 29953,
    20739 => 29952,
    20740 => 29951,
    20741 => 29950,
    20742 => 29948,
    20743 => 29947,
    20744 => 29946,
    20745 => 29944,
    20746 => 29943,
    20747 => 29942,
    20748 => 29941,
    20749 => 29939,
    20750 => 29938,
    20751 => 29937,
    20752 => 29936,
    20753 => 29934,
    20754 => 29933,
    20755 => 29932,
    20756 => 29930,
    20757 => 29929,
    20758 => 29928,
    20759 => 29927,
    20760 => 29925,
    20761 => 29924,
    20762 => 29923,
    20763 => 29921,
    20764 => 29920,
    20765 => 29919,
    20766 => 29918,
    20767 => 29916,
    20768 => 29915,
    20769 => 29914,
    20770 => 29912,
    20771 => 29911,
    20772 => 29910,
    20773 => 29909,
    20774 => 29907,
    20775 => 29906,
    20776 => 29905,
    20777 => 29903,
    20778 => 29902,
    20779 => 29901,
    20780 => 29900,
    20781 => 29898,
    20782 => 29897,
    20783 => 29896,
    20784 => 29894,
    20785 => 29893,
    20786 => 29892,
    20787 => 29891,
    20788 => 29889,
    20789 => 29888,
    20790 => 29887,
    20791 => 29885,
    20792 => 29884,
    20793 => 29883,
    20794 => 29882,
    20795 => 29880,
    20796 => 29879,
    20797 => 29878,
    20798 => 29876,
    20799 => 29875,
    20800 => 29874,
    20801 => 29873,
    20802 => 29871,
    20803 => 29870,
    20804 => 29869,
    20805 => 29867,
    20806 => 29866,
    20807 => 29865,
    20808 => 29864,
    20809 => 29862,
    20810 => 29861,
    20811 => 29860,
    20812 => 29858,
    20813 => 29857,
    20814 => 29856,
    20815 => 29854,
    20816 => 29853,
    20817 => 29852,
    20818 => 29851,
    20819 => 29849,
    20820 => 29848,
    20821 => 29847,
    20822 => 29845,
    20823 => 29844,
    20824 => 29843,
    20825 => 29842,
    20826 => 29840,
    20827 => 29839,
    20828 => 29838,
    20829 => 29836,
    20830 => 29835,
    20831 => 29834,
    20832 => 29832,
    20833 => 29831,
    20834 => 29830,
    20835 => 29829,
    20836 => 29827,
    20837 => 29826,
    20838 => 29825,
    20839 => 29823,
    20840 => 29822,
    20841 => 29821,
    20842 => 29819,
    20843 => 29818,
    20844 => 29817,
    20845 => 29816,
    20846 => 29814,
    20847 => 29813,
    20848 => 29812,
    20849 => 29810,
    20850 => 29809,
    20851 => 29808,
    20852 => 29806,
    20853 => 29805,
    20854 => 29804,
    20855 => 29802,
    20856 => 29801,
    20857 => 29800,
    20858 => 29799,
    20859 => 29797,
    20860 => 29796,
    20861 => 29795,
    20862 => 29793,
    20863 => 29792,
    20864 => 29791,
    20865 => 29789,
    20866 => 29788,
    20867 => 29787,
    20868 => 29785,
    20869 => 29784,
    20870 => 29783,
    20871 => 29782,
    20872 => 29780,
    20873 => 29779,
    20874 => 29778,
    20875 => 29776,
    20876 => 29775,
    20877 => 29774,
    20878 => 29772,
    20879 => 29771,
    20880 => 29770,
    20881 => 29768,
    20882 => 29767,
    20883 => 29766,
    20884 => 29764,
    20885 => 29763,
    20886 => 29762,
    20887 => 29761,
    20888 => 29759,
    20889 => 29758,
    20890 => 29757,
    20891 => 29755,
    20892 => 29754,
    20893 => 29753,
    20894 => 29751,
    20895 => 29750,
    20896 => 29749,
    20897 => 29747,
    20898 => 29746,
    20899 => 29745,
    20900 => 29743,
    20901 => 29742,
    20902 => 29741,
    20903 => 29739,
    20904 => 29738,
    20905 => 29737,
    20906 => 29736,
    20907 => 29734,
    20908 => 29733,
    20909 => 29732,
    20910 => 29730,
    20911 => 29729,
    20912 => 29728,
    20913 => 29726,
    20914 => 29725,
    20915 => 29724,
    20916 => 29722,
    20917 => 29721,
    20918 => 29720,
    20919 => 29718,
    20920 => 29717,
    20921 => 29716,
    20922 => 29714,
    20923 => 29713,
    20924 => 29712,
    20925 => 29710,
    20926 => 29709,
    20927 => 29708,
    20928 => 29706,
    20929 => 29705,
    20930 => 29704,
    20931 => 29702,
    20932 => 29701,
    20933 => 29700,
    20934 => 29698,
    20935 => 29697,
    20936 => 29696,
    20937 => 29694,
    20938 => 29693,
    20939 => 29692,
    20940 => 29690,
    20941 => 29689,
    20942 => 29688,
    20943 => 29687,
    20944 => 29685,
    20945 => 29684,
    20946 => 29683,
    20947 => 29681,
    20948 => 29680,
    20949 => 29679,
    20950 => 29677,
    20951 => 29676,
    20952 => 29675,
    20953 => 29673,
    20954 => 29672,
    20955 => 29671,
    20956 => 29669,
    20957 => 29668,
    20958 => 29667,
    20959 => 29665,
    20960 => 29664,
    20961 => 29663,
    20962 => 29661,
    20963 => 29660,
    20964 => 29659,
    20965 => 29657,
    20966 => 29656,
    20967 => 29655,
    20968 => 29653,
    20969 => 29652,
    20970 => 29651,
    20971 => 29649,
    20972 => 29648,
    20973 => 29646,
    20974 => 29645,
    20975 => 29644,
    20976 => 29642,
    20977 => 29641,
    20978 => 29640,
    20979 => 29638,
    20980 => 29637,
    20981 => 29636,
    20982 => 29634,
    20983 => 29633,
    20984 => 29632,
    20985 => 29630,
    20986 => 29629,
    20987 => 29628,
    20988 => 29626,
    20989 => 29625,
    20990 => 29624,
    20991 => 29622,
    20992 => 29621,
    20993 => 29620,
    20994 => 29618,
    20995 => 29617,
    20996 => 29616,
    20997 => 29614,
    20998 => 29613,
    20999 => 29612,
    21000 => 29610,
    21001 => 29609,
    21002 => 29608,
    21003 => 29606,
    21004 => 29605,
    21005 => 29604,
    21006 => 29602,
    21007 => 29601,
    21008 => 29599,
    21009 => 29598,
    21010 => 29597,
    21011 => 29595,
    21012 => 29594,
    21013 => 29593,
    21014 => 29591,
    21015 => 29590,
    21016 => 29589,
    21017 => 29587,
    21018 => 29586,
    21019 => 29585,
    21020 => 29583,
    21021 => 29582,
    21022 => 29581,
    21023 => 29579,
    21024 => 29578,
    21025 => 29577,
    21026 => 29575,
    21027 => 29574,
    21028 => 29572,
    21029 => 29571,
    21030 => 29570,
    21031 => 29568,
    21032 => 29567,
    21033 => 29566,
    21034 => 29564,
    21035 => 29563,
    21036 => 29562,
    21037 => 29560,
    21038 => 29559,
    21039 => 29558,
    21040 => 29556,
    21041 => 29555,
    21042 => 29554,
    21043 => 29552,
    21044 => 29551,
    21045 => 29549,
    21046 => 29548,
    21047 => 29547,
    21048 => 29545,
    21049 => 29544,
    21050 => 29543,
    21051 => 29541,
    21052 => 29540,
    21053 => 29539,
    21054 => 29537,
    21055 => 29536,
    21056 => 29534,
    21057 => 29533,
    21058 => 29532,
    21059 => 29530,
    21060 => 29529,
    21061 => 29528,
    21062 => 29526,
    21063 => 29525,
    21064 => 29524,
    21065 => 29522,
    21066 => 29521,
    21067 => 29520,
    21068 => 29518,
    21069 => 29517,
    21070 => 29515,
    21071 => 29514,
    21072 => 29513,
    21073 => 29511,
    21074 => 29510,
    21075 => 29509,
    21076 => 29507,
    21077 => 29506,
    21078 => 29504,
    21079 => 29503,
    21080 => 29502,
    21081 => 29500,
    21082 => 29499,
    21083 => 29498,
    21084 => 29496,
    21085 => 29495,
    21086 => 29494,
    21087 => 29492,
    21088 => 29491,
    21089 => 29489,
    21090 => 29488,
    21091 => 29487,
    21092 => 29485,
    21093 => 29484,
    21094 => 29483,
    21095 => 29481,
    21096 => 29480,
    21097 => 29478,
    21098 => 29477,
    21099 => 29476,
    21100 => 29474,
    21101 => 29473,
    21102 => 29472,
    21103 => 29470,
    21104 => 29469,
    21105 => 29468,
    21106 => 29466,
    21107 => 29465,
    21108 => 29463,
    21109 => 29462,
    21110 => 29461,
    21111 => 29459,
    21112 => 29458,
    21113 => 29457,
    21114 => 29455,
    21115 => 29454,
    21116 => 29452,
    21117 => 29451,
    21118 => 29450,
    21119 => 29448,
    21120 => 29447,
    21121 => 29445,
    21122 => 29444,
    21123 => 29443,
    21124 => 29441,
    21125 => 29440,
    21126 => 29439,
    21127 => 29437,
    21128 => 29436,
    21129 => 29434,
    21130 => 29433,
    21131 => 29432,
    21132 => 29430,
    21133 => 29429,
    21134 => 29428,
    21135 => 29426,
    21136 => 29425,
    21137 => 29423,
    21138 => 29422,
    21139 => 29421,
    21140 => 29419,
    21141 => 29418,
    21142 => 29416,
    21143 => 29415,
    21144 => 29414,
    21145 => 29412,
    21146 => 29411,
    21147 => 29410,
    21148 => 29408,
    21149 => 29407,
    21150 => 29405,
    21151 => 29404,
    21152 => 29403,
    21153 => 29401,
    21154 => 29400,
    21155 => 29398,
    21156 => 29397,
    21157 => 29396,
    21158 => 29394,
    21159 => 29393,
    21160 => 29392,
    21161 => 29390,
    21162 => 29389,
    21163 => 29387,
    21164 => 29386,
    21165 => 29385,
    21166 => 29383,
    21167 => 29382,
    21168 => 29380,
    21169 => 29379,
    21170 => 29378,
    21171 => 29376,
    21172 => 29375,
    21173 => 29373,
    21174 => 29372,
    21175 => 29371,
    21176 => 29369,
    21177 => 29368,
    21178 => 29366,
    21179 => 29365,
    21180 => 29364,
    21181 => 29362,
    21182 => 29361,
    21183 => 29360,
    21184 => 29358,
    21185 => 29357,
    21186 => 29355,
    21187 => 29354,
    21188 => 29353,
    21189 => 29351,
    21190 => 29350,
    21191 => 29348,
    21192 => 29347,
    21193 => 29346,
    21194 => 29344,
    21195 => 29343,
    21196 => 29341,
    21197 => 29340,
    21198 => 29339,
    21199 => 29337,
    21200 => 29336,
    21201 => 29334,
    21202 => 29333,
    21203 => 29332,
    21204 => 29330,
    21205 => 29329,
    21206 => 29327,
    21207 => 29326,
    21208 => 29325,
    21209 => 29323,
    21210 => 29322,
    21211 => 29320,
    21212 => 29319,
    21213 => 29318,
    21214 => 29316,
    21215 => 29315,
    21216 => 29313,
    21217 => 29312,
    21218 => 29311,
    21219 => 29309,
    21220 => 29308,
    21221 => 29306,
    21222 => 29305,
    21223 => 29304,
    21224 => 29302,
    21225 => 29301,
    21226 => 29299,
    21227 => 29298,
    21228 => 29296,
    21229 => 29295,
    21230 => 29294,
    21231 => 29292,
    21232 => 29291,
    21233 => 29289,
    21234 => 29288,
    21235 => 29287,
    21236 => 29285,
    21237 => 29284,
    21238 => 29282,
    21239 => 29281,
    21240 => 29280,
    21241 => 29278,
    21242 => 29277,
    21243 => 29275,
    21244 => 29274,
    21245 => 29273,
    21246 => 29271,
    21247 => 29270,
    21248 => 29268,
    21249 => 29267,
    21250 => 29265,
    21251 => 29264,
    21252 => 29263,
    21253 => 29261,
    21254 => 29260,
    21255 => 29258,
    21256 => 29257,
    21257 => 29256,
    21258 => 29254,
    21259 => 29253,
    21260 => 29251,
    21261 => 29250,
    21262 => 29248,
    21263 => 29247,
    21264 => 29246,
    21265 => 29244,
    21266 => 29243,
    21267 => 29241,
    21268 => 29240,
    21269 => 29239,
    21270 => 29237,
    21271 => 29236,
    21272 => 29234,
    21273 => 29233,
    21274 => 29231,
    21275 => 29230,
    21276 => 29229,
    21277 => 29227,
    21278 => 29226,
    21279 => 29224,
    21280 => 29223,
    21281 => 29222,
    21282 => 29220,
    21283 => 29219,
    21284 => 29217,
    21285 => 29216,
    21286 => 29214,
    21287 => 29213,
    21288 => 29212,
    21289 => 29210,
    21290 => 29209,
    21291 => 29207,
    21292 => 29206,
    21293 => 29204,
    21294 => 29203,
    21295 => 29202,
    21296 => 29200,
    21297 => 29199,
    21298 => 29197,
    21299 => 29196,
    21300 => 29194,
    21301 => 29193,
    21302 => 29192,
    21303 => 29190,
    21304 => 29189,
    21305 => 29187,
    21306 => 29186,
    21307 => 29184,
    21308 => 29183,
    21309 => 29182,
    21310 => 29180,
    21311 => 29179,
    21312 => 29177,
    21313 => 29176,
    21314 => 29174,
    21315 => 29173,
    21316 => 29172,
    21317 => 29170,
    21318 => 29169,
    21319 => 29167,
    21320 => 29166,
    21321 => 29164,
    21322 => 29163,
    21323 => 29162,
    21324 => 29160,
    21325 => 29159,
    21326 => 29157,
    21327 => 29156,
    21328 => 29154,
    21329 => 29153,
    21330 => 29152,
    21331 => 29150,
    21332 => 29149,
    21333 => 29147,
    21334 => 29146,
    21335 => 29144,
    21336 => 29143,
    21337 => 29142,
    21338 => 29140,
    21339 => 29139,
    21340 => 29137,
    21341 => 29136,
    21342 => 29134,
    21343 => 29133,
    21344 => 29131,
    21345 => 29130,
    21346 => 29129,
    21347 => 29127,
    21348 => 29126,
    21349 => 29124,
    21350 => 29123,
    21351 => 29121,
    21352 => 29120,
    21353 => 29118,
    21354 => 29117,
    21355 => 29116,
    21356 => 29114,
    21357 => 29113,
    21358 => 29111,
    21359 => 29110,
    21360 => 29108,
    21361 => 29107,
    21362 => 29106,
    21363 => 29104,
    21364 => 29103,
    21365 => 29101,
    21366 => 29100,
    21367 => 29098,
    21368 => 29097,
    21369 => 29095,
    21370 => 29094,
    21371 => 29093,
    21372 => 29091,
    21373 => 29090,
    21374 => 29088,
    21375 => 29087,
    21376 => 29085,
    21377 => 29084,
    21378 => 29082,
    21379 => 29081,
    21380 => 29079,
    21381 => 29078,
    21382 => 29077,
    21383 => 29075,
    21384 => 29074,
    21385 => 29072,
    21386 => 29071,
    21387 => 29069,
    21388 => 29068,
    21389 => 29066,
    21390 => 29065,
    21391 => 29064,
    21392 => 29062,
    21393 => 29061,
    21394 => 29059,
    21395 => 29058,
    21396 => 29056,
    21397 => 29055,
    21398 => 29053,
    21399 => 29052,
    21400 => 29050,
    21401 => 29049,
    21402 => 29048,
    21403 => 29046,
    21404 => 29045,
    21405 => 29043,
    21406 => 29042,
    21407 => 29040,
    21408 => 29039,
    21409 => 29037,
    21410 => 29036,
    21411 => 29034,
    21412 => 29033,
    21413 => 29032,
    21414 => 29030,
    21415 => 29029,
    21416 => 29027,
    21417 => 29026,
    21418 => 29024,
    21419 => 29023,
    21420 => 29021,
    21421 => 29020,
    21422 => 29018,
    21423 => 29017,
    21424 => 29016,
    21425 => 29014,
    21426 => 29013,
    21427 => 29011,
    21428 => 29010,
    21429 => 29008,
    21430 => 29007,
    21431 => 29005,
    21432 => 29004,
    21433 => 29002,
    21434 => 29001,
    21435 => 28999,
    21436 => 28998,
    21437 => 28997,
    21438 => 28995,
    21439 => 28994,
    21440 => 28992,
    21441 => 28991,
    21442 => 28989,
    21443 => 28988,
    21444 => 28986,
    21445 => 28985,
    21446 => 28983,
    21447 => 28982,
    21448 => 28980,
    21449 => 28979,
    21450 => 28977,
    21451 => 28976,
    21452 => 28975,
    21453 => 28973,
    21454 => 28972,
    21455 => 28970,
    21456 => 28969,
    21457 => 28967,
    21458 => 28966,
    21459 => 28964,
    21460 => 28963,
    21461 => 28961,
    21462 => 28960,
    21463 => 28958,
    21464 => 28957,
    21465 => 28955,
    21466 => 28954,
    21467 => 28953,
    21468 => 28951,
    21469 => 28950,
    21470 => 28948,
    21471 => 28947,
    21472 => 28945,
    21473 => 28944,
    21474 => 28942,
    21475 => 28941,
    21476 => 28939,
    21477 => 28938,
    21478 => 28936,
    21479 => 28935,
    21480 => 28933,
    21481 => 28932,
    21482 => 28930,
    21483 => 28929,
    21484 => 28927,
    21485 => 28926,
    21486 => 28925,
    21487 => 28923,
    21488 => 28922,
    21489 => 28920,
    21490 => 28919,
    21491 => 28917,
    21492 => 28916,
    21493 => 28914,
    21494 => 28913,
    21495 => 28911,
    21496 => 28910,
    21497 => 28908,
    21498 => 28907,
    21499 => 28905,
    21500 => 28904,
    21501 => 28902,
    21502 => 28901,
    21503 => 28899,
    21504 => 28898,
    21505 => 28896,
    21506 => 28895,
    21507 => 28893,
    21508 => 28892,
    21509 => 28891,
    21510 => 28889,
    21511 => 28888,
    21512 => 28886,
    21513 => 28885,
    21514 => 28883,
    21515 => 28882,
    21516 => 28880,
    21517 => 28879,
    21518 => 28877,
    21519 => 28876,
    21520 => 28874,
    21521 => 28873,
    21522 => 28871,
    21523 => 28870,
    21524 => 28868,
    21525 => 28867,
    21526 => 28865,
    21527 => 28864,
    21528 => 28862,
    21529 => 28861,
    21530 => 28859,
    21531 => 28858,
    21532 => 28856,
    21533 => 28855,
    21534 => 28853,
    21535 => 28852,
    21536 => 28850,
    21537 => 28849,
    21538 => 28847,
    21539 => 28846,
    21540 => 28844,
    21541 => 28843,
    21542 => 28841,
    21543 => 28840,
    21544 => 28838,
    21545 => 28837,
    21546 => 28835,
    21547 => 28834,
    21548 => 28832,
    21549 => 28831,
    21550 => 28830,
    21551 => 28828,
    21552 => 28827,
    21553 => 28825,
    21554 => 28824,
    21555 => 28822,
    21556 => 28821,
    21557 => 28819,
    21558 => 28818,
    21559 => 28816,
    21560 => 28815,
    21561 => 28813,
    21562 => 28812,
    21563 => 28810,
    21564 => 28809,
    21565 => 28807,
    21566 => 28806,
    21567 => 28804,
    21568 => 28803,
    21569 => 28801,
    21570 => 28800,
    21571 => 28798,
    21572 => 28797,
    21573 => 28795,
    21574 => 28794,
    21575 => 28792,
    21576 => 28791,
    21577 => 28789,
    21578 => 28788,
    21579 => 28786,
    21580 => 28785,
    21581 => 28783,
    21582 => 28782,
    21583 => 28780,
    21584 => 28779,
    21585 => 28777,
    21586 => 28776,
    21587 => 28774,
    21588 => 28773,
    21589 => 28771,
    21590 => 28770,
    21591 => 28768,
    21592 => 28767,
    21593 => 28765,
    21594 => 28764,
    21595 => 28762,
    21596 => 28761,
    21597 => 28759,
    21598 => 28758,
    21599 => 28756,
    21600 => 28755,
    21601 => 28753,
    21602 => 28752,
    21603 => 28750,
    21604 => 28748,
    21605 => 28747,
    21606 => 28745,
    21607 => 28744,
    21608 => 28742,
    21609 => 28741,
    21610 => 28739,
    21611 => 28738,
    21612 => 28736,
    21613 => 28735,
    21614 => 28733,
    21615 => 28732,
    21616 => 28730,
    21617 => 28729,
    21618 => 28727,
    21619 => 28726,
    21620 => 28724,
    21621 => 28723,
    21622 => 28721,
    21623 => 28720,
    21624 => 28718,
    21625 => 28717,
    21626 => 28715,
    21627 => 28714,
    21628 => 28712,
    21629 => 28711,
    21630 => 28709,
    21631 => 28708,
    21632 => 28706,
    21633 => 28705,
    21634 => 28703,
    21635 => 28702,
    21636 => 28700,
    21637 => 28699,
    21638 => 28697,
    21639 => 28696,
    21640 => 28694,
    21641 => 28693,
    21642 => 28691,
    21643 => 28690,
    21644 => 28688,
    21645 => 28686,
    21646 => 28685,
    21647 => 28683,
    21648 => 28682,
    21649 => 28680,
    21650 => 28679,
    21651 => 28677,
    21652 => 28676,
    21653 => 28674,
    21654 => 28673,
    21655 => 28671,
    21656 => 28670,
    21657 => 28668,
    21658 => 28667,
    21659 => 28665,
    21660 => 28664,
    21661 => 28662,
    21662 => 28661,
    21663 => 28659,
    21664 => 28658,
    21665 => 28656,
    21666 => 28655,
    21667 => 28653,
    21668 => 28651,
    21669 => 28650,
    21670 => 28648,
    21671 => 28647,
    21672 => 28645,
    21673 => 28644,
    21674 => 28642,
    21675 => 28641,
    21676 => 28639,
    21677 => 28638,
    21678 => 28636,
    21679 => 28635,
    21680 => 28633,
    21681 => 28632,
    21682 => 28630,
    21683 => 28629,
    21684 => 28627,
    21685 => 28626,
    21686 => 28624,
    21687 => 28622,
    21688 => 28621,
    21689 => 28619,
    21690 => 28618,
    21691 => 28616,
    21692 => 28615,
    21693 => 28613,
    21694 => 28612,
    21695 => 28610,
    21696 => 28609,
    21697 => 28607,
    21698 => 28606,
    21699 => 28604,
    21700 => 28603,
    21701 => 28601,
    21702 => 28600,
    21703 => 28598,
    21704 => 28596,
    21705 => 28595,
    21706 => 28593,
    21707 => 28592,
    21708 => 28590,
    21709 => 28589,
    21710 => 28587,
    21711 => 28586,
    21712 => 28584,
    21713 => 28583,
    21714 => 28581,
    21715 => 28580,
    21716 => 28578,
    21717 => 28576,
    21718 => 28575,
    21719 => 28573,
    21720 => 28572,
    21721 => 28570,
    21722 => 28569,
    21723 => 28567,
    21724 => 28566,
    21725 => 28564,
    21726 => 28563,
    21727 => 28561,
    21728 => 28560,
    21729 => 28558,
    21730 => 28556,
    21731 => 28555,
    21732 => 28553,
    21733 => 28552,
    21734 => 28550,
    21735 => 28549,
    21736 => 28547,
    21737 => 28546,
    21738 => 28544,
    21739 => 28543,
    21740 => 28541,
    21741 => 28540,
    21742 => 28538,
    21743 => 28536,
    21744 => 28535,
    21745 => 28533,
    21746 => 28532,
    21747 => 28530,
    21748 => 28529,
    21749 => 28527,
    21750 => 28526,
    21751 => 28524,
    21752 => 28523,
    21753 => 28521,
    21754 => 28519,
    21755 => 28518,
    21756 => 28516,
    21757 => 28515,
    21758 => 28513,
    21759 => 28512,
    21760 => 28510,
    21761 => 28509,
    21762 => 28507,
    21763 => 28505,
    21764 => 28504,
    21765 => 28502,
    21766 => 28501,
    21767 => 28499,
    21768 => 28498,
    21769 => 28496,
    21770 => 28495,
    21771 => 28493,
    21772 => 28492,
    21773 => 28490,
    21774 => 28488,
    21775 => 28487,
    21776 => 28485,
    21777 => 28484,
    21778 => 28482,
    21779 => 28481,
    21780 => 28479,
    21781 => 28478,
    21782 => 28476,
    21783 => 28474,
    21784 => 28473,
    21785 => 28471,
    21786 => 28470,
    21787 => 28468,
    21788 => 28467,
    21789 => 28465,
    21790 => 28464,
    21791 => 28462,
    21792 => 28460,
    21793 => 28459,
    21794 => 28457,
    21795 => 28456,
    21796 => 28454,
    21797 => 28453,
    21798 => 28451,
    21799 => 28450,
    21800 => 28448,
    21801 => 28446,
    21802 => 28445,
    21803 => 28443,
    21804 => 28442,
    21805 => 28440,
    21806 => 28439,
    21807 => 28437,
    21808 => 28436,
    21809 => 28434,
    21810 => 28432,
    21811 => 28431,
    21812 => 28429,
    21813 => 28428,
    21814 => 28426,
    21815 => 28425,
    21816 => 28423,
    21817 => 28421,
    21818 => 28420,
    21819 => 28418,
    21820 => 28417,
    21821 => 28415,
    21822 => 28414,
    21823 => 28412,
    21824 => 28411,
    21825 => 28409,
    21826 => 28407,
    21827 => 28406,
    21828 => 28404,
    21829 => 28403,
    21830 => 28401,
    21831 => 28400,
    21832 => 28398,
    21833 => 28396,
    21834 => 28395,
    21835 => 28393,
    21836 => 28392,
    21837 => 28390,
    21838 => 28389,
    21839 => 28387,
    21840 => 28385,
    21841 => 28384,
    21842 => 28382,
    21843 => 28381,
    21844 => 28379,
    21845 => 28378,
    21846 => 28376,
    21847 => 28374,
    21848 => 28373,
    21849 => 28371,
    21850 => 28370,
    21851 => 28368,
    21852 => 28367,
    21853 => 28365,
    21854 => 28363,
    21855 => 28362,
    21856 => 28360,
    21857 => 28359,
    21858 => 28357,
    21859 => 28356,
    21860 => 28354,
    21861 => 28352,
    21862 => 28351,
    21863 => 28349,
    21864 => 28348,
    21865 => 28346,
    21866 => 28345,
    21867 => 28343,
    21868 => 28341,
    21869 => 28340,
    21870 => 28338,
    21871 => 28337,
    21872 => 28335,
    21873 => 28333,
    21874 => 28332,
    21875 => 28330,
    21876 => 28329,
    21877 => 28327,
    21878 => 28326,
    21879 => 28324,
    21880 => 28322,
    21881 => 28321,
    21882 => 28319,
    21883 => 28318,
    21884 => 28316,
    21885 => 28315,
    21886 => 28313,
    21887 => 28311,
    21888 => 28310,
    21889 => 28308,
    21890 => 28307,
    21891 => 28305,
    21892 => 28303,
    21893 => 28302,
    21894 => 28300,
    21895 => 28299,
    21896 => 28297,
    21897 => 28296,
    21898 => 28294,
    21899 => 28292,
    21900 => 28291,
    21901 => 28289,
    21902 => 28288,
    21903 => 28286,
    21904 => 28284,
    21905 => 28283,
    21906 => 28281,
    21907 => 28280,
    21908 => 28278,
    21909 => 28277,
    21910 => 28275,
    21911 => 28273,
    21912 => 28272,
    21913 => 28270,
    21914 => 28269,
    21915 => 28267,
    21916 => 28265,
    21917 => 28264,
    21918 => 28262,
    21919 => 28261,
    21920 => 28259,
    21921 => 28257,
    21922 => 28256,
    21923 => 28254,
    21924 => 28253,
    21925 => 28251,
    21926 => 28249,
    21927 => 28248,
    21928 => 28246,
    21929 => 28245,
    21930 => 28243,
    21931 => 28242,
    21932 => 28240,
    21933 => 28238,
    21934 => 28237,
    21935 => 28235,
    21936 => 28234,
    21937 => 28232,
    21938 => 28230,
    21939 => 28229,
    21940 => 28227,
    21941 => 28226,
    21942 => 28224,
    21943 => 28222,
    21944 => 28221,
    21945 => 28219,
    21946 => 28218,
    21947 => 28216,
    21948 => 28214,
    21949 => 28213,
    21950 => 28211,
    21951 => 28210,
    21952 => 28208,
    21953 => 28206,
    21954 => 28205,
    21955 => 28203,
    21956 => 28202,
    21957 => 28200,
    21958 => 28198,
    21959 => 28197,
    21960 => 28195,
    21961 => 28194,
    21962 => 28192,
    21963 => 28190,
    21964 => 28189,
    21965 => 28187,
    21966 => 28186,
    21967 => 28184,
    21968 => 28182,
    21969 => 28181,
    21970 => 28179,
    21971 => 28178,
    21972 => 28176,
    21973 => 28174,
    21974 => 28173,
    21975 => 28171,
    21976 => 28170,
    21977 => 28168,
    21978 => 28166,
    21979 => 28165,
    21980 => 28163,
    21981 => 28162,
    21982 => 28160,
    21983 => 28158,
    21984 => 28157,
    21985 => 28155,
    21986 => 28154,
    21987 => 28152,
    21988 => 28150,
    21989 => 28149,
    21990 => 28147,
    21991 => 28145,
    21992 => 28144,
    21993 => 28142,
    21994 => 28141,
    21995 => 28139,
    21996 => 28137,
    21997 => 28136,
    21998 => 28134,
    21999 => 28133,
    22000 => 28131,
    22001 => 28129,
    22002 => 28128,
    22003 => 28126,
    22004 => 28125,
    22005 => 28123,
    22006 => 28121,
    22007 => 28120,
    22008 => 28118,
    22009 => 28116,
    22010 => 28115,
    22011 => 28113,
    22012 => 28112,
    22013 => 28110,
    22014 => 28108,
    22015 => 28107,
    22016 => 28105,
    22017 => 28104,
    22018 => 28102,
    22019 => 28100,
    22020 => 28099,
    22021 => 28097,
    22022 => 28095,
    22023 => 28094,
    22024 => 28092,
    22025 => 28091,
    22026 => 28089,
    22027 => 28087,
    22028 => 28086,
    22029 => 28084,
    22030 => 28083,
    22031 => 28081,
    22032 => 28079,
    22033 => 28078,
    22034 => 28076,
    22035 => 28074,
    22036 => 28073,
    22037 => 28071,
    22038 => 28070,
    22039 => 28068,
    22040 => 28066,
    22041 => 28065,
    22042 => 28063,
    22043 => 28061,
    22044 => 28060,
    22045 => 28058,
    22046 => 28057,
    22047 => 28055,
    22048 => 28053,
    22049 => 28052,
    22050 => 28050,
    22051 => 28049,
    22052 => 28047,
    22053 => 28045,
    22054 => 28044,
    22055 => 28042,
    22056 => 28040,
    22057 => 28039,
    22058 => 28037,
    22059 => 28036,
    22060 => 28034,
    22061 => 28032,
    22062 => 28031,
    22063 => 28029,
    22064 => 28027,
    22065 => 28026,
    22066 => 28024,
    22067 => 28022,
    22068 => 28021,
    22069 => 28019,
    22070 => 28018,
    22071 => 28016,
    22072 => 28014,
    22073 => 28013,
    22074 => 28011,
    22075 => 28009,
    22076 => 28008,
    22077 => 28006,
    22078 => 28005,
    22079 => 28003,
    22080 => 28001,
    22081 => 28000,
    22082 => 27998,
    22083 => 27996,
    22084 => 27995,
    22085 => 27993,
    22086 => 27992,
    22087 => 27990,
    22088 => 27988,
    22089 => 27987,
    22090 => 27985,
    22091 => 27983,
    22092 => 27982,
    22093 => 27980,
    22094 => 27978,
    22095 => 27977,
    22096 => 27975,
    22097 => 27974,
    22098 => 27972,
    22099 => 27970,
    22100 => 27969,
    22101 => 27967,
    22102 => 27965,
    22103 => 27964,
    22104 => 27962,
    22105 => 27960,
    22106 => 27959,
    22107 => 27957,
    22108 => 27956,
    22109 => 27954,
    22110 => 27952,
    22111 => 27951,
    22112 => 27949,
    22113 => 27947,
    22114 => 27946,
    22115 => 27944,
    22116 => 27942,
    22117 => 27941,
    22118 => 27939,
    22119 => 27937,
    22120 => 27936,
    22121 => 27934,
    22122 => 27933,
    22123 => 27931,
    22124 => 27929,
    22125 => 27928,
    22126 => 27926,
    22127 => 27924,
    22128 => 27923,
    22129 => 27921,
    22130 => 27919,
    22131 => 27918,
    22132 => 27916,
    22133 => 27914,
    22134 => 27913,
    22135 => 27911,
    22136 => 27910,
    22137 => 27908,
    22138 => 27906,
    22139 => 27905,
    22140 => 27903,
    22141 => 27901,
    22142 => 27900,
    22143 => 27898,
    22144 => 27896,
    22145 => 27895,
    22146 => 27893,
    22147 => 27891,
    22148 => 27890,
    22149 => 27888,
    22150 => 27886,
    22151 => 27885,
    22152 => 27883,
    22153 => 27882,
    22154 => 27880,
    22155 => 27878,
    22156 => 27877,
    22157 => 27875,
    22158 => 27873,
    22159 => 27872,
    22160 => 27870,
    22161 => 27868,
    22162 => 27867,
    22163 => 27865,
    22164 => 27863,
    22165 => 27862,
    22166 => 27860,
    22167 => 27858,
    22168 => 27857,
    22169 => 27855,
    22170 => 27853,
    22171 => 27852,
    22172 => 27850,
    22173 => 27848,
    22174 => 27847,
    22175 => 27845,
    22176 => 27843,
    22177 => 27842,
    22178 => 27840,
    22179 => 27839,
    22180 => 27837,
    22181 => 27835,
    22182 => 27834,
    22183 => 27832,
    22184 => 27830,
    22185 => 27829,
    22186 => 27827,
    22187 => 27825,
    22188 => 27824,
    22189 => 27822,
    22190 => 27820,
    22191 => 27819,
    22192 => 27817,
    22193 => 27815,
    22194 => 27814,
    22195 => 27812,
    22196 => 27810,
    22197 => 27809,
    22198 => 27807,
    22199 => 27805,
    22200 => 27804,
    22201 => 27802,
    22202 => 27800,
    22203 => 27799,
    22204 => 27797,
    22205 => 27795,
    22206 => 27794,
    22207 => 27792,
    22208 => 27790,
    22209 => 27789,
    22210 => 27787,
    22211 => 27785,
    22212 => 27784,
    22213 => 27782,
    22214 => 27780,
    22215 => 27779,
    22216 => 27777,
    22217 => 27775,
    22218 => 27774,
    22219 => 27772,
    22220 => 27770,
    22221 => 27769,
    22222 => 27767,
    22223 => 27765,
    22224 => 27764,
    22225 => 27762,
    22226 => 27760,
    22227 => 27759,
    22228 => 27757,
    22229 => 27755,
    22230 => 27754,
    22231 => 27752,
    22232 => 27750,
    22233 => 27749,
    22234 => 27747,
    22235 => 27745,
    22236 => 27744,
    22237 => 27742,
    22238 => 27740,
    22239 => 27739,
    22240 => 27737,
    22241 => 27735,
    22242 => 27734,
    22243 => 27732,
    22244 => 27730,
    22245 => 27729,
    22246 => 27727,
    22247 => 27725,
    22248 => 27724,
    22249 => 27722,
    22250 => 27720,
    22251 => 27719,
    22252 => 27717,
    22253 => 27715,
    22254 => 27714,
    22255 => 27712,
    22256 => 27710,
    22257 => 27708,
    22258 => 27707,
    22259 => 27705,
    22260 => 27703,
    22261 => 27702,
    22262 => 27700,
    22263 => 27698,
    22264 => 27697,
    22265 => 27695,
    22266 => 27693,
    22267 => 27692,
    22268 => 27690,
    22269 => 27688,
    22270 => 27687,
    22271 => 27685,
    22272 => 27683,
    22273 => 27682,
    22274 => 27680,
    22275 => 27678,
    22276 => 27677,
    22277 => 27675,
    22278 => 27673,
    22279 => 27672,
    22280 => 27670,
    22281 => 27668,
    22282 => 27666,
    22283 => 27665,
    22284 => 27663,
    22285 => 27661,
    22286 => 27660,
    22287 => 27658,
    22288 => 27656,
    22289 => 27655,
    22290 => 27653,
    22291 => 27651,
    22292 => 27650,
    22293 => 27648,
    22294 => 27646,
    22295 => 27645,
    22296 => 27643,
    22297 => 27641,
    22298 => 27640,
    22299 => 27638,
    22300 => 27636,
    22301 => 27634,
    22302 => 27633,
    22303 => 27631,
    22304 => 27629,
    22305 => 27628,
    22306 => 27626,
    22307 => 27624,
    22308 => 27623,
    22309 => 27621,
    22310 => 27619,
    22311 => 27618,
    22312 => 27616,
    22313 => 27614,
    22314 => 27613,
    22315 => 27611,
    22316 => 27609,
    22317 => 27607,
    22318 => 27606,
    22319 => 27604,
    22320 => 27602,
    22321 => 27601,
    22322 => 27599,
    22323 => 27597,
    22324 => 27596,
    22325 => 27594,
    22326 => 27592,
    22327 => 27590,
    22328 => 27589,
    22329 => 27587,
    22330 => 27585,
    22331 => 27584,
    22332 => 27582,
    22333 => 27580,
    22334 => 27579,
    22335 => 27577,
    22336 => 27575,
    22337 => 27574,
    22338 => 27572,
    22339 => 27570,
    22340 => 27568,
    22341 => 27567,
    22342 => 27565,
    22343 => 27563,
    22344 => 27562,
    22345 => 27560,
    22346 => 27558,
    22347 => 27557,
    22348 => 27555,
    22349 => 27553,
    22350 => 27551,
    22351 => 27550,
    22352 => 27548,
    22353 => 27546,
    22354 => 27545,
    22355 => 27543,
    22356 => 27541,
    22357 => 27540,
    22358 => 27538,
    22359 => 27536,
    22360 => 27534,
    22361 => 27533,
    22362 => 27531,
    22363 => 27529,
    22364 => 27528,
    22365 => 27526,
    22366 => 27524,
    22367 => 27523,
    22368 => 27521,
    22369 => 27519,
    22370 => 27517,
    22371 => 27516,
    22372 => 27514,
    22373 => 27512,
    22374 => 27511,
    22375 => 27509,
    22376 => 27507,
    22377 => 27505,
    22378 => 27504,
    22379 => 27502,
    22380 => 27500,
    22381 => 27499,
    22382 => 27497,
    22383 => 27495,
    22384 => 27493,
    22385 => 27492,
    22386 => 27490,
    22387 => 27488,
    22388 => 27487,
    22389 => 27485,
    22390 => 27483,
    22391 => 27482,
    22392 => 27480,
    22393 => 27478,
    22394 => 27476,
    22395 => 27475,
    22396 => 27473,
    22397 => 27471,
    22398 => 27470,
    22399 => 27468,
    22400 => 27466,
    22401 => 27464,
    22402 => 27463,
    22403 => 27461,
    22404 => 27459,
    22405 => 27458,
    22406 => 27456,
    22407 => 27454,
    22408 => 27452,
    22409 => 27451,
    22410 => 27449,
    22411 => 27447,
    22412 => 27446,
    22413 => 27444,
    22414 => 27442,
    22415 => 27440,
    22416 => 27439,
    22417 => 27437,
    22418 => 27435,
    22419 => 27434,
    22420 => 27432,
    22421 => 27430,
    22422 => 27428,
    22423 => 27427,
    22424 => 27425,
    22425 => 27423,
    22426 => 27421,
    22427 => 27420,
    22428 => 27418,
    22429 => 27416,
    22430 => 27415,
    22431 => 27413,
    22432 => 27411,
    22433 => 27409,
    22434 => 27408,
    22435 => 27406,
    22436 => 27404,
    22437 => 27403,
    22438 => 27401,
    22439 => 27399,
    22440 => 27397,
    22441 => 27396,
    22442 => 27394,
    22443 => 27392,
    22444 => 27390,
    22445 => 27389,
    22446 => 27387,
    22447 => 27385,
    22448 => 27384,
    22449 => 27382,
    22450 => 27380,
    22451 => 27378,
    22452 => 27377,
    22453 => 27375,
    22454 => 27373,
    22455 => 27372,
    22456 => 27370,
    22457 => 27368,
    22458 => 27366,
    22459 => 27365,
    22460 => 27363,
    22461 => 27361,
    22462 => 27359,
    22463 => 27358,
    22464 => 27356,
    22465 => 27354,
    22466 => 27352,
    22467 => 27351,
    22468 => 27349,
    22469 => 27347,
    22470 => 27346,
    22471 => 27344,
    22472 => 27342,
    22473 => 27340,
    22474 => 27339,
    22475 => 27337,
    22476 => 27335,
    22477 => 27333,
    22478 => 27332,
    22479 => 27330,
    22480 => 27328,
    22481 => 27327,
    22482 => 27325,
    22483 => 27323,
    22484 => 27321,
    22485 => 27320,
    22486 => 27318,
    22487 => 27316,
    22488 => 27314,
    22489 => 27313,
    22490 => 27311,
    22491 => 27309,
    22492 => 27307,
    22493 => 27306,
    22494 => 27304,
    22495 => 27302,
    22496 => 27300,
    22497 => 27299,
    22498 => 27297,
    22499 => 27295,
    22500 => 27294,
    22501 => 27292,
    22502 => 27290,
    22503 => 27288,
    22504 => 27287,
    22505 => 27285,
    22506 => 27283,
    22507 => 27281,
    22508 => 27280,
    22509 => 27278,
    22510 => 27276,
    22511 => 27274,
    22512 => 27273,
    22513 => 27271,
    22514 => 27269,
    22515 => 27267,
    22516 => 27266,
    22517 => 27264,
    22518 => 27262,
    22519 => 27260,
    22520 => 27259,
    22521 => 27257,
    22522 => 27255,
    22523 => 27253,
    22524 => 27252,
    22525 => 27250,
    22526 => 27248,
    22527 => 27247,
    22528 => 27245,
    22529 => 27243,
    22530 => 27241,
    22531 => 27240,
    22532 => 27238,
    22533 => 27236,
    22534 => 27234,
    22535 => 27233,
    22536 => 27231,
    22537 => 27229,
    22538 => 27227,
    22539 => 27226,
    22540 => 27224,
    22541 => 27222,
    22542 => 27220,
    22543 => 27219,
    22544 => 27217,
    22545 => 27215,
    22546 => 27213,
    22547 => 27212,
    22548 => 27210,
    22549 => 27208,
    22550 => 27206,
    22551 => 27205,
    22552 => 27203,
    22553 => 27201,
    22554 => 27199,
    22555 => 27198,
    22556 => 27196,
    22557 => 27194,
    22558 => 27192,
    22559 => 27191,
    22560 => 27189,
    22561 => 27187,
    22562 => 27185,
    22563 => 27184,
    22564 => 27182,
    22565 => 27180,
    22566 => 27178,
    22567 => 27177,
    22568 => 27175,
    22569 => 27173,
    22570 => 27171,
    22571 => 27169,
    22572 => 27168,
    22573 => 27166,
    22574 => 27164,
    22575 => 27162,
    22576 => 27161,
    22577 => 27159,
    22578 => 27157,
    22579 => 27155,
    22580 => 27154,
    22581 => 27152,
    22582 => 27150,
    22583 => 27148,
    22584 => 27147,
    22585 => 27145,
    22586 => 27143,
    22587 => 27141,
    22588 => 27140,
    22589 => 27138,
    22590 => 27136,
    22591 => 27134,
    22592 => 27133,
    22593 => 27131,
    22594 => 27129,
    22595 => 27127,
    22596 => 27126,
    22597 => 27124,
    22598 => 27122,
    22599 => 27120,
    22600 => 27118,
    22601 => 27117,
    22602 => 27115,
    22603 => 27113,
    22604 => 27111,
    22605 => 27110,
    22606 => 27108,
    22607 => 27106,
    22608 => 27104,
    22609 => 27103,
    22610 => 27101,
    22611 => 27099,
    22612 => 27097,
    22613 => 27096,
    22614 => 27094,
    22615 => 27092,
    22616 => 27090,
    22617 => 27088,
    22618 => 27087,
    22619 => 27085,
    22620 => 27083,
    22621 => 27081,
    22622 => 27080,
    22623 => 27078,
    22624 => 27076,
    22625 => 27074,
    22626 => 27073,
    22627 => 27071,
    22628 => 27069,
    22629 => 27067,
    22630 => 27065,
    22631 => 27064,
    22632 => 27062,
    22633 => 27060,
    22634 => 27058,
    22635 => 27057,
    22636 => 27055,
    22637 => 27053,
    22638 => 27051,
    22639 => 27049,
    22640 => 27048,
    22641 => 27046,
    22642 => 27044,
    22643 => 27042,
    22644 => 27041,
    22645 => 27039,
    22646 => 27037,
    22647 => 27035,
    22648 => 27034,
    22649 => 27032,
    22650 => 27030,
    22651 => 27028,
    22652 => 27026,
    22653 => 27025,
    22654 => 27023,
    22655 => 27021,
    22656 => 27019,
    22657 => 27018,
    22658 => 27016,
    22659 => 27014,
    22660 => 27012,
    22661 => 27010,
    22662 => 27009,
    22663 => 27007,
    22664 => 27005,
    22665 => 27003,
    22666 => 27002,
    22667 => 27000,
    22668 => 26998,
    22669 => 26996,
    22670 => 26994,
    22671 => 26993,
    22672 => 26991,
    22673 => 26989,
    22674 => 26987,
    22675 => 26986,
    22676 => 26984,
    22677 => 26982,
    22678 => 26980,
    22679 => 26978,
    22680 => 26977,
    22681 => 26975,
    22682 => 26973,
    22683 => 26971,
    22684 => 26969,
    22685 => 26968,
    22686 => 26966,
    22687 => 26964,
    22688 => 26962,
    22689 => 26961,
    22690 => 26959,
    22691 => 26957,
    22692 => 26955,
    22693 => 26953,
    22694 => 26952,
    22695 => 26950,
    22696 => 26948,
    22697 => 26946,
    22698 => 26944,
    22699 => 26943,
    22700 => 26941,
    22701 => 26939,
    22702 => 26937,
    22703 => 26936,
    22704 => 26934,
    22705 => 26932,
    22706 => 26930,
    22707 => 26928,
    22708 => 26927,
    22709 => 26925,
    22710 => 26923,
    22711 => 26921,
    22712 => 26919,
    22713 => 26918,
    22714 => 26916,
    22715 => 26914,
    22716 => 26912,
    22717 => 26910,
    22718 => 26909,
    22719 => 26907,
    22720 => 26905,
    22721 => 26903,
    22722 => 26901,
    22723 => 26900,
    22724 => 26898,
    22725 => 26896,
    22726 => 26894,
    22727 => 26893,
    22728 => 26891,
    22729 => 26889,
    22730 => 26887,
    22731 => 26885,
    22732 => 26884,
    22733 => 26882,
    22734 => 26880,
    22735 => 26878,
    22736 => 26876,
    22737 => 26875,
    22738 => 26873,
    22739 => 26871,
    22740 => 26869,
    22741 => 26867,
    22742 => 26866,
    22743 => 26864,
    22744 => 26862,
    22745 => 26860,
    22746 => 26858,
    22747 => 26857,
    22748 => 26855,
    22749 => 26853,
    22750 => 26851,
    22751 => 26849,
    22752 => 26848,
    22753 => 26846,
    22754 => 26844,
    22755 => 26842,
    22756 => 26840,
    22757 => 26839,
    22758 => 26837,
    22759 => 26835,
    22760 => 26833,
    22761 => 26831,
    22762 => 26830,
    22763 => 26828,
    22764 => 26826,
    22765 => 26824,
    22766 => 26822,
    22767 => 26821,
    22768 => 26819,
    22769 => 26817,
    22770 => 26815,
    22771 => 26813,
    22772 => 26811,
    22773 => 26810,
    22774 => 26808,
    22775 => 26806,
    22776 => 26804,
    22777 => 26802,
    22778 => 26801,
    22779 => 26799,
    22780 => 26797,
    22781 => 26795,
    22782 => 26793,
    22783 => 26792,
    22784 => 26790,
    22785 => 26788,
    22786 => 26786,
    22787 => 26784,
    22788 => 26783,
    22789 => 26781,
    22790 => 26779,
    22791 => 26777,
    22792 => 26775,
    22793 => 26774,
    22794 => 26772,
    22795 => 26770,
    22796 => 26768,
    22797 => 26766,
    22798 => 26764,
    22799 => 26763,
    22800 => 26761,
    22801 => 26759,
    22802 => 26757,
    22803 => 26755,
    22804 => 26754,
    22805 => 26752,
    22806 => 26750,
    22807 => 26748,
    22808 => 26746,
    22809 => 26745,
    22810 => 26743,
    22811 => 26741,
    22812 => 26739,
    22813 => 26737,
    22814 => 26735,
    22815 => 26734,
    22816 => 26732,
    22817 => 26730,
    22818 => 26728,
    22819 => 26726,
    22820 => 26725,
    22821 => 26723,
    22822 => 26721,
    22823 => 26719,
    22824 => 26717,
    22825 => 26715,
    22826 => 26714,
    22827 => 26712,
    22828 => 26710,
    22829 => 26708,
    22830 => 26706,
    22831 => 26705,
    22832 => 26703,
    22833 => 26701,
    22834 => 26699,
    22835 => 26697,
    22836 => 26695,
    22837 => 26694,
    22838 => 26692,
    22839 => 26690,
    22840 => 26688,
    22841 => 26686,
    22842 => 26684,
    22843 => 26683,
    22844 => 26681,
    22845 => 26679,
    22846 => 26677,
    22847 => 26675,
    22848 => 26674,
    22849 => 26672,
    22850 => 26670,
    22851 => 26668,
    22852 => 26666,
    22853 => 26664,
    22854 => 26663,
    22855 => 26661,
    22856 => 26659,
    22857 => 26657,
    22858 => 26655,
    22859 => 26653,
    22860 => 26652,
    22861 => 26650,
    22862 => 26648,
    22863 => 26646,
    22864 => 26644,
    22865 => 26642,
    22866 => 26641,
    22867 => 26639,
    22868 => 26637,
    22869 => 26635,
    22870 => 26633,
    22871 => 26631,
    22872 => 26630,
    22873 => 26628,
    22874 => 26626,
    22875 => 26624,
    22876 => 26622,
    22877 => 26621,
    22878 => 26619,
    22879 => 26617,
    22880 => 26615,
    22881 => 26613,
    22882 => 26611,
    22883 => 26610,
    22884 => 26608,
    22885 => 26606,
    22886 => 26604,
    22887 => 26602,
    22888 => 26600,
    22889 => 26599,
    22890 => 26597,
    22891 => 26595,
    22892 => 26593,
    22893 => 26591,
    22894 => 26589,
    22895 => 26588,
    22896 => 26586,
    22897 => 26584,
    22898 => 26582,
    22899 => 26580,
    22900 => 26578,
    22901 => 26576,
    22902 => 26575,
    22903 => 26573,
    22904 => 26571,
    22905 => 26569,
    22906 => 26567,
    22907 => 26565,
    22908 => 26564,
    22909 => 26562,
    22910 => 26560,
    22911 => 26558,
    22912 => 26556,
    22913 => 26554,
    22914 => 26553,
    22915 => 26551,
    22916 => 26549,
    22917 => 26547,
    22918 => 26545,
    22919 => 26543,
    22920 => 26542,
    22921 => 26540,
    22922 => 26538,
    22923 => 26536,
    22924 => 26534,
    22925 => 26532,
    22926 => 26530,
    22927 => 26529,
    22928 => 26527,
    22929 => 26525,
    22930 => 26523,
    22931 => 26521,
    22932 => 26519,
    22933 => 26518,
    22934 => 26516,
    22935 => 26514,
    22936 => 26512,
    22937 => 26510,
    22938 => 26508,
    22939 => 26506,
    22940 => 26505,
    22941 => 26503,
    22942 => 26501,
    22943 => 26499,
    22944 => 26497,
    22945 => 26495,
    22946 => 26494,
    22947 => 26492,
    22948 => 26490,
    22949 => 26488,
    22950 => 26486,
    22951 => 26484,
    22952 => 26482,
    22953 => 26481,
    22954 => 26479,
    22955 => 26477,
    22956 => 26475,
    22957 => 26473,
    22958 => 26471,
    22959 => 26469,
    22960 => 26468,
    22961 => 26466,
    22962 => 26464,
    22963 => 26462,
    22964 => 26460,
    22965 => 26458,
    22966 => 26457,
    22967 => 26455,
    22968 => 26453,
    22969 => 26451,
    22970 => 26449,
    22971 => 26447,
    22972 => 26445,
    22973 => 26444,
    22974 => 26442,
    22975 => 26440,
    22976 => 26438,
    22977 => 26436,
    22978 => 26434,
    22979 => 26432,
    22980 => 26431,
    22981 => 26429,
    22982 => 26427,
    22983 => 26425,
    22984 => 26423,
    22985 => 26421,
    22986 => 26419,
    22987 => 26418,
    22988 => 26416,
    22989 => 26414,
    22990 => 26412,
    22991 => 26410,
    22992 => 26408,
    22993 => 26406,
    22994 => 26405,
    22995 => 26403,
    22996 => 26401,
    22997 => 26399,
    22998 => 26397,
    22999 => 26395,
    23000 => 26393,
    23001 => 26392,
    23002 => 26390,
    23003 => 26388,
    23004 => 26386,
    23005 => 26384,
    23006 => 26382,
    23007 => 26380,
    23008 => 26378,
    23009 => 26377,
    23010 => 26375,
    23011 => 26373,
    23012 => 26371,
    23013 => 26369,
    23014 => 26367,
    23015 => 26365,
    23016 => 26364,
    23017 => 26362,
    23018 => 26360,
    23019 => 26358,
    23020 => 26356,
    23021 => 26354,
    23022 => 26352,
    23023 => 26350,
    23024 => 26349,
    23025 => 26347,
    23026 => 26345,
    23027 => 26343,
    23028 => 26341,
    23029 => 26339,
    23030 => 26337,
    23031 => 26336,
    23032 => 26334,
    23033 => 26332,
    23034 => 26330,
    23035 => 26328,
    23036 => 26326,
    23037 => 26324,
    23038 => 26322,
    23039 => 26321,
    23040 => 26319,
    23041 => 26317,
    23042 => 26315,
    23043 => 26313,
    23044 => 26311,
    23045 => 26309,
    23046 => 26307,
    23047 => 26306,
    23048 => 26304,
    23049 => 26302,
    23050 => 26300,
    23051 => 26298,
    23052 => 26296,
    23053 => 26294,
    23054 => 26292,
    23055 => 26291,
    23056 => 26289,
    23057 => 26287,
    23058 => 26285,
    23059 => 26283,
    23060 => 26281,
    23061 => 26279,
    23062 => 26277,
    23063 => 26276,
    23064 => 26274,
    23065 => 26272,
    23066 => 26270,
    23067 => 26268,
    23068 => 26266,
    23069 => 26264,
    23070 => 26262,
    23071 => 26261,
    23072 => 26259,
    23073 => 26257,
    23074 => 26255,
    23075 => 26253,
    23076 => 26251,
    23077 => 26249,
    23078 => 26247,
    23079 => 26246,
    23080 => 26244,
    23081 => 26242,
    23082 => 26240,
    23083 => 26238,
    23084 => 26236,
    23085 => 26234,
    23086 => 26232,
    23087 => 26230,
    23088 => 26229,
    23089 => 26227,
    23090 => 26225,
    23091 => 26223,
    23092 => 26221,
    23093 => 26219,
    23094 => 26217,
    23095 => 26215,
    23096 => 26214,
    23097 => 26212,
    23098 => 26210,
    23099 => 26208,
    23100 => 26206,
    23101 => 26204,
    23102 => 26202,
    23103 => 26200,
    23104 => 26198,
    23105 => 26197,
    23106 => 26195,
    23107 => 26193,
    23108 => 26191,
    23109 => 26189,
    23110 => 26187,
    23111 => 26185,
    23112 => 26183,
    23113 => 26181,
    23114 => 26180,
    23115 => 26178,
    23116 => 26176,
    23117 => 26174,
    23118 => 26172,
    23119 => 26170,
    23120 => 26168,
    23121 => 26166,
    23122 => 26164,
    23123 => 26163,
    23124 => 26161,
    23125 => 26159,
    23126 => 26157,
    23127 => 26155,
    23128 => 26153,
    23129 => 26151,
    23130 => 26149,
    23131 => 26147,
    23132 => 26146,
    23133 => 26144,
    23134 => 26142,
    23135 => 26140,
    23136 => 26138,
    23137 => 26136,
    23138 => 26134,
    23139 => 26132,
    23140 => 26130,
    23141 => 26128,
    23142 => 26127,
    23143 => 26125,
    23144 => 26123,
    23145 => 26121,
    23146 => 26119,
    23147 => 26117,
    23148 => 26115,
    23149 => 26113,
    23150 => 26111,
    23151 => 26109,
    23152 => 26108,
    23153 => 26106,
    23154 => 26104,
    23155 => 26102,
    23156 => 26100,
    23157 => 26098,
    23158 => 26096,
    23159 => 26094,
    23160 => 26092,
    23161 => 26090,
    23162 => 26089,
    23163 => 26087,
    23164 => 26085,
    23165 => 26083,
    23166 => 26081,
    23167 => 26079,
    23168 => 26077,
    23169 => 26075,
    23170 => 26073,
    23171 => 26071,
    23172 => 26070,
    23173 => 26068,
    23174 => 26066,
    23175 => 26064,
    23176 => 26062,
    23177 => 26060,
    23178 => 26058,
    23179 => 26056,
    23180 => 26054,
    23181 => 26052,
    23182 => 26051,
    23183 => 26049,
    23184 => 26047,
    23185 => 26045,
    23186 => 26043,
    23187 => 26041,
    23188 => 26039,
    23189 => 26037,
    23190 => 26035,
    23191 => 26033,
    23192 => 26031,
    23193 => 26030,
    23194 => 26028,
    23195 => 26026,
    23196 => 26024,
    23197 => 26022,
    23198 => 26020,
    23199 => 26018,
    23200 => 26016,
    23201 => 26014,
    23202 => 26012,
    23203 => 26010,
    23204 => 26009,
    23205 => 26007,
    23206 => 26005,
    23207 => 26003,
    23208 => 26001,
    23209 => 25999,
    23210 => 25997,
    23211 => 25995,
    23212 => 25993,
    23213 => 25991,
    23214 => 25989,
    23215 => 25988,
    23216 => 25986,
    23217 => 25984,
    23218 => 25982,
    23219 => 25980,
    23220 => 25978,
    23221 => 25976,
    23222 => 25974,
    23223 => 25972,
    23224 => 25970,
    23225 => 25968,
    23226 => 25966,
    23227 => 25965,
    23228 => 25963,
    23229 => 25961,
    23230 => 25959,
    23231 => 25957,
    23232 => 25955,
    23233 => 25953,
    23234 => 25951,
    23235 => 25949,
    23236 => 25947,
    23237 => 25945,
    23238 => 25943,
    23239 => 25942,
    23240 => 25940,
    23241 => 25938,
    23242 => 25936,
    23243 => 25934,
    23244 => 25932,
    23245 => 25930,
    23246 => 25928,
    23247 => 25926,
    23248 => 25924,
    23249 => 25922,
    23250 => 25920,
    23251 => 25918,
    23252 => 25917,
    23253 => 25915,
    23254 => 25913,
    23255 => 25911,
    23256 => 25909,
    23257 => 25907,
    23258 => 25905,
    23259 => 25903,
    23260 => 25901,
    23261 => 25899,
    23262 => 25897,
    23263 => 25895,
    23264 => 25893,
    23265 => 25892,
    23266 => 25890,
    23267 => 25888,
    23268 => 25886,
    23269 => 25884,
    23270 => 25882,
    23271 => 25880,
    23272 => 25878,
    23273 => 25876,
    23274 => 25874,
    23275 => 25872,
    23276 => 25870,
    23277 => 25868,
    23278 => 25866,
    23279 => 25865,
    23280 => 25863,
    23281 => 25861,
    23282 => 25859,
    23283 => 25857,
    23284 => 25855,
    23285 => 25853,
    23286 => 25851,
    23287 => 25849,
    23288 => 25847,
    23289 => 25845,
    23290 => 25843,
    23291 => 25841,
    23292 => 25839,
    23293 => 25838,
    23294 => 25836,
    23295 => 25834,
    23296 => 25832,
    23297 => 25830,
    23298 => 25828,
    23299 => 25826,
    23300 => 25824,
    23301 => 25822,
    23302 => 25820,
    23303 => 25818,
    23304 => 25816,
    23305 => 25814,
    23306 => 25812,
    23307 => 25810,
    23308 => 25809,
    23309 => 25807,
    23310 => 25805,
    23311 => 25803,
    23312 => 25801,
    23313 => 25799,
    23314 => 25797,
    23315 => 25795,
    23316 => 25793,
    23317 => 25791,
    23318 => 25789,
    23319 => 25787,
    23320 => 25785,
    23321 => 25783,
    23322 => 25781,
    23323 => 25779,
    23324 => 25778,
    23325 => 25776,
    23326 => 25774,
    23327 => 25772,
    23328 => 25770,
    23329 => 25768,
    23330 => 25766,
    23331 => 25764,
    23332 => 25762,
    23333 => 25760,
    23334 => 25758,
    23335 => 25756,
    23336 => 25754,
    23337 => 25752,
    23338 => 25750,
    23339 => 25748,
    23340 => 25746,
    23341 => 25745,
    23342 => 25743,
    23343 => 25741,
    23344 => 25739,
    23345 => 25737,
    23346 => 25735,
    23347 => 25733,
    23348 => 25731,
    23349 => 25729,
    23350 => 25727,
    23351 => 25725,
    23352 => 25723,
    23353 => 25721,
    23354 => 25719,
    23355 => 25717,
    23356 => 25715,
    23357 => 25713,
    23358 => 25711,
    23359 => 25710,
    23360 => 25708,
    23361 => 25706,
    23362 => 25704,
    23363 => 25702,
    23364 => 25700,
    23365 => 25698,
    23366 => 25696,
    23367 => 25694,
    23368 => 25692,
    23369 => 25690,
    23370 => 25688,
    23371 => 25686,
    23372 => 25684,
    23373 => 25682,
    23374 => 25680,
    23375 => 25678,
    23376 => 25676,
    23377 => 25674,
    23378 => 25672,
    23379 => 25671,
    23380 => 25669,
    23381 => 25667,
    23382 => 25665,
    23383 => 25663,
    23384 => 25661,
    23385 => 25659,
    23386 => 25657,
    23387 => 25655,
    23388 => 25653,
    23389 => 25651,
    23390 => 25649,
    23391 => 25647,
    23392 => 25645,
    23393 => 25643,
    23394 => 25641,
    23395 => 25639,
    23396 => 25637,
    23397 => 25635,
    23398 => 25633,
    23399 => 25631,
    23400 => 25629,
    23401 => 25628,
    23402 => 25626,
    23403 => 25624,
    23404 => 25622,
    23405 => 25620,
    23406 => 25618,
    23407 => 25616,
    23408 => 25614,
    23409 => 25612,
    23410 => 25610,
    23411 => 25608,
    23412 => 25606,
    23413 => 25604,
    23414 => 25602,
    23415 => 25600,
    23416 => 25598,
    23417 => 25596,
    23418 => 25594,
    23419 => 25592,
    23420 => 25590,
    23421 => 25588,
    23422 => 25586,
    23423 => 25584,
    23424 => 25582,
    23425 => 25580,
    23426 => 25578,
    23427 => 25577,
    23428 => 25575,
    23429 => 25573,
    23430 => 25571,
    23431 => 25569,
    23432 => 25567,
    23433 => 25565,
    23434 => 25563,
    23435 => 25561,
    23436 => 25559,
    23437 => 25557,
    23438 => 25555,
    23439 => 25553,
    23440 => 25551,
    23441 => 25549,
    23442 => 25547,
    23443 => 25545,
    23444 => 25543,
    23445 => 25541,
    23446 => 25539,
    23447 => 25537,
    23448 => 25535,
    23449 => 25533,
    23450 => 25531,
    23451 => 25529,
    23452 => 25527,
    23453 => 25525,
    23454 => 25523,
    23455 => 25521,
    23456 => 25519,
    23457 => 25518,
    23458 => 25516,
    23459 => 25514,
    23460 => 25512,
    23461 => 25510,
    23462 => 25508,
    23463 => 25506,
    23464 => 25504,
    23465 => 25502,
    23466 => 25500,
    23467 => 25498,
    23468 => 25496,
    23469 => 25494,
    23470 => 25492,
    23471 => 25490,
    23472 => 25488,
    23473 => 25486,
    23474 => 25484,
    23475 => 25482,
    23476 => 25480,
    23477 => 25478,
    23478 => 25476,
    23479 => 25474,
    23480 => 25472,
    23481 => 25470,
    23482 => 25468,
    23483 => 25466,
    23484 => 25464,
    23485 => 25462,
    23486 => 25460,
    23487 => 25458,
    23488 => 25456,
    23489 => 25454,
    23490 => 25452,
    23491 => 25450,
    23492 => 25448,
    23493 => 25446,
    23494 => 25444,
    23495 => 25442,
    23496 => 25440,
    23497 => 25438,
    23498 => 25437,
    23499 => 25435,
    23500 => 25433,
    23501 => 25431,
    23502 => 25429,
    23503 => 25427,
    23504 => 25425,
    23505 => 25423,
    23506 => 25421,
    23507 => 25419,
    23508 => 25417,
    23509 => 25415,
    23510 => 25413,
    23511 => 25411,
    23512 => 25409,
    23513 => 25407,
    23514 => 25405,
    23515 => 25403,
    23516 => 25401,
    23517 => 25399,
    23518 => 25397,
    23519 => 25395,
    23520 => 25393,
    23521 => 25391,
    23522 => 25389,
    23523 => 25387,
    23524 => 25385,
    23525 => 25383,
    23526 => 25381,
    23527 => 25379,
    23528 => 25377,
    23529 => 25375,
    23530 => 25373,
    23531 => 25371,
    23532 => 25369,
    23533 => 25367,
    23534 => 25365,
    23535 => 25363,
    23536 => 25361,
    23537 => 25359,
    23538 => 25357,
    23539 => 25355,
    23540 => 25353,
    23541 => 25351,
    23542 => 25349,
    23543 => 25347,
    23544 => 25345,
    23545 => 25343,
    23546 => 25341,
    23547 => 25339,
    23548 => 25337,
    23549 => 25335,
    23550 => 25333,
    23551 => 25331,
    23552 => 25329,
    23553 => 25327,
    23554 => 25325,
    23555 => 25323,
    23556 => 25321,
    23557 => 25319,
    23558 => 25317,
    23559 => 25315,
    23560 => 25313,
    23561 => 25311,
    23562 => 25309,
    23563 => 25307,
    23564 => 25305,
    23565 => 25303,
    23566 => 25301,
    23567 => 25299,
    23568 => 25297,
    23569 => 25295,
    23570 => 25293,
    23571 => 25291,
    23572 => 25289,
    23573 => 25287,
    23574 => 25285,
    23575 => 25283,
    23576 => 25281,
    23577 => 25279,
    23578 => 25277,
    23579 => 25275,
    23580 => 25273,
    23581 => 25271,
    23582 => 25269,
    23583 => 25267,
    23584 => 25265,
    23585 => 25263,
    23586 => 25261,
    23587 => 25259,
    23588 => 25257,
    23589 => 25255,
    23590 => 25253,
    23591 => 25251,
    23592 => 25249,
    23593 => 25247,
    23594 => 25245,
    23595 => 25243,
    23596 => 25241,
    23597 => 25239,
    23598 => 25237,
    23599 => 25235,
    23600 => 25233,
    23601 => 25231,
    23602 => 25229,
    23603 => 25227,
    23604 => 25225,
    23605 => 25223,
    23606 => 25221,
    23607 => 25219,
    23608 => 25217,
    23609 => 25215,
    23610 => 25213,
    23611 => 25211,
    23612 => 25209,
    23613 => 25207,
    23614 => 25205,
    23615 => 25203,
    23616 => 25201,
    23617 => 25199,
    23618 => 25197,
    23619 => 25195,
    23620 => 25193,
    23621 => 25191,
    23622 => 25189,
    23623 => 25187,
    23624 => 25185,
    23625 => 25183,
    23626 => 25181,
    23627 => 25179,
    23628 => 25177,
    23629 => 25175,
    23630 => 25173,
    23631 => 25171,
    23632 => 25169,
    23633 => 25167,
    23634 => 25165,
    23635 => 25163,
    23636 => 25161,
    23637 => 25159,
    23638 => 25157,
    23639 => 25155,
    23640 => 25153,
    23641 => 25151,
    23642 => 25149,
    23643 => 25147,
    23644 => 25145,
    23645 => 25143,
    23646 => 25141,
    23647 => 25139,
    23648 => 25137,
    23649 => 25135,
    23650 => 25133,
    23651 => 25131,
    23652 => 25129,
    23653 => 25127,
    23654 => 25125,
    23655 => 25123,
    23656 => 25121,
    23657 => 25119,
    23658 => 25117,
    23659 => 25115,
    23660 => 25113,
    23661 => 25111,
    23662 => 25109,
    23663 => 25107,
    23664 => 25105,
    23665 => 25103,
    23666 => 25101,
    23667 => 25099,
    23668 => 25096,
    23669 => 25094,
    23670 => 25092,
    23671 => 25090,
    23672 => 25088,
    23673 => 25086,
    23674 => 25084,
    23675 => 25082,
    23676 => 25080,
    23677 => 25078,
    23678 => 25076,
    23679 => 25074,
    23680 => 25072,
    23681 => 25070,
    23682 => 25068,
    23683 => 25066,
    23684 => 25064,
    23685 => 25062,
    23686 => 25060,
    23687 => 25058,
    23688 => 25056,
    23689 => 25054,
    23690 => 25052,
    23691 => 25050,
    23692 => 25048,
    23693 => 25046,
    23694 => 25044,
    23695 => 25042,
    23696 => 25040,
    23697 => 25038,
    23698 => 25036,
    23699 => 25034,
    23700 => 25032,
    23701 => 25030,
    23702 => 25028,
    23703 => 25026,
    23704 => 25024,
    23705 => 25022,
    23706 => 25020,
    23707 => 25018,
    23708 => 25016,
    23709 => 25013,
    23710 => 25011,
    23711 => 25009,
    23712 => 25007,
    23713 => 25005,
    23714 => 25003,
    23715 => 25001,
    23716 => 24999,
    23717 => 24997,
    23718 => 24995,
    23719 => 24993,
    23720 => 24991,
    23721 => 24989,
    23722 => 24987,
    23723 => 24985,
    23724 => 24983,
    23725 => 24981,
    23726 => 24979,
    23727 => 24977,
    23728 => 24975,
    23729 => 24973,
    23730 => 24971,
    23731 => 24969,
    23732 => 24967,
    23733 => 24965,
    23734 => 24963,
    23735 => 24961,
    23736 => 24959,
    23737 => 24957,
    23738 => 24955,
    23739 => 24953,
    23740 => 24950,
    23741 => 24948,
    23742 => 24946,
    23743 => 24944,
    23744 => 24942,
    23745 => 24940,
    23746 => 24938,
    23747 => 24936,
    23748 => 24934,
    23749 => 24932,
    23750 => 24930,
    23751 => 24928,
    23752 => 24926,
    23753 => 24924,
    23754 => 24922,
    23755 => 24920,
    23756 => 24918,
    23757 => 24916,
    23758 => 24914,
    23759 => 24912,
    23760 => 24910,
    23761 => 24908,
    23762 => 24906,
    23763 => 24904,
    23764 => 24902,
    23765 => 24899,
    23766 => 24897,
    23767 => 24895,
    23768 => 24893,
    23769 => 24891,
    23770 => 24889,
    23771 => 24887,
    23772 => 24885,
    23773 => 24883,
    23774 => 24881,
    23775 => 24879,
    23776 => 24877,
    23777 => 24875,
    23778 => 24873,
    23779 => 24871,
    23780 => 24869,
    23781 => 24867,
    23782 => 24865,
    23783 => 24863,
    23784 => 24861,
    23785 => 24859,
    23786 => 24857,
    23787 => 24855,
    23788 => 24852,
    23789 => 24850,
    23790 => 24848,
    23791 => 24846,
    23792 => 24844,
    23793 => 24842,
    23794 => 24840,
    23795 => 24838,
    23796 => 24836,
    23797 => 24834,
    23798 => 24832,
    23799 => 24830,
    23800 => 24828,
    23801 => 24826,
    23802 => 24824,
    23803 => 24822,
    23804 => 24820,
    23805 => 24818,
    23806 => 24816,
    23807 => 24814,
    23808 => 24811,
    23809 => 24809,
    23810 => 24807,
    23811 => 24805,
    23812 => 24803,
    23813 => 24801,
    23814 => 24799,
    23815 => 24797,
    23816 => 24795,
    23817 => 24793,
    23818 => 24791,
    23819 => 24789,
    23820 => 24787,
    23821 => 24785,
    23822 => 24783,
    23823 => 24781,
    23824 => 24779,
    23825 => 24777,
    23826 => 24774,
    23827 => 24772,
    23828 => 24770,
    23829 => 24768,
    23830 => 24766,
    23831 => 24764,
    23832 => 24762,
    23833 => 24760,
    23834 => 24758,
    23835 => 24756,
    23836 => 24754,
    23837 => 24752,
    23838 => 24750,
    23839 => 24748,
    23840 => 24746,
    23841 => 24744,
    23842 => 24742,
    23843 => 24740,
    23844 => 24737,
    23845 => 24735,
    23846 => 24733,
    23847 => 24731,
    23848 => 24729,
    23849 => 24727,
    23850 => 24725,
    23851 => 24723,
    23852 => 24721,
    23853 => 24719,
    23854 => 24717,
    23855 => 24715,
    23856 => 24713,
    23857 => 24711,
    23858 => 24709,
    23859 => 24707,
    23860 => 24704,
    23861 => 24702,
    23862 => 24700,
    23863 => 24698,
    23864 => 24696,
    23865 => 24694,
    23866 => 24692,
    23867 => 24690,
    23868 => 24688,
    23869 => 24686,
    23870 => 24684,
    23871 => 24682,
    23872 => 24680,
    23873 => 24678,
    23874 => 24676,
    23875 => 24673,
    23876 => 24671,
    23877 => 24669,
    23878 => 24667,
    23879 => 24665,
    23880 => 24663,
    23881 => 24661,
    23882 => 24659,
    23883 => 24657,
    23884 => 24655,
    23885 => 24653,
    23886 => 24651,
    23887 => 24649,
    23888 => 24647,
    23889 => 24645,
    23890 => 24642,
    23891 => 24640,
    23892 => 24638,
    23893 => 24636,
    23894 => 24634,
    23895 => 24632,
    23896 => 24630,
    23897 => 24628,
    23898 => 24626,
    23899 => 24624,
    23900 => 24622,
    23901 => 24620,
    23902 => 24618,
    23903 => 24616,
    23904 => 24613,
    23905 => 24611,
    23906 => 24609,
    23907 => 24607,
    23908 => 24605,
    23909 => 24603,
    23910 => 24601,
    23911 => 24599,
    23912 => 24597,
    23913 => 24595,
    23914 => 24593,
    23915 => 24591,
    23916 => 24589,
    23917 => 24586,
    23918 => 24584,
    23919 => 24582,
    23920 => 24580,
    23921 => 24578,
    23922 => 24576,
    23923 => 24574,
    23924 => 24572,
    23925 => 24570,
    23926 => 24568,
    23927 => 24566,
    23928 => 24564,
    23929 => 24562,
    23930 => 24559,
    23931 => 24557,
    23932 => 24555,
    23933 => 24553,
    23934 => 24551,
    23935 => 24549,
    23936 => 24547,
    23937 => 24545,
    23938 => 24543,
    23939 => 24541,
    23940 => 24539,
    23941 => 24537,
    23942 => 24534,
    23943 => 24532,
    23944 => 24530,
    23945 => 24528,
    23946 => 24526,
    23947 => 24524,
    23948 => 24522,
    23949 => 24520,
    23950 => 24518,
    23951 => 24516,
    23952 => 24514,
    23953 => 24512,
    23954 => 24509,
    23955 => 24507,
    23956 => 24505,
    23957 => 24503,
    23958 => 24501,
    23959 => 24499,
    23960 => 24497,
    23961 => 24495,
    23962 => 24493,
    23963 => 24491,
    23964 => 24489,
    23965 => 24487,
    23966 => 24484,
    23967 => 24482,
    23968 => 24480,
    23969 => 24478,
    23970 => 24476,
    23971 => 24474,
    23972 => 24472,
    23973 => 24470,
    23974 => 24468,
    23975 => 24466,
    23976 => 24464,
    23977 => 24461,
    23978 => 24459,
    23979 => 24457,
    23980 => 24455,
    23981 => 24453,
    23982 => 24451,
    23983 => 24449,
    23984 => 24447,
    23985 => 24445,
    23986 => 24443,
    23987 => 24441,
    23988 => 24438,
    23989 => 24436,
    23990 => 24434,
    23991 => 24432,
    23992 => 24430,
    23993 => 24428,
    23994 => 24426,
    23995 => 24424,
    23996 => 24422,
    23997 => 24420,
    23998 => 24417,
    23999 => 24415,
    24000 => 24413,
    24001 => 24411,
    24002 => 24409,
    24003 => 24407,
    24004 => 24405,
    24005 => 24403,
    24006 => 24401,
    24007 => 24399,
    24008 => 24397,
    24009 => 24394,
    24010 => 24392,
    24011 => 24390,
    24012 => 24388,
    24013 => 24386,
    24014 => 24384,
    24015 => 24382,
    24016 => 24380,
    24017 => 24378,
    24018 => 24376,
    24019 => 24373,
    24020 => 24371,
    24021 => 24369,
    24022 => 24367,
    24023 => 24365,
    24024 => 24363,
    24025 => 24361,
    24026 => 24359,
    24027 => 24357,
    24028 => 24355,
    24029 => 24352,
    24030 => 24350,
    24031 => 24348,
    24032 => 24346,
    24033 => 24344,
    24034 => 24342,
    24035 => 24340,
    24036 => 24338,
    24037 => 24336,
    24038 => 24334,
    24039 => 24331,
    24040 => 24329,
    24041 => 24327,
    24042 => 24325,
    24043 => 24323,
    24044 => 24321,
    24045 => 24319,
    24046 => 24317,
    24047 => 24315,
    24048 => 24312,
    24049 => 24310,
    24050 => 24308,
    24051 => 24306,
    24052 => 24304,
    24053 => 24302,
    24054 => 24300,
    24055 => 24298,
    24056 => 24296,
    24057 => 24294,
    24058 => 24291,
    24059 => 24289,
    24060 => 24287,
    24061 => 24285,
    24062 => 24283,
    24063 => 24281,
    24064 => 24279,
    24065 => 24277,
    24066 => 24275,
    24067 => 24272,
    24068 => 24270,
    24069 => 24268,
    24070 => 24266,
    24071 => 24264,
    24072 => 24262,
    24073 => 24260,
    24074 => 24258,
    24075 => 24256,
    24076 => 24253,
    24077 => 24251,
    24078 => 24249,
    24079 => 24247,
    24080 => 24245,
    24081 => 24243,
    24082 => 24241,
    24083 => 24239,
    24084 => 24237,
    24085 => 24234,
    24086 => 24232,
    24087 => 24230,
    24088 => 24228,
    24089 => 24226,
    24090 => 24224,
    24091 => 24222,
    24092 => 24220,
    24093 => 24217,
    24094 => 24215,
    24095 => 24213,
    24096 => 24211,
    24097 => 24209,
    24098 => 24207,
    24099 => 24205,
    24100 => 24203,
    24101 => 24201,
    24102 => 24198,
    24103 => 24196,
    24104 => 24194,
    24105 => 24192,
    24106 => 24190,
    24107 => 24188,
    24108 => 24186,
    24109 => 24184,
    24110 => 24181,
    24111 => 24179,
    24112 => 24177,
    24113 => 24175,
    24114 => 24173,
    24115 => 24171,
    24116 => 24169,
    24117 => 24167,
    24118 => 24164,
    24119 => 24162,
    24120 => 24160,
    24121 => 24158,
    24122 => 24156,
    24123 => 24154,
    24124 => 24152,
    24125 => 24150,
    24126 => 24148,
    24127 => 24145,
    24128 => 24143,
    24129 => 24141,
    24130 => 24139,
    24131 => 24137,
    24132 => 24135,
    24133 => 24133,
    24134 => 24131,
    24135 => 24128,
    24136 => 24126,
    24137 => 24124,
    24138 => 24122,
    24139 => 24120,
    24140 => 24118,
    24141 => 24116,
    24142 => 24114,
    24143 => 24111,
    24144 => 24109,
    24145 => 24107,
    24146 => 24105,
    24147 => 24103,
    24148 => 24101,
    24149 => 24099,
    24150 => 24096,
    24151 => 24094,
    24152 => 24092,
    24153 => 24090,
    24154 => 24088,
    24155 => 24086,
    24156 => 24084,
    24157 => 24082,
    24158 => 24079,
    24159 => 24077,
    24160 => 24075,
    24161 => 24073,
    24162 => 24071,
    24163 => 24069,
    24164 => 24067,
    24165 => 24065,
    24166 => 24062,
    24167 => 24060,
    24168 => 24058,
    24169 => 24056,
    24170 => 24054,
    24171 => 24052,
    24172 => 24050,
    24173 => 24047,
    24174 => 24045,
    24175 => 24043,
    24176 => 24041,
    24177 => 24039,
    24178 => 24037,
    24179 => 24035,
    24180 => 24033,
    24181 => 24030,
    24182 => 24028,
    24183 => 24026,
    24184 => 24024,
    24185 => 24022,
    24186 => 24020,
    24187 => 24018,
    24188 => 24015,
    24189 => 24013,
    24190 => 24011,
    24191 => 24009,
    24192 => 24007,
    24193 => 24005,
    24194 => 24003,
    24195 => 24000,
    24196 => 23998,
    24197 => 23996,
    24198 => 23994,
    24199 => 23992,
    24200 => 23990,
    24201 => 23988,
    24202 => 23985,
    24203 => 23983,
    24204 => 23981,
    24205 => 23979,
    24206 => 23977,
    24207 => 23975,
    24208 => 23973,
    24209 => 23971,
    24210 => 23968,
    24211 => 23966,
    24212 => 23964,
    24213 => 23962,
    24214 => 23960,
    24215 => 23958,
    24216 => 23956,
    24217 => 23953,
    24218 => 23951,
    24219 => 23949,
    24220 => 23947,
    24221 => 23945,
    24222 => 23943,
    24223 => 23940,
    24224 => 23938,
    24225 => 23936,
    24226 => 23934,
    24227 => 23932,
    24228 => 23930,
    24229 => 23928,
    24230 => 23925,
    24231 => 23923,
    24232 => 23921,
    24233 => 23919,
    24234 => 23917,
    24235 => 23915,
    24236 => 23913,
    24237 => 23910,
    24238 => 23908,
    24239 => 23906,
    24240 => 23904,
    24241 => 23902,
    24242 => 23900,
    24243 => 23898,
    24244 => 23895,
    24245 => 23893,
    24246 => 23891,
    24247 => 23889,
    24248 => 23887,
    24249 => 23885,
    24250 => 23883,
    24251 => 23880,
    24252 => 23878,
    24253 => 23876,
    24254 => 23874,
    24255 => 23872,
    24256 => 23870,
    24257 => 23867,
    24258 => 23865,
    24259 => 23863,
    24260 => 23861,
    24261 => 23859,
    24262 => 23857,
    24263 => 23855,
    24264 => 23852,
    24265 => 23850,
    24266 => 23848,
    24267 => 23846,
    24268 => 23844,
    24269 => 23842,
    24270 => 23839,
    24271 => 23837,
    24272 => 23835,
    24273 => 23833,
    24274 => 23831,
    24275 => 23829,
    24276 => 23827,
    24277 => 23824,
    24278 => 23822,
    24279 => 23820,
    24280 => 23818,
    24281 => 23816,
    24282 => 23814,
    24283 => 23811,
    24284 => 23809,
    24285 => 23807,
    24286 => 23805,
    24287 => 23803,
    24288 => 23801,
    24289 => 23798,
    24290 => 23796,
    24291 => 23794,
    24292 => 23792,
    24293 => 23790,
    24294 => 23788,
    24295 => 23785,
    24296 => 23783,
    24297 => 23781,
    24298 => 23779,
    24299 => 23777,
    24300 => 23775,
    24301 => 23773,
    24302 => 23770,
    24303 => 23768,
    24304 => 23766,
    24305 => 23764,
    24306 => 23762,
    24307 => 23760,
    24308 => 23757,
    24309 => 23755,
    24310 => 23753,
    24311 => 23751,
    24312 => 23749,
    24313 => 23747,
    24314 => 23744,
    24315 => 23742,
    24316 => 23740,
    24317 => 23738,
    24318 => 23736,
    24319 => 23734,
    24320 => 23731,
    24321 => 23729,
    24322 => 23727,
    24323 => 23725,
    24324 => 23723,
    24325 => 23721,
    24326 => 23718,
    24327 => 23716,
    24328 => 23714,
    24329 => 23712,
    24330 => 23710,
    24331 => 23708,
    24332 => 23705,
    24333 => 23703,
    24334 => 23701,
    24335 => 23699,
    24336 => 23697,
    24337 => 23695,
    24338 => 23692,
    24339 => 23690,
    24340 => 23688,
    24341 => 23686,
    24342 => 23684,
    24343 => 23682,
    24344 => 23679,
    24345 => 23677,
    24346 => 23675,
    24347 => 23673,
    24348 => 23671,
    24349 => 23668,
    24350 => 23666,
    24351 => 23664,
    24352 => 23662,
    24353 => 23660,
    24354 => 23658,
    24355 => 23655,
    24356 => 23653,
    24357 => 23651,
    24358 => 23649,
    24359 => 23647,
    24360 => 23645,
    24361 => 23642,
    24362 => 23640,
    24363 => 23638,
    24364 => 23636,
    24365 => 23634,
    24366 => 23632,
    24367 => 23629,
    24368 => 23627,
    24369 => 23625,
    24370 => 23623,
    24371 => 23621,
    24372 => 23618,
    24373 => 23616,
    24374 => 23614,
    24375 => 23612,
    24376 => 23610,
    24377 => 23608,
    24378 => 23605,
    24379 => 23603,
    24380 => 23601,
    24381 => 23599,
    24382 => 23597,
    24383 => 23595,
    24384 => 23592,
    24385 => 23590,
    24386 => 23588,
    24387 => 23586,
    24388 => 23584,
    24389 => 23581,
    24390 => 23579,
    24391 => 23577,
    24392 => 23575,
    24393 => 23573,
    24394 => 23571,
    24395 => 23568,
    24396 => 23566,
    24397 => 23564,
    24398 => 23562,
    24399 => 23560,
    24400 => 23557,
    24401 => 23555,
    24402 => 23553,
    24403 => 23551,
    24404 => 23549,
    24405 => 23546,
    24406 => 23544,
    24407 => 23542,
    24408 => 23540,
    24409 => 23538,
    24410 => 23536,
    24411 => 23533,
    24412 => 23531,
    24413 => 23529,
    24414 => 23527,
    24415 => 23525,
    24416 => 23522,
    24417 => 23520,
    24418 => 23518,
    24419 => 23516,
    24420 => 23514,
    24421 => 23512,
    24422 => 23509,
    24423 => 23507,
    24424 => 23505,
    24425 => 23503,
    24426 => 23501,
    24427 => 23498,
    24428 => 23496,
    24429 => 23494,
    24430 => 23492,
    24431 => 23490,
    24432 => 23487,
    24433 => 23485,
    24434 => 23483,
    24435 => 23481,
    24436 => 23479,
    24437 => 23476,
    24438 => 23474,
    24439 => 23472,
    24440 => 23470,
    24441 => 23468,
    24442 => 23466,
    24443 => 23463,
    24444 => 23461,
    24445 => 23459,
    24446 => 23457,
    24447 => 23455,
    24448 => 23452,
    24449 => 23450,
    24450 => 23448,
    24451 => 23446,
    24452 => 23444,
    24453 => 23441,
    24454 => 23439,
    24455 => 23437,
    24456 => 23435,
    24457 => 23433,
    24458 => 23430,
    24459 => 23428,
    24460 => 23426,
    24461 => 23424,
    24462 => 23422,
    24463 => 23419,
    24464 => 23417,
    24465 => 23415,
    24466 => 23413,
    24467 => 23411,
    24468 => 23408,
    24469 => 23406,
    24470 => 23404,
    24471 => 23402,
    24472 => 23400,
    24473 => 23397,
    24474 => 23395,
    24475 => 23393,
    24476 => 23391,
    24477 => 23389,
    24478 => 23386,
    24479 => 23384,
    24480 => 23382,
    24481 => 23380,
    24482 => 23378,
    24483 => 23375,
    24484 => 23373,
    24485 => 23371,
    24486 => 23369,
    24487 => 23367,
    24488 => 23364,
    24489 => 23362,
    24490 => 23360,
    24491 => 23358,
    24492 => 23356,
    24493 => 23353,
    24494 => 23351,
    24495 => 23349,
    24496 => 23347,
    24497 => 23345,
    24498 => 23342,
    24499 => 23340,
    24500 => 23338,
    24501 => 23336,
    24502 => 23334,
    24503 => 23331,
    24504 => 23329,
    24505 => 23327,
    24506 => 23325,
    24507 => 23323,
    24508 => 23320,
    24509 => 23318,
    24510 => 23316,
    24511 => 23314,
    24512 => 23311,
    24513 => 23309,
    24514 => 23307,
    24515 => 23305,
    24516 => 23303,
    24517 => 23300,
    24518 => 23298,
    24519 => 23296,
    24520 => 23294,
    24521 => 23292,
    24522 => 23289,
    24523 => 23287,
    24524 => 23285,
    24525 => 23283,
    24526 => 23281,
    24527 => 23278,
    24528 => 23276,
    24529 => 23274,
    24530 => 23272,
    24531 => 23270,
    24532 => 23267,
    24533 => 23265,
    24534 => 23263,
    24535 => 23261,
    24536 => 23258,
    24537 => 23256,
    24538 => 23254,
    24539 => 23252,
    24540 => 23250,
    24541 => 23247,
    24542 => 23245,
    24543 => 23243,
    24544 => 23241,
    24545 => 23239,
    24546 => 23236,
    24547 => 23234,
    24548 => 23232,
    24549 => 23230,
    24550 => 23227,
    24551 => 23225,
    24552 => 23223,
    24553 => 23221,
    24554 => 23219,
    24555 => 23216,
    24556 => 23214,
    24557 => 23212,
    24558 => 23210,
    24559 => 23208,
    24560 => 23205,
    24561 => 23203,
    24562 => 23201,
    24563 => 23199,
    24564 => 23196,
    24565 => 23194,
    24566 => 23192,
    24567 => 23190,
    24568 => 23188,
    24569 => 23185,
    24570 => 23183,
    24571 => 23181,
    24572 => 23179,
    24573 => 23176,
    24574 => 23174,
    24575 => 23172,
    24576 => 23170,
    24577 => 23168,
    24578 => 23165,
    24579 => 23163,
    24580 => 23161,
    24581 => 23159,
    24582 => 23156,
    24583 => 23154,
    24584 => 23152,
    24585 => 23150,
    24586 => 23148,
    24587 => 23145,
    24588 => 23143,
    24589 => 23141,
    24590 => 23139,
    24591 => 23136,
    24592 => 23134,
    24593 => 23132,
    24594 => 23130,
    24595 => 23128,
    24596 => 23125,
    24597 => 23123,
    24598 => 23121,
    24599 => 23119,
    24600 => 23116,
    24601 => 23114,
    24602 => 23112,
    24603 => 23110,
    24604 => 23107,
    24605 => 23105,
    24606 => 23103,
    24607 => 23101,
    24608 => 23099,
    24609 => 23096,
    24610 => 23094,
    24611 => 23092,
    24612 => 23090,
    24613 => 23087,
    24614 => 23085,
    24615 => 23083,
    24616 => 23081,
    24617 => 23079,
    24618 => 23076,
    24619 => 23074,
    24620 => 23072,
    24621 => 23070,
    24622 => 23067,
    24623 => 23065,
    24624 => 23063,
    24625 => 23061,
    24626 => 23058,
    24627 => 23056,
    24628 => 23054,
    24629 => 23052,
    24630 => 23050,
    24631 => 23047,
    24632 => 23045,
    24633 => 23043,
    24634 => 23041,
    24635 => 23038,
    24636 => 23036,
    24637 => 23034,
    24638 => 23032,
    24639 => 23029,
    24640 => 23027,
    24641 => 23025,
    24642 => 23023,
    24643 => 23020,
    24644 => 23018,
    24645 => 23016,
    24646 => 23014,
    24647 => 23012,
    24648 => 23009,
    24649 => 23007,
    24650 => 23005,
    24651 => 23003,
    24652 => 23000,
    24653 => 22998,
    24654 => 22996,
    24655 => 22994,
    24656 => 22991,
    24657 => 22989,
    24658 => 22987,
    24659 => 22985,
    24660 => 22982,
    24661 => 22980,
    24662 => 22978,
    24663 => 22976,
    24664 => 22973,
    24665 => 22971,
    24666 => 22969,
    24667 => 22967,
    24668 => 22965,
    24669 => 22962,
    24670 => 22960,
    24671 => 22958,
    24672 => 22956,
    24673 => 22953,
    24674 => 22951,
    24675 => 22949,
    24676 => 22947,
    24677 => 22944,
    24678 => 22942,
    24679 => 22940,
    24680 => 22938,
    24681 => 22935,
    24682 => 22933,
    24683 => 22931,
    24684 => 22929,
    24685 => 22926,
    24686 => 22924,
    24687 => 22922,
    24688 => 22920,
    24689 => 22917,
    24690 => 22915,
    24691 => 22913,
    24692 => 22911,
    24693 => 22908,
    24694 => 22906,
    24695 => 22904,
    24696 => 22902,
    24697 => 22899,
    24698 => 22897,
    24699 => 22895,
    24700 => 22893,
    24701 => 22890,
    24702 => 22888,
    24703 => 22886,
    24704 => 22884,
    24705 => 22881,
    24706 => 22879,
    24707 => 22877,
    24708 => 22875,
    24709 => 22872,
    24710 => 22870,
    24711 => 22868,
    24712 => 22866,
    24713 => 22863,
    24714 => 22861,
    24715 => 22859,
    24716 => 22857,
    24717 => 22854,
    24718 => 22852,
    24719 => 22850,
    24720 => 22848,
    24721 => 22845,
    24722 => 22843,
    24723 => 22841,
    24724 => 22839,
    24725 => 22836,
    24726 => 22834,
    24727 => 22832,
    24728 => 22830,
    24729 => 22827,
    24730 => 22825,
    24731 => 22823,
    24732 => 22821,
    24733 => 22818,
    24734 => 22816,
    24735 => 22814,
    24736 => 22812,
    24737 => 22809,
    24738 => 22807,
    24739 => 22805,
    24740 => 22803,
    24741 => 22800,
    24742 => 22798,
    24743 => 22796,
    24744 => 22794,
    24745 => 22791,
    24746 => 22789,
    24747 => 22787,
    24748 => 22785,
    24749 => 22782,
    24750 => 22780,
    24751 => 22778,
    24752 => 22776,
    24753 => 22773,
    24754 => 22771,
    24755 => 22769,
    24756 => 22766,
    24757 => 22764,
    24758 => 22762,
    24759 => 22760,
    24760 => 22757,
    24761 => 22755,
    24762 => 22753,
    24763 => 22751,
    24764 => 22748,
    24765 => 22746,
    24766 => 22744,
    24767 => 22742,
    24768 => 22739,
    24769 => 22737,
    24770 => 22735,
    24771 => 22733,
    24772 => 22730,
    24773 => 22728,
    24774 => 22726,
    24775 => 22724,
    24776 => 22721,
    24777 => 22719,
    24778 => 22717,
    24779 => 22714,
    24780 => 22712,
    24781 => 22710,
    24782 => 22708,
    24783 => 22705,
    24784 => 22703,
    24785 => 22701,
    24786 => 22699,
    24787 => 22696,
    24788 => 22694,
    24789 => 22692,
    24790 => 22690,
    24791 => 22687,
    24792 => 22685,
    24793 => 22683,
    24794 => 22680,
    24795 => 22678,
    24796 => 22676,
    24797 => 22674,
    24798 => 22671,
    24799 => 22669,
    24800 => 22667,
    24801 => 22665,
    24802 => 22662,
    24803 => 22660,
    24804 => 22658,
    24805 => 22656,
    24806 => 22653,
    24807 => 22651,
    24808 => 22649,
    24809 => 22646,
    24810 => 22644,
    24811 => 22642,
    24812 => 22640,
    24813 => 22637,
    24814 => 22635,
    24815 => 22633,
    24816 => 22631,
    24817 => 22628,
    24818 => 22626,
    24819 => 22624,
    24820 => 22621,
    24821 => 22619,
    24822 => 22617,
    24823 => 22615,
    24824 => 22612,
    24825 => 22610,
    24826 => 22608,
    24827 => 22606,
    24828 => 22603,
    24829 => 22601,
    24830 => 22599,
    24831 => 22596,
    24832 => 22594,
    24833 => 22592,
    24834 => 22590,
    24835 => 22587,
    24836 => 22585,
    24837 => 22583,
    24838 => 22581,
    24839 => 22578,
    24840 => 22576,
    24841 => 22574,
    24842 => 22571,
    24843 => 22569,
    24844 => 22567,
    24845 => 22565,
    24846 => 22562,
    24847 => 22560,
    24848 => 22558,
    24849 => 22555,
    24850 => 22553,
    24851 => 22551,
    24852 => 22549,
    24853 => 22546,
    24854 => 22544,
    24855 => 22542,
    24856 => 22540,
    24857 => 22537,
    24858 => 22535,
    24859 => 22533,
    24860 => 22530,
    24861 => 22528,
    24862 => 22526,
    24863 => 22524,
    24864 => 22521,
    24865 => 22519,
    24866 => 22517,
    24867 => 22514,
    24868 => 22512,
    24869 => 22510,
    24870 => 22508,
    24871 => 22505,
    24872 => 22503,
    24873 => 22501,
    24874 => 22498,
    24875 => 22496,
    24876 => 22494,
    24877 => 22492,
    24878 => 22489,
    24879 => 22487,
    24880 => 22485,
    24881 => 22482,
    24882 => 22480,
    24883 => 22478,
    24884 => 22476,
    24885 => 22473,
    24886 => 22471,
    24887 => 22469,
    24888 => 22466,
    24889 => 22464,
    24890 => 22462,
    24891 => 22460,
    24892 => 22457,
    24893 => 22455,
    24894 => 22453,
    24895 => 22450,
    24896 => 22448,
    24897 => 22446,
    24898 => 22444,
    24899 => 22441,
    24900 => 22439,
    24901 => 22437,
    24902 => 22434,
    24903 => 22432,
    24904 => 22430,
    24905 => 22428,
    24906 => 22425,
    24907 => 22423,
    24908 => 22421,
    24909 => 22418,
    24910 => 22416,
    24911 => 22414,
    24912 => 22411,
    24913 => 22409,
    24914 => 22407,
    24915 => 22405,
    24916 => 22402,
    24917 => 22400,
    24918 => 22398,
    24919 => 22395,
    24920 => 22393,
    24921 => 22391,
    24922 => 22389,
    24923 => 22386,
    24924 => 22384,
    24925 => 22382,
    24926 => 22379,
    24927 => 22377,
    24928 => 22375,
    24929 => 22373,
    24930 => 22370,
    24931 => 22368,
    24932 => 22366,
    24933 => 22363,
    24934 => 22361,
    24935 => 22359,
    24936 => 22356,
    24937 => 22354,
    24938 => 22352,
    24939 => 22350,
    24940 => 22347,
    24941 => 22345,
    24942 => 22343,
    24943 => 22340,
    24944 => 22338,
    24945 => 22336,
    24946 => 22333,
    24947 => 22331,
    24948 => 22329,
    24949 => 22327,
    24950 => 22324,
    24951 => 22322,
    24952 => 22320,
    24953 => 22317,
    24954 => 22315,
    24955 => 22313,
    24956 => 22310,
    24957 => 22308,
    24958 => 22306,
    24959 => 22304,
    24960 => 22301,
    24961 => 22299,
    24962 => 22297,
    24963 => 22294,
    24964 => 22292,
    24965 => 22290,
    24966 => 22287,
    24967 => 22285,
    24968 => 22283,
    24969 => 22281,
    24970 => 22278,
    24971 => 22276,
    24972 => 22274,
    24973 => 22271,
    24974 => 22269,
    24975 => 22267,
    24976 => 22264,
    24977 => 22262,
    24978 => 22260,
    24979 => 22257,
    24980 => 22255,
    24981 => 22253,
    24982 => 22251,
    24983 => 22248,
    24984 => 22246,
    24985 => 22244,
    24986 => 22241,
    24987 => 22239,
    24988 => 22237,
    24989 => 22234,
    24990 => 22232,
    24991 => 22230,
    24992 => 22227,
    24993 => 22225,
    24994 => 22223,
    24995 => 22221,
    24996 => 22218,
    24997 => 22216,
    24998 => 22214,
    24999 => 22211,
    25000 => 22209,
    25001 => 22207,
    25002 => 22204,
    25003 => 22202,
    25004 => 22200,
    25005 => 22197,
    25006 => 22195,
    25007 => 22193,
    25008 => 22191,
    25009 => 22188,
    25010 => 22186,
    25011 => 22184,
    25012 => 22181,
    25013 => 22179,
    25014 => 22177,
    25015 => 22174,
    25016 => 22172,
    25017 => 22170,
    25018 => 22167,
    25019 => 22165,
    25020 => 22163,
    25021 => 22160,
    25022 => 22158,
    25023 => 22156,
    25024 => 22154,
    25025 => 22151,
    25026 => 22149,
    25027 => 22147,
    25028 => 22144,
    25029 => 22142,
    25030 => 22140,
    25031 => 22137,
    25032 => 22135,
    25033 => 22133,
    25034 => 22130,
    25035 => 22128,
    25036 => 22126,
    25037 => 22123,
    25038 => 22121,
    25039 => 22119,
    25040 => 22116,
    25041 => 22114,
    25042 => 22112,
    25043 => 22110,
    25044 => 22107,
    25045 => 22105,
    25046 => 22103,
    25047 => 22100,
    25048 => 22098,
    25049 => 22096,
    25050 => 22093,
    25051 => 22091,
    25052 => 22089,
    25053 => 22086,
    25054 => 22084,
    25055 => 22082,
    25056 => 22079,
    25057 => 22077,
    25058 => 22075,
    25059 => 22072,
    25060 => 22070,
    25061 => 22068,
    25062 => 22065,
    25063 => 22063,
    25064 => 22061,
    25065 => 22058,
    25066 => 22056,
    25067 => 22054,
    25068 => 22051,
    25069 => 22049,
    25070 => 22047,
    25071 => 22045,
    25072 => 22042,
    25073 => 22040,
    25074 => 22038,
    25075 => 22035,
    25076 => 22033,
    25077 => 22031,
    25078 => 22028,
    25079 => 22026,
    25080 => 22024,
    25081 => 22021,
    25082 => 22019,
    25083 => 22017,
    25084 => 22014,
    25085 => 22012,
    25086 => 22010,
    25087 => 22007,
    25088 => 22005,
    25089 => 22003,
    25090 => 22000,
    25091 => 21998,
    25092 => 21996,
    25093 => 21993,
    25094 => 21991,
    25095 => 21989,
    25096 => 21986,
    25097 => 21984,
    25098 => 21982,
    25099 => 21979,
    25100 => 21977,
    25101 => 21975,
    25102 => 21972,
    25103 => 21970,
    25104 => 21968,
    25105 => 21965,
    25106 => 21963,
    25107 => 21961,
    25108 => 21958,
    25109 => 21956,
    25110 => 21954,
    25111 => 21951,
    25112 => 21949,
    25113 => 21947,
    25114 => 21944,
    25115 => 21942,
    25116 => 21940,
    25117 => 21937,
    25118 => 21935,
    25119 => 21933,
    25120 => 21930,
    25121 => 21928,
    25122 => 21926,
    25123 => 21923,
    25124 => 21921,
    25125 => 21919,
    25126 => 21916,
    25127 => 21914,
    25128 => 21912,
    25129 => 21909,
    25130 => 21907,
    25131 => 21905,
    25132 => 21902,
    25133 => 21900,
    25134 => 21898,
    25135 => 21895,
    25136 => 21893,
    25137 => 21891,
    25138 => 21888,
    25139 => 21886,
    25140 => 21884,
    25141 => 21881,
    25142 => 21879,
    25143 => 21877,
    25144 => 21874,
    25145 => 21872,
    25146 => 21870,
    25147 => 21867,
    25148 => 21865,
    25149 => 21863,
    25150 => 21860,
    25151 => 21858,
    25152 => 21856,
    25153 => 21853,
    25154 => 21851,
    25155 => 21849,
    25156 => 21846,
    25157 => 21844,
    25158 => 21842,
    25159 => 21839,
    25160 => 21837,
    25161 => 21835,
    25162 => 21832,
    25163 => 21830,
    25164 => 21827,
    25165 => 21825,
    25166 => 21823,
    25167 => 21820,
    25168 => 21818,
    25169 => 21816,
    25170 => 21813,
    25171 => 21811,
    25172 => 21809,
    25173 => 21806,
    25174 => 21804,
    25175 => 21802,
    25176 => 21799,
    25177 => 21797,
    25178 => 21795,
    25179 => 21792,
    25180 => 21790,
    25181 => 21788,
    25182 => 21785,
    25183 => 21783,
    25184 => 21781,
    25185 => 21778,
    25186 => 21776,
    25187 => 21774,
    25188 => 21771,
    25189 => 21769,
    25190 => 21766,
    25191 => 21764,
    25192 => 21762,
    25193 => 21759,
    25194 => 21757,
    25195 => 21755,
    25196 => 21752,
    25197 => 21750,
    25198 => 21748,
    25199 => 21745,
    25200 => 21743,
    25201 => 21741,
    25202 => 21738,
    25203 => 21736,
    25204 => 21734,
    25205 => 21731,
    25206 => 21729,
    25207 => 21727,
    25208 => 21724,
    25209 => 21722,
    25210 => 21719,
    25211 => 21717,
    25212 => 21715,
    25213 => 21712,
    25214 => 21710,
    25215 => 21708,
    25216 => 21705,
    25217 => 21703,
    25218 => 21701,
    25219 => 21698,
    25220 => 21696,
    25221 => 21694,
    25222 => 21691,
    25223 => 21689,
    25224 => 21687,
    25225 => 21684,
    25226 => 21682,
    25227 => 21679,
    25228 => 21677,
    25229 => 21675,
    25230 => 21672,
    25231 => 21670,
    25232 => 21668,
    25233 => 21665,
    25234 => 21663,
    25235 => 21661,
    25236 => 21658,
    25237 => 21656,
    25238 => 21654,
    25239 => 21651,
    25240 => 21649,
    25241 => 21646,
    25242 => 21644,
    25243 => 21642,
    25244 => 21639,
    25245 => 21637,
    25246 => 21635,
    25247 => 21632,
    25248 => 21630,
    25249 => 21628,
    25250 => 21625,
    25251 => 21623,
    25252 => 21621,
    25253 => 21618,
    25254 => 21616,
    25255 => 21613,
    25256 => 21611,
    25257 => 21609,
    25258 => 21606,
    25259 => 21604,
    25260 => 21602,
    25261 => 21599,
    25262 => 21597,
    25263 => 21595,
    25264 => 21592,
    25265 => 21590,
    25266 => 21587,
    25267 => 21585,
    25268 => 21583,
    25269 => 21580,
    25270 => 21578,
    25271 => 21576,
    25272 => 21573,
    25273 => 21571,
    25274 => 21569,
    25275 => 21566,
    25276 => 21564,
    25277 => 21561,
    25278 => 21559,
    25279 => 21557,
    25280 => 21554,
    25281 => 21552,
    25282 => 21550,
    25283 => 21547,
    25284 => 21545,
    25285 => 21543,
    25286 => 21540,
    25287 => 21538,
    25288 => 21535,
    25289 => 21533,
    25290 => 21531,
    25291 => 21528,
    25292 => 21526,
    25293 => 21524,
    25294 => 21521,
    25295 => 21519,
    25296 => 21516,
    25297 => 21514,
    25298 => 21512,
    25299 => 21509,
    25300 => 21507,
    25301 => 21505,
    25302 => 21502,
    25303 => 21500,
    25304 => 21498,
    25305 => 21495,
    25306 => 21493,
    25307 => 21490,
    25308 => 21488,
    25309 => 21486,
    25310 => 21483,
    25311 => 21481,
    25312 => 21479,
    25313 => 21476,
    25314 => 21474,
    25315 => 21471,
    25316 => 21469,
    25317 => 21467,
    25318 => 21464,
    25319 => 21462,
    25320 => 21460,
    25321 => 21457,
    25322 => 21455,
    25323 => 21452,
    25324 => 21450,
    25325 => 21448,
    25326 => 21445,
    25327 => 21443,
    25328 => 21441,
    25329 => 21438,
    25330 => 21436,
    25331 => 21433,
    25332 => 21431,
    25333 => 21429,
    25334 => 21426,
    25335 => 21424,
    25336 => 21422,
    25337 => 21419,
    25338 => 21417,
    25339 => 21414,
    25340 => 21412,
    25341 => 21410,
    25342 => 21407,
    25343 => 21405,
    25344 => 21403,
    25345 => 21400,
    25346 => 21398,
    25347 => 21395,
    25348 => 21393,
    25349 => 21391,
    25350 => 21388,
    25351 => 21386,
    25352 => 21383,
    25353 => 21381,
    25354 => 21379,
    25355 => 21376,
    25356 => 21374,
    25357 => 21372,
    25358 => 21369,
    25359 => 21367,
    25360 => 21364,
    25361 => 21362,
    25362 => 21360,
    25363 => 21357,
    25364 => 21355,
    25365 => 21353,
    25366 => 21350,
    25367 => 21348,
    25368 => 21345,
    25369 => 21343,
    25370 => 21341,
    25371 => 21338,
    25372 => 21336,
    25373 => 21333,
    25374 => 21331,
    25375 => 21329,
    25376 => 21326,
    25377 => 21324,
    25378 => 21322,
    25379 => 21319,
    25380 => 21317,
    25381 => 21314,
    25382 => 21312,
    25383 => 21310,
    25384 => 21307,
    25385 => 21305,
    25386 => 21302,
    25387 => 21300,
    25388 => 21298,
    25389 => 21295,
    25390 => 21293,
    25391 => 21290,
    25392 => 21288,
    25393 => 21286,
    25394 => 21283,
    25395 => 21281,
    25396 => 21279,
    25397 => 21276,
    25398 => 21274,
    25399 => 21271,
    25400 => 21269,
    25401 => 21267,
    25402 => 21264,
    25403 => 21262,
    25404 => 21259,
    25405 => 21257,
    25406 => 21255,
    25407 => 21252,
    25408 => 21250,
    25409 => 21247,
    25410 => 21245,
    25411 => 21243,
    25412 => 21240,
    25413 => 21238,
    25414 => 21236,
    25415 => 21233,
    25416 => 21231,
    25417 => 21228,
    25418 => 21226,
    25419 => 21224,
    25420 => 21221,
    25421 => 21219,
    25422 => 21216,
    25423 => 21214,
    25424 => 21212,
    25425 => 21209,
    25426 => 21207,
    25427 => 21204,
    25428 => 21202,
    25429 => 21200,
    25430 => 21197,
    25431 => 21195,
    25432 => 21192,
    25433 => 21190,
    25434 => 21188,
    25435 => 21185,
    25436 => 21183,
    25437 => 21180,
    25438 => 21178,
    25439 => 21176,
    25440 => 21173,
    25441 => 21171,
    25442 => 21168,
    25443 => 21166,
    25444 => 21164,
    25445 => 21161,
    25446 => 21159,
    25447 => 21156,
    25448 => 21154,
    25449 => 21152,
    25450 => 21149,
    25451 => 21147,
    25452 => 21144,
    25453 => 21142,
    25454 => 21140,
    25455 => 21137,
    25456 => 21135,
    25457 => 21132,
    25458 => 21130,
    25459 => 21128,
    25460 => 21125,
    25461 => 21123,
    25462 => 21120,
    25463 => 21118,
    25464 => 21116,
    25465 => 21113,
    25466 => 21111,
    25467 => 21108,
    25468 => 21106,
    25469 => 21104,
    25470 => 21101,
    25471 => 21099,
    25472 => 21096,
    25473 => 21094,
    25474 => 21092,
    25475 => 21089,
    25476 => 21087,
    25477 => 21084,
    25478 => 21082,
    25479 => 21080,
    25480 => 21077,
    25481 => 21075,
    25482 => 21072,
    25483 => 21070,
    25484 => 21068,
    25485 => 21065,
    25486 => 21063,
    25487 => 21060,
    25488 => 21058,
    25489 => 21056,
    25490 => 21053,
    25491 => 21051,
    25492 => 21048,
    25493 => 21046,
    25494 => 21043,
    25495 => 21041,
    25496 => 21039,
    25497 => 21036,
    25498 => 21034,
    25499 => 21031,
    25500 => 21029,
    25501 => 21027,
    25502 => 21024,
    25503 => 21022,
    25504 => 21019,
    25505 => 21017,
    25506 => 21015,
    25507 => 21012,
    25508 => 21010,
    25509 => 21007,
    25510 => 21005,
    25511 => 21003,
    25512 => 21000,
    25513 => 20998,
    25514 => 20995,
    25515 => 20993,
    25516 => 20990,
    25517 => 20988,
    25518 => 20986,
    25519 => 20983,
    25520 => 20981,
    25521 => 20978,
    25522 => 20976,
    25523 => 20974,
    25524 => 20971,
    25525 => 20969,
    25526 => 20966,
    25527 => 20964,
    25528 => 20962,
    25529 => 20959,
    25530 => 20957,
    25531 => 20954,
    25532 => 20952,
    25533 => 20949,
    25534 => 20947,
    25535 => 20945,
    25536 => 20942,
    25537 => 20940,
    25538 => 20937,
    25539 => 20935,
    25540 => 20933,
    25541 => 20930,
    25542 => 20928,
    25543 => 20925,
    25544 => 20923,
    25545 => 20920,
    25546 => 20918,
    25547 => 20916,
    25548 => 20913,
    25549 => 20911,
    25550 => 20908,
    25551 => 20906,
    25552 => 20904,
    25553 => 20901,
    25554 => 20899,
    25555 => 20896,
    25556 => 20894,
    25557 => 20891,
    25558 => 20889,
    25559 => 20887,
    25560 => 20884,
    25561 => 20882,
    25562 => 20879,
    25563 => 20877,
    25564 => 20874,
    25565 => 20872,
    25566 => 20870,
    25567 => 20867,
    25568 => 20865,
    25569 => 20862,
    25570 => 20860,
    25571 => 20858,
    25572 => 20855,
    25573 => 20853,
    25574 => 20850,
    25575 => 20848,
    25576 => 20845,
    25577 => 20843,
    25578 => 20841,
    25579 => 20838,
    25580 => 20836,
    25581 => 20833,
    25582 => 20831,
    25583 => 20828,
    25584 => 20826,
    25585 => 20824,
    25586 => 20821,
    25587 => 20819,
    25588 => 20816,
    25589 => 20814,
    25590 => 20811,
    25591 => 20809,
    25592 => 20807,
    25593 => 20804,
    25594 => 20802,
    25595 => 20799,
    25596 => 20797,
    25597 => 20794,
    25598 => 20792,
    25599 => 20790,
    25600 => 20787,
    25601 => 20785,
    25602 => 20782,
    25603 => 20780,
    25604 => 20777,
    25605 => 20775,
    25606 => 20773,
    25607 => 20770,
    25608 => 20768,
    25609 => 20765,
    25610 => 20763,
    25611 => 20760,
    25612 => 20758,
    25613 => 20756,
    25614 => 20753,
    25615 => 20751,
    25616 => 20748,
    25617 => 20746,
    25618 => 20743,
    25619 => 20741,
    25620 => 20739,
    25621 => 20736,
    25622 => 20734,
    25623 => 20731,
    25624 => 20729,
    25625 => 20726,
    25626 => 20724,
    25627 => 20722,
    25628 => 20719,
    25629 => 20717,
    25630 => 20714,
    25631 => 20712,
    25632 => 20709,
    25633 => 20707,
    25634 => 20704,
    25635 => 20702,
    25636 => 20700,
    25637 => 20697,
    25638 => 20695,
    25639 => 20692,
    25640 => 20690,
    25641 => 20687,
    25642 => 20685,
    25643 => 20683,
    25644 => 20680,
    25645 => 20678,
    25646 => 20675,
    25647 => 20673,
    25648 => 20670,
    25649 => 20668,
    25650 => 20666,
    25651 => 20663,
    25652 => 20661,
    25653 => 20658,
    25654 => 20656,
    25655 => 20653,
    25656 => 20651,
    25657 => 20648,
    25658 => 20646,
    25659 => 20644,
    25660 => 20641,
    25661 => 20639,
    25662 => 20636,
    25663 => 20634,
    25664 => 20631,
    25665 => 20629,
    25666 => 20626,
    25667 => 20624,
    25668 => 20622,
    25669 => 20619,
    25670 => 20617,
    25671 => 20614,
    25672 => 20612,
    25673 => 20609,
    25674 => 20607,
    25675 => 20604,
    25676 => 20602,
    25677 => 20600,
    25678 => 20597,
    25679 => 20595,
    25680 => 20592,
    25681 => 20590,
    25682 => 20587,
    25683 => 20585,
    25684 => 20583,
    25685 => 20580,
    25686 => 20578,
    25687 => 20575,
    25688 => 20573,
    25689 => 20570,
    25690 => 20568,
    25691 => 20565,
    25692 => 20563,
    25693 => 20560,
    25694 => 20558,
    25695 => 20556,
    25696 => 20553,
    25697 => 20551,
    25698 => 20548,
    25699 => 20546,
    25700 => 20543,
    25701 => 20541,
    25702 => 20538,
    25703 => 20536,
    25704 => 20534,
    25705 => 20531,
    25706 => 20529,
    25707 => 20526,
    25708 => 20524,
    25709 => 20521,
    25710 => 20519,
    25711 => 20516,
    25712 => 20514,
    25713 => 20512,
    25714 => 20509,
    25715 => 20507,
    25716 => 20504,
    25717 => 20502,
    25718 => 20499,
    25719 => 20497,
    25720 => 20494,
    25721 => 20492,
    25722 => 20489,
    25723 => 20487,
    25724 => 20485,
    25725 => 20482,
    25726 => 20480,
    25727 => 20477,
    25728 => 20475,
    25729 => 20472,
    25730 => 20470,
    25731 => 20467,
    25732 => 20465,
    25733 => 20463,
    25734 => 20460,
    25735 => 20458,
    25736 => 20455,
    25737 => 20453,
    25738 => 20450,
    25739 => 20448,
    25740 => 20445,
    25741 => 20443,
    25742 => 20440,
    25743 => 20438,
    25744 => 20436,
    25745 => 20433,
    25746 => 20431,
    25747 => 20428,
    25748 => 20426,
    25749 => 20423,
    25750 => 20421,
    25751 => 20418,
    25752 => 20416,
    25753 => 20413,
    25754 => 20411,
    25755 => 20408,
    25756 => 20406,
    25757 => 20404,
    25758 => 20401,
    25759 => 20399,
    25760 => 20396,
    25761 => 20394,
    25762 => 20391,
    25763 => 20389,
    25764 => 20386,
    25765 => 20384,
    25766 => 20381,
    25767 => 20379,
    25768 => 20377,
    25769 => 20374,
    25770 => 20372,
    25771 => 20369,
    25772 => 20367,
    25773 => 20364,
    25774 => 20362,
    25775 => 20359,
    25776 => 20357,
    25777 => 20354,
    25778 => 20352,
    25779 => 20349,
    25780 => 20347,
    25781 => 20345,
    25782 => 20342,
    25783 => 20340,
    25784 => 20337,
    25785 => 20335,
    25786 => 20332,
    25787 => 20330,
    25788 => 20327,
    25789 => 20325,
    25790 => 20322,
    25791 => 20320,
    25792 => 20317,
    25793 => 20315,
    25794 => 20312,
    25795 => 20310,
    25796 => 20308,
    25797 => 20305,
    25798 => 20303,
    25799 => 20300,
    25800 => 20298,
    25801 => 20295,
    25802 => 20293,
    25803 => 20290,
    25804 => 20288,
    25805 => 20285,
    25806 => 20283,
    25807 => 20280,
    25808 => 20278,
    25809 => 20275,
    25810 => 20273,
    25811 => 20271,
    25812 => 20268,
    25813 => 20266,
    25814 => 20263,
    25815 => 20261,
    25816 => 20258,
    25817 => 20256,
    25818 => 20253,
    25819 => 20251,
    25820 => 20248,
    25821 => 20246,
    25822 => 20243,
    25823 => 20241,
    25824 => 20238,
    25825 => 20236,
    25826 => 20234,
    25827 => 20231,
    25828 => 20229,
    25829 => 20226,
    25830 => 20224,
    25831 => 20221,
    25832 => 20219,
    25833 => 20216,
    25834 => 20214,
    25835 => 20211,
    25836 => 20209,
    25837 => 20206,
    25838 => 20204,
    25839 => 20201,
    25840 => 20199,
    25841 => 20196,
    25842 => 20194,
    25843 => 20191,
    25844 => 20189,
    25845 => 20187,
    25846 => 20184,
    25847 => 20182,
    25848 => 20179,
    25849 => 20177,
    25850 => 20174,
    25851 => 20172,
    25852 => 20169,
    25853 => 20167,
    25854 => 20164,
    25855 => 20162,
    25856 => 20159,
    25857 => 20157,
    25858 => 20154,
    25859 => 20152,
    25860 => 20149,
    25861 => 20147,
    25862 => 20144,
    25863 => 20142,
    25864 => 20139,
    25865 => 20137,
    25866 => 20135,
    25867 => 20132,
    25868 => 20130,
    25869 => 20127,
    25870 => 20125,
    25871 => 20122,
    25872 => 20120,
    25873 => 20117,
    25874 => 20115,
    25875 => 20112,
    25876 => 20110,
    25877 => 20107,
    25878 => 20105,
    25879 => 20102,
    25880 => 20100,
    25881 => 20097,
    25882 => 20095,
    25883 => 20092,
    25884 => 20090,
    25885 => 20087,
    25886 => 20085,
    25887 => 20082,
    25888 => 20080,
    25889 => 20077,
    25890 => 20075,
    25891 => 20072,
    25892 => 20070,
    25893 => 20068,
    25894 => 20065,
    25895 => 20063,
    25896 => 20060,
    25897 => 20058,
    25898 => 20055,
    25899 => 20053,
    25900 => 20050,
    25901 => 20048,
    25902 => 20045,
    25903 => 20043,
    25904 => 20040,
    25905 => 20038,
    25906 => 20035,
    25907 => 20033,
    25908 => 20030,
    25909 => 20028,
    25910 => 20025,
    25911 => 20023,
    25912 => 20020,
    25913 => 20018,
    25914 => 20015,
    25915 => 20013,
    25916 => 20010,
    25917 => 20008,
    25918 => 20005,
    25919 => 20003,
    25920 => 20000,
    25921 => 19998,
    25922 => 19995,
    25923 => 19993,
    25924 => 19990,
    25925 => 19988,
    25926 => 19985,
    25927 => 19983,
    25928 => 19981,
    25929 => 19978,
    25930 => 19976,
    25931 => 19973,
    25932 => 19971,
    25933 => 19968,
    25934 => 19966,
    25935 => 19963,
    25936 => 19961,
    25937 => 19958,
    25938 => 19956,
    25939 => 19953,
    25940 => 19951,
    25941 => 19948,
    25942 => 19946,
    25943 => 19943,
    25944 => 19941,
    25945 => 19938,
    25946 => 19936,
    25947 => 19933,
    25948 => 19931,
    25949 => 19928,
    25950 => 19926,
    25951 => 19923,
    25952 => 19921,
    25953 => 19918,
    25954 => 19916,
    25955 => 19913,
    25956 => 19911,
    25957 => 19908,
    25958 => 19906,
    25959 => 19903,
    25960 => 19901,
    25961 => 19898,
    25962 => 19896,
    25963 => 19893,
    25964 => 19891,
    25965 => 19888,
    25966 => 19886,
    25967 => 19883,
    25968 => 19881,
    25969 => 19878,
    25970 => 19876,
    25971 => 19873,
    25972 => 19871,
    25973 => 19868,
    25974 => 19866,
    25975 => 19863,
    25976 => 19861,
    25977 => 19858,
    25978 => 19856,
    25979 => 19853,
    25980 => 19851,
    25981 => 19848,
    25982 => 19846,
    25983 => 19843,
    25984 => 19841,
    25985 => 19838,
    25986 => 19836,
    25987 => 19833,
    25988 => 19831,
    25989 => 19828,
    25990 => 19826,
    25991 => 19823,
    25992 => 19821,
    25993 => 19818,
    25994 => 19816,
    25995 => 19813,
    25996 => 19811,
    25997 => 19808,
    25998 => 19806,
    25999 => 19803,
    26000 => 19801,
    26001 => 19798,
    26002 => 19796,
    26003 => 19793,
    26004 => 19791,
    26005 => 19788,
    26006 => 19786,
    26007 => 19783,
    26008 => 19781,
    26009 => 19778,
    26010 => 19776,
    26011 => 19773,
    26012 => 19771,
    26013 => 19768,
    26014 => 19766,
    26015 => 19763,
    26016 => 19761,
    26017 => 19758,
    26018 => 19756,
    26019 => 19753,
    26020 => 19751,
    26021 => 19748,
    26022 => 19746,
    26023 => 19743,
    26024 => 19741,
    26025 => 19738,
    26026 => 19736,
    26027 => 19733,
    26028 => 19731,
    26029 => 19728,
    26030 => 19726,
    26031 => 19723,
    26032 => 19721,
    26033 => 19718,
    26034 => 19716,
    26035 => 19713,
    26036 => 19711,
    26037 => 19708,
    26038 => 19706,
    26039 => 19703,
    26040 => 19700,
    26041 => 19698,
    26042 => 19695,
    26043 => 19693,
    26044 => 19690,
    26045 => 19688,
    26046 => 19685,
    26047 => 19683,
    26048 => 19680,
    26049 => 19678,
    26050 => 19675,
    26051 => 19673,
    26052 => 19670,
    26053 => 19668,
    26054 => 19665,
    26055 => 19663,
    26056 => 19660,
    26057 => 19658,
    26058 => 19655,
    26059 => 19653,
    26060 => 19650,
    26061 => 19648,
    26062 => 19645,
    26063 => 19643,
    26064 => 19640,
    26065 => 19638,
    26066 => 19635,
    26067 => 19633,
    26068 => 19630,
    26069 => 19628,
    26070 => 19625,
    26071 => 19623,
    26072 => 19620,
    26073 => 19618,
    26074 => 19615,
    26075 => 19613,
    26076 => 19610,
    26077 => 19607,
    26078 => 19605,
    26079 => 19602,
    26080 => 19600,
    26081 => 19597,
    26082 => 19595,
    26083 => 19592,
    26084 => 19590,
    26085 => 19587,
    26086 => 19585,
    26087 => 19582,
    26088 => 19580,
    26089 => 19577,
    26090 => 19575,
    26091 => 19572,
    26092 => 19570,
    26093 => 19567,
    26094 => 19565,
    26095 => 19562,
    26096 => 19560,
    26097 => 19557,
    26098 => 19555,
    26099 => 19552,
    26100 => 19550,
    26101 => 19547,
    26102 => 19545,
    26103 => 19542,
    26104 => 19539,
    26105 => 19537,
    26106 => 19534,
    26107 => 19532,
    26108 => 19529,
    26109 => 19527,
    26110 => 19524,
    26111 => 19522,
    26112 => 19519,
    26113 => 19517,
    26114 => 19514,
    26115 => 19512,
    26116 => 19509,
    26117 => 19507,
    26118 => 19504,
    26119 => 19502,
    26120 => 19499,
    26121 => 19497,
    26122 => 19494,
    26123 => 19492,
    26124 => 19489,
    26125 => 19486,
    26126 => 19484,
    26127 => 19481,
    26128 => 19479,
    26129 => 19476,
    26130 => 19474,
    26131 => 19471,
    26132 => 19469,
    26133 => 19466,
    26134 => 19464,
    26135 => 19461,
    26136 => 19459,
    26137 => 19456,
    26138 => 19454,
    26139 => 19451,
    26140 => 19449,
    26141 => 19446,
    26142 => 19444,
    26143 => 19441,
    26144 => 19438,
    26145 => 19436,
    26146 => 19433,
    26147 => 19431,
    26148 => 19428,
    26149 => 19426,
    26150 => 19423,
    26151 => 19421,
    26152 => 19418,
    26153 => 19416,
    26154 => 19413,
    26155 => 19411,
    26156 => 19408,
    26157 => 19406,
    26158 => 19403,
    26159 => 19400,
    26160 => 19398,
    26161 => 19395,
    26162 => 19393,
    26163 => 19390,
    26164 => 19388,
    26165 => 19385,
    26166 => 19383,
    26167 => 19380,
    26168 => 19378,
    26169 => 19375,
    26170 => 19373,
    26171 => 19370,
    26172 => 19368,
    26173 => 19365,
    26174 => 19362,
    26175 => 19360,
    26176 => 19357,
    26177 => 19355,
    26178 => 19352,
    26179 => 19350,
    26180 => 19347,
    26181 => 19345,
    26182 => 19342,
    26183 => 19340,
    26184 => 19337,
    26185 => 19335,
    26186 => 19332,
    26187 => 19330,
    26188 => 19327,
    26189 => 19324,
    26190 => 19322,
    26191 => 19319,
    26192 => 19317,
    26193 => 19314,
    26194 => 19312,
    26195 => 19309,
    26196 => 19307,
    26197 => 19304,
    26198 => 19302,
    26199 => 19299,
    26200 => 19297,
    26201 => 19294,
    26202 => 19291,
    26203 => 19289,
    26204 => 19286,
    26205 => 19284,
    26206 => 19281,
    26207 => 19279,
    26208 => 19276,
    26209 => 19274,
    26210 => 19271,
    26211 => 19269,
    26212 => 19266,
    26213 => 19264,
    26214 => 19261,
    26215 => 19258,
    26216 => 19256,
    26217 => 19253,
    26218 => 19251,
    26219 => 19248,
    26220 => 19246,
    26221 => 19243,
    26222 => 19241,
    26223 => 19238,
    26224 => 19236,
    26225 => 19233,
    26226 => 19230,
    26227 => 19228,
    26228 => 19225,
    26229 => 19223,
    26230 => 19220,
    26231 => 19218,
    26232 => 19215,
    26233 => 19213,
    26234 => 19210,
    26235 => 19208,
    26236 => 19205,
    26237 => 19202,
    26238 => 19200,
    26239 => 19197,
    26240 => 19195,
    26241 => 19192,
    26242 => 19190,
    26243 => 19187,
    26244 => 19185,
    26245 => 19182,
    26246 => 19180,
    26247 => 19177,
    26248 => 19174,
    26249 => 19172,
    26250 => 19169,
    26251 => 19167,
    26252 => 19164,
    26253 => 19162,
    26254 => 19159,
    26255 => 19157,
    26256 => 19154,
    26257 => 19152,
    26258 => 19149,
    26259 => 19146,
    26260 => 19144,
    26261 => 19141,
    26262 => 19139,
    26263 => 19136,
    26264 => 19134,
    26265 => 19131,
    26266 => 19129,
    26267 => 19126,
    26268 => 19123,
    26269 => 19121,
    26270 => 19118,
    26271 => 19116,
    26272 => 19113,
    26273 => 19111,
    26274 => 19108,
    26275 => 19106,
    26276 => 19103,
    26277 => 19101,
    26278 => 19098,
    26279 => 19095,
    26280 => 19093,
    26281 => 19090,
    26282 => 19088,
    26283 => 19085,
    26284 => 19083,
    26285 => 19080,
    26286 => 19078,
    26287 => 19075,
    26288 => 19072,
    26289 => 19070,
    26290 => 19067,
    26291 => 19065,
    26292 => 19062,
    26293 => 19060,
    26294 => 19057,
    26295 => 19055,
    26296 => 19052,
    26297 => 19049,
    26298 => 19047,
    26299 => 19044,
    26300 => 19042,
    26301 => 19039,
    26302 => 19037,
    26303 => 19034,
    26304 => 19032,
    26305 => 19029,
    26306 => 19026,
    26307 => 19024,
    26308 => 19021,
    26309 => 19019,
    26310 => 19016,
    26311 => 19014,
    26312 => 19011,
    26313 => 19009,
    26314 => 19006,
    26315 => 19003,
    26316 => 19001,
    26317 => 18998,
    26318 => 18996,
    26319 => 18993,
    26320 => 18991,
    26321 => 18988,
    26322 => 18985,
    26323 => 18983,
    26324 => 18980,
    26325 => 18978,
    26326 => 18975,
    26327 => 18973,
    26328 => 18970,
    26329 => 18968,
    26330 => 18965,
    26331 => 18962,
    26332 => 18960,
    26333 => 18957,
    26334 => 18955,
    26335 => 18952,
    26336 => 18950,
    26337 => 18947,
    26338 => 18944,
    26339 => 18942,
    26340 => 18939,
    26341 => 18937,
    26342 => 18934,
    26343 => 18932,
    26344 => 18929,
    26345 => 18927,
    26346 => 18924,
    26347 => 18921,
    26348 => 18919,
    26349 => 18916,
    26350 => 18914,
    26351 => 18911,
    26352 => 18909,
    26353 => 18906,
    26354 => 18903,
    26355 => 18901,
    26356 => 18898,
    26357 => 18896,
    26358 => 18893,
    26359 => 18891,
    26360 => 18888,
    26361 => 18885,
    26362 => 18883,
    26363 => 18880,
    26364 => 18878,
    26365 => 18875,
    26366 => 18873,
    26367 => 18870,
    26368 => 18868,
    26369 => 18865,
    26370 => 18862,
    26371 => 18860,
    26372 => 18857,
    26373 => 18855,
    26374 => 18852,
    26375 => 18850,
    26376 => 18847,
    26377 => 18844,
    26378 => 18842,
    26379 => 18839,
    26380 => 18837,
    26381 => 18834,
    26382 => 18832,
    26383 => 18829,
    26384 => 18826,
    26385 => 18824,
    26386 => 18821,
    26387 => 18819,
    26388 => 18816,
    26389 => 18814,
    26390 => 18811,
    26391 => 18808,
    26392 => 18806,
    26393 => 18803,
    26394 => 18801,
    26395 => 18798,
    26396 => 18796,
    26397 => 18793,
    26398 => 18790,
    26399 => 18788,
    26400 => 18785,
    26401 => 18783,
    26402 => 18780,
    26403 => 18778,
    26404 => 18775,
    26405 => 18772,
    26406 => 18770,
    26407 => 18767,
    26408 => 18765,
    26409 => 18762,
    26410 => 18759,
    26411 => 18757,
    26412 => 18754,
    26413 => 18752,
    26414 => 18749,
    26415 => 18747,
    26416 => 18744,
    26417 => 18741,
    26418 => 18739,
    26419 => 18736,
    26420 => 18734,
    26421 => 18731,
    26422 => 18729,
    26423 => 18726,
    26424 => 18723,
    26425 => 18721,
    26426 => 18718,
    26427 => 18716,
    26428 => 18713,
    26429 => 18711,
    26430 => 18708,
    26431 => 18705,
    26432 => 18703,
    26433 => 18700,
    26434 => 18698,
    26435 => 18695,
    26436 => 18692,
    26437 => 18690,
    26438 => 18687,
    26439 => 18685,
    26440 => 18682,
    26441 => 18680,
    26442 => 18677,
    26443 => 18674,
    26444 => 18672,
    26445 => 18669,
    26446 => 18667,
    26447 => 18664,
    26448 => 18661,
    26449 => 18659,
    26450 => 18656,
    26451 => 18654,
    26452 => 18651,
    26453 => 18649,
    26454 => 18646,
    26455 => 18643,
    26456 => 18641,
    26457 => 18638,
    26458 => 18636,
    26459 => 18633,
    26460 => 18630,
    26461 => 18628,
    26462 => 18625,
    26463 => 18623,
    26464 => 18620,
    26465 => 18618,
    26466 => 18615,
    26467 => 18612,
    26468 => 18610,
    26469 => 18607,
    26470 => 18605,
    26471 => 18602,
    26472 => 18599,
    26473 => 18597,
    26474 => 18594,
    26475 => 18592,
    26476 => 18589,
    26477 => 18587,
    26478 => 18584,
    26479 => 18581,
    26480 => 18579,
    26481 => 18576,
    26482 => 18574,
    26483 => 18571,
    26484 => 18568,
    26485 => 18566,
    26486 => 18563,
    26487 => 18561,
    26488 => 18558,
    26489 => 18555,
    26490 => 18553,
    26491 => 18550,
    26492 => 18548,
    26493 => 18545,
    26494 => 18543,
    26495 => 18540,
    26496 => 18537,
    26497 => 18535,
    26498 => 18532,
    26499 => 18530,
    26500 => 18527,
    26501 => 18524,
    26502 => 18522,
    26503 => 18519,
    26504 => 18517,
    26505 => 18514,
    26506 => 18511,
    26507 => 18509,
    26508 => 18506,
    26509 => 18504,
    26510 => 18501,
    26511 => 18498,
    26512 => 18496,
    26513 => 18493,
    26514 => 18491,
    26515 => 18488,
    26516 => 18485,
    26517 => 18483,
    26518 => 18480,
    26519 => 18478,
    26520 => 18475,
    26521 => 18473,
    26522 => 18470,
    26523 => 18467,
    26524 => 18465,
    26525 => 18462,
    26526 => 18460,
    26527 => 18457,
    26528 => 18454,
    26529 => 18452,
    26530 => 18449,
    26531 => 18447,
    26532 => 18444,
    26533 => 18441,
    26534 => 18439,
    26535 => 18436,
    26536 => 18434,
    26537 => 18431,
    26538 => 18428,
    26539 => 18426,
    26540 => 18423,
    26541 => 18421,
    26542 => 18418,
    26543 => 18415,
    26544 => 18413,
    26545 => 18410,
    26546 => 18408,
    26547 => 18405,
    26548 => 18402,
    26549 => 18400,
    26550 => 18397,
    26551 => 18395,
    26552 => 18392,
    26553 => 18389,
    26554 => 18387,
    26555 => 18384,
    26556 => 18382,
    26557 => 18379,
    26558 => 18376,
    26559 => 18374,
    26560 => 18371,
    26561 => 18369,
    26562 => 18366,
    26563 => 18363,
    26564 => 18361,
    26565 => 18358,
    26566 => 18356,
    26567 => 18353,
    26568 => 18350,
    26569 => 18348,
    26570 => 18345,
    26571 => 18343,
    26572 => 18340,
    26573 => 18337,
    26574 => 18335,
    26575 => 18332,
    26576 => 18330,
    26577 => 18327,
    26578 => 18324,
    26579 => 18322,
    26580 => 18319,
    26581 => 18317,
    26582 => 18314,
    26583 => 18311,
    26584 => 18309,
    26585 => 18306,
    26586 => 18304,
    26587 => 18301,
    26588 => 18298,
    26589 => 18296,
    26590 => 18293,
    26591 => 18290,
    26592 => 18288,
    26593 => 18285,
    26594 => 18283,
    26595 => 18280,
    26596 => 18277,
    26597 => 18275,
    26598 => 18272,
    26599 => 18270,
    26600 => 18267,
    26601 => 18264,
    26602 => 18262,
    26603 => 18259,
    26604 => 18257,
    26605 => 18254,
    26606 => 18251,
    26607 => 18249,
    26608 => 18246,
    26609 => 18244,
    26610 => 18241,
    26611 => 18238,
    26612 => 18236,
    26613 => 18233,
    26614 => 18230,
    26615 => 18228,
    26616 => 18225,
    26617 => 18223,
    26618 => 18220,
    26619 => 18217,
    26620 => 18215,
    26621 => 18212,
    26622 => 18210,
    26623 => 18207,
    26624 => 18204,
    26625 => 18202,
    26626 => 18199,
    26627 => 18197,
    26628 => 18194,
    26629 => 18191,
    26630 => 18189,
    26631 => 18186,
    26632 => 18183,
    26633 => 18181,
    26634 => 18178,
    26635 => 18176,
    26636 => 18173,
    26637 => 18170,
    26638 => 18168,
    26639 => 18165,
    26640 => 18163,
    26641 => 18160,
    26642 => 18157,
    26643 => 18155,
    26644 => 18152,
    26645 => 18149,
    26646 => 18147,
    26647 => 18144,
    26648 => 18142,
    26649 => 18139,
    26650 => 18136,
    26651 => 18134,
    26652 => 18131,
    26653 => 18129,
    26654 => 18126,
    26655 => 18123,
    26656 => 18121,
    26657 => 18118,
    26658 => 18115,
    26659 => 18113,
    26660 => 18110,
    26661 => 18108,
    26662 => 18105,
    26663 => 18102,
    26664 => 18100,
    26665 => 18097,
    26666 => 18095,
    26667 => 18092,
    26668 => 18089,
    26669 => 18087,
    26670 => 18084,
    26671 => 18081,
    26672 => 18079,
    26673 => 18076,
    26674 => 18074,
    26675 => 18071,
    26676 => 18068,
    26677 => 18066,
    26678 => 18063,
    26679 => 18060,
    26680 => 18058,
    26681 => 18055,
    26682 => 18053,
    26683 => 18050,
    26684 => 18047,
    26685 => 18045,
    26686 => 18042,
    26687 => 18039,
    26688 => 18037,
    26689 => 18034,
    26690 => 18032,
    26691 => 18029,
    26692 => 18026,
    26693 => 18024,
    26694 => 18021,
    26695 => 18018,
    26696 => 18016,
    26697 => 18013,
    26698 => 18011,
    26699 => 18008,
    26700 => 18005,
    26701 => 18003,
    26702 => 18000,
    26703 => 17997,
    26704 => 17995,
    26705 => 17992,
    26706 => 17990,
    26707 => 17987,
    26708 => 17984,
    26709 => 17982,
    26710 => 17979,
    26711 => 17976,
    26712 => 17974,
    26713 => 17971,
    26714 => 17969,
    26715 => 17966,
    26716 => 17963,
    26717 => 17961,
    26718 => 17958,
    26719 => 17955,
    26720 => 17953,
    26721 => 17950,
    26722 => 17948,
    26723 => 17945,
    26724 => 17942,
    26725 => 17940,
    26726 => 17937,
    26727 => 17934,
    26728 => 17932,
    26729 => 17929,
    26730 => 17927,
    26731 => 17924,
    26732 => 17921,
    26733 => 17919,
    26734 => 17916,
    26735 => 17913,
    26736 => 17911,
    26737 => 17908,
    26738 => 17906,
    26739 => 17903,
    26740 => 17900,
    26741 => 17898,
    26742 => 17895,
    26743 => 17892,
    26744 => 17890,
    26745 => 17887,
    26746 => 17884,
    26747 => 17882,
    26748 => 17879,
    26749 => 17877,
    26750 => 17874,
    26751 => 17871,
    26752 => 17869,
    26753 => 17866,
    26754 => 17863,
    26755 => 17861,
    26756 => 17858,
    26757 => 17855,
    26758 => 17853,
    26759 => 17850,
    26760 => 17848,
    26761 => 17845,
    26762 => 17842,
    26763 => 17840,
    26764 => 17837,
    26765 => 17834,
    26766 => 17832,
    26767 => 17829,
    26768 => 17827,
    26769 => 17824,
    26770 => 17821,
    26771 => 17819,
    26772 => 17816,
    26773 => 17813,
    26774 => 17811,
    26775 => 17808,
    26776 => 17805,
    26777 => 17803,
    26778 => 17800,
    26779 => 17798,
    26780 => 17795,
    26781 => 17792,
    26782 => 17790,
    26783 => 17787,
    26784 => 17784,
    26785 => 17782,
    26786 => 17779,
    26787 => 17776,
    26788 => 17774,
    26789 => 17771,
    26790 => 17768,
    26791 => 17766,
    26792 => 17763,
    26793 => 17761,
    26794 => 17758,
    26795 => 17755,
    26796 => 17753,
    26797 => 17750,
    26798 => 17747,
    26799 => 17745,
    26800 => 17742,
    26801 => 17739,
    26802 => 17737,
    26803 => 17734,
    26804 => 17732,
    26805 => 17729,
    26806 => 17726,
    26807 => 17724,
    26808 => 17721,
    26809 => 17718,
    26810 => 17716,
    26811 => 17713,
    26812 => 17710,
    26813 => 17708,
    26814 => 17705,
    26815 => 17702,
    26816 => 17700,
    26817 => 17697,
    26818 => 17695,
    26819 => 17692,
    26820 => 17689,
    26821 => 17687,
    26822 => 17684,
    26823 => 17681,
    26824 => 17679,
    26825 => 17676,
    26826 => 17673,
    26827 => 17671,
    26828 => 17668,
    26829 => 17665,
    26830 => 17663,
    26831 => 17660,
    26832 => 17657,
    26833 => 17655,
    26834 => 17652,
    26835 => 17650,
    26836 => 17647,
    26837 => 17644,
    26838 => 17642,
    26839 => 17639,
    26840 => 17636,
    26841 => 17634,
    26842 => 17631,
    26843 => 17628,
    26844 => 17626,
    26845 => 17623,
    26846 => 17620,
    26847 => 17618,
    26848 => 17615,
    26849 => 17612,
    26850 => 17610,
    26851 => 17607,
    26852 => 17605,
    26853 => 17602,
    26854 => 17599,
    26855 => 17597,
    26856 => 17594,
    26857 => 17591,
    26858 => 17589,
    26859 => 17586,
    26860 => 17583,
    26861 => 17581,
    26862 => 17578,
    26863 => 17575,
    26864 => 17573,
    26865 => 17570,
    26866 => 17567,
    26867 => 17565,
    26868 => 17562,
    26869 => 17559,
    26870 => 17557,
    26871 => 17554,
    26872 => 17551,
    26873 => 17549,
    26874 => 17546,
    26875 => 17544,
    26876 => 17541,
    26877 => 17538,
    26878 => 17536,
    26879 => 17533,
    26880 => 17530,
    26881 => 17528,
    26882 => 17525,
    26883 => 17522,
    26884 => 17520,
    26885 => 17517,
    26886 => 17514,
    26887 => 17512,
    26888 => 17509,
    26889 => 17506,
    26890 => 17504,
    26891 => 17501,
    26892 => 17498,
    26893 => 17496,
    26894 => 17493,
    26895 => 17490,
    26896 => 17488,
    26897 => 17485,
    26898 => 17482,
    26899 => 17480,
    26900 => 17477,
    26901 => 17474,
    26902 => 17472,
    26903 => 17469,
    26904 => 17467,
    26905 => 17464,
    26906 => 17461,
    26907 => 17459,
    26908 => 17456,
    26909 => 17453,
    26910 => 17451,
    26911 => 17448,
    26912 => 17445,
    26913 => 17443,
    26914 => 17440,
    26915 => 17437,
    26916 => 17435,
    26917 => 17432,
    26918 => 17429,
    26919 => 17427,
    26920 => 17424,
    26921 => 17421,
    26922 => 17419,
    26923 => 17416,
    26924 => 17413,
    26925 => 17411,
    26926 => 17408,
    26927 => 17405,
    26928 => 17403,
    26929 => 17400,
    26930 => 17397,
    26931 => 17395,
    26932 => 17392,
    26933 => 17389,
    26934 => 17387,
    26935 => 17384,
    26936 => 17381,
    26937 => 17379,
    26938 => 17376,
    26939 => 17373,
    26940 => 17371,
    26941 => 17368,
    26942 => 17365,
    26943 => 17363,
    26944 => 17360,
    26945 => 17357,
    26946 => 17355,
    26947 => 17352,
    26948 => 17349,
    26949 => 17347,
    26950 => 17344,
    26951 => 17341,
    26952 => 17339,
    26953 => 17336,
    26954 => 17333,
    26955 => 17331,
    26956 => 17328,
    26957 => 17325,
    26958 => 17323,
    26959 => 17320,
    26960 => 17317,
    26961 => 17315,
    26962 => 17312,
    26963 => 17309,
    26964 => 17307,
    26965 => 17304,
    26966 => 17301,
    26967 => 17299,
    26968 => 17296,
    26969 => 17293,
    26970 => 17291,
    26971 => 17288,
    26972 => 17285,
    26973 => 17283,
    26974 => 17280,
    26975 => 17277,
    26976 => 17275,
    26977 => 17272,
    26978 => 17269,
    26979 => 17267,
    26980 => 17264,
    26981 => 17261,
    26982 => 17259,
    26983 => 17256,
    26984 => 17253,
    26985 => 17251,
    26986 => 17248,
    26987 => 17245,
    26988 => 17243,
    26989 => 17240,
    26990 => 17237,
    26991 => 17235,
    26992 => 17232,
    26993 => 17229,
    26994 => 17227,
    26995 => 17224,
    26996 => 17221,
    26997 => 17219,
    26998 => 17216,
    26999 => 17213,
    27000 => 17211,
    27001 => 17208,
    27002 => 17205,
    27003 => 17203,
    27004 => 17200,
    27005 => 17197,
    27006 => 17195,
    27007 => 17192,
    27008 => 17189,
    27009 => 17187,
    27010 => 17184,
    27011 => 17181,
    27012 => 17179,
    27013 => 17176,
    27014 => 17173,
    27015 => 17171,
    27016 => 17168,
    27017 => 17165,
    27018 => 17162,
    27019 => 17160,
    27020 => 17157,
    27021 => 17154,
    27022 => 17152,
    27023 => 17149,
    27024 => 17146,
    27025 => 17144,
    27026 => 17141,
    27027 => 17138,
    27028 => 17136,
    27029 => 17133,
    27030 => 17130,
    27031 => 17128,
    27032 => 17125,
    27033 => 17122,
    27034 => 17120,
    27035 => 17117,
    27036 => 17114,
    27037 => 17112,
    27038 => 17109,
    27039 => 17106,
    27040 => 17104,
    27041 => 17101,
    27042 => 17098,
    27043 => 17096,
    27044 => 17093,
    27045 => 17090,
    27046 => 17087,
    27047 => 17085,
    27048 => 17082,
    27049 => 17079,
    27050 => 17077,
    27051 => 17074,
    27052 => 17071,
    27053 => 17069,
    27054 => 17066,
    27055 => 17063,
    27056 => 17061,
    27057 => 17058,
    27058 => 17055,
    27059 => 17053,
    27060 => 17050,
    27061 => 17047,
    27062 => 17045,
    27063 => 17042,
    27064 => 17039,
    27065 => 17037,
    27066 => 17034,
    27067 => 17031,
    27068 => 17028,
    27069 => 17026,
    27070 => 17023,
    27071 => 17020,
    27072 => 17018,
    27073 => 17015,
    27074 => 17012,
    27075 => 17010,
    27076 => 17007,
    27077 => 17004,
    27078 => 17002,
    27079 => 16999,
    27080 => 16996,
    27081 => 16994,
    27082 => 16991,
    27083 => 16988,
    27084 => 16986,
    27085 => 16983,
    27086 => 16980,
    27087 => 16977,
    27088 => 16975,
    27089 => 16972,
    27090 => 16969,
    27091 => 16967,
    27092 => 16964,
    27093 => 16961,
    27094 => 16959,
    27095 => 16956,
    27096 => 16953,
    27097 => 16951,
    27098 => 16948,
    27099 => 16945,
    27100 => 16943,
    27101 => 16940,
    27102 => 16937,
    27103 => 16934,
    27104 => 16932,
    27105 => 16929,
    27106 => 16926,
    27107 => 16924,
    27108 => 16921,
    27109 => 16918,
    27110 => 16916,
    27111 => 16913,
    27112 => 16910,
    27113 => 16908,
    27114 => 16905,
    27115 => 16902,
    27116 => 16899,
    27117 => 16897,
    27118 => 16894,
    27119 => 16891,
    27120 => 16889,
    27121 => 16886,
    27122 => 16883,
    27123 => 16881,
    27124 => 16878,
    27125 => 16875,
    27126 => 16873,
    27127 => 16870,
    27128 => 16867,
    27129 => 16864,
    27130 => 16862,
    27131 => 16859,
    27132 => 16856,
    27133 => 16854,
    27134 => 16851,
    27135 => 16848,
    27136 => 16846,
    27137 => 16843,
    27138 => 16840,
    27139 => 16838,
    27140 => 16835,
    27141 => 16832,
    27142 => 16829,
    27143 => 16827,
    27144 => 16824,
    27145 => 16821,
    27146 => 16819,
    27147 => 16816,
    27148 => 16813,
    27149 => 16811,
    27150 => 16808,
    27151 => 16805,
    27152 => 16802,
    27153 => 16800,
    27154 => 16797,
    27155 => 16794,
    27156 => 16792,
    27157 => 16789,
    27158 => 16786,
    27159 => 16784,
    27160 => 16781,
    27161 => 16778,
    27162 => 16775,
    27163 => 16773,
    27164 => 16770,
    27165 => 16767,
    27166 => 16765,
    27167 => 16762,
    27168 => 16759,
    27169 => 16757,
    27170 => 16754,
    27171 => 16751,
    27172 => 16749,
    27173 => 16746,
    27174 => 16743,
    27175 => 16740,
    27176 => 16738,
    27177 => 16735,
    27178 => 16732,
    27179 => 16730,
    27180 => 16727,
    27181 => 16724,
    27182 => 16721,
    27183 => 16719,
    27184 => 16716,
    27185 => 16713,
    27186 => 16711,
    27187 => 16708,
    27188 => 16705,
    27189 => 16703,
    27190 => 16700,
    27191 => 16697,
    27192 => 16694,
    27193 => 16692,
    27194 => 16689,
    27195 => 16686,
    27196 => 16684,
    27197 => 16681,
    27198 => 16678,
    27199 => 16676,
    27200 => 16673,
    27201 => 16670,
    27202 => 16667,
    27203 => 16665,
    27204 => 16662,
    27205 => 16659,
    27206 => 16657,
    27207 => 16654,
    27208 => 16651,
    27209 => 16648,
    27210 => 16646,
    27211 => 16643,
    27212 => 16640,
    27213 => 16638,
    27214 => 16635,
    27215 => 16632,
    27216 => 16630,
    27217 => 16627,
    27218 => 16624,
    27219 => 16621,
    27220 => 16619,
    27221 => 16616,
    27222 => 16613,
    27223 => 16611,
    27224 => 16608,
    27225 => 16605,
    27226 => 16602,
    27227 => 16600,
    27228 => 16597,
    27229 => 16594,
    27230 => 16592,
    27231 => 16589,
    27232 => 16586,
    27233 => 16584,
    27234 => 16581,
    27235 => 16578,
    27236 => 16575,
    27237 => 16573,
    27238 => 16570,
    27239 => 16567,
    27240 => 16565,
    27241 => 16562,
    27242 => 16559,
    27243 => 16556,
    27244 => 16554,
    27245 => 16551,
    27246 => 16548,
    27247 => 16546,
    27248 => 16543,
    27249 => 16540,
    27250 => 16537,
    27251 => 16535,
    27252 => 16532,
    27253 => 16529,
    27254 => 16527,
    27255 => 16524,
    27256 => 16521,
    27257 => 16518,
    27258 => 16516,
    27259 => 16513,
    27260 => 16510,
    27261 => 16508,
    27262 => 16505,
    27263 => 16502,
    27264 => 16499,
    27265 => 16497,
    27266 => 16494,
    27267 => 16491,
    27268 => 16489,
    27269 => 16486,
    27270 => 16483,
    27271 => 16480,
    27272 => 16478,
    27273 => 16475,
    27274 => 16472,
    27275 => 16470,
    27276 => 16467,
    27277 => 16464,
    27278 => 16461,
    27279 => 16459,
    27280 => 16456,
    27281 => 16453,
    27282 => 16451,
    27283 => 16448,
    27284 => 16445,
    27285 => 16442,
    27286 => 16440,
    27287 => 16437,
    27288 => 16434,
    27289 => 16432,
    27290 => 16429,
    27291 => 16426,
    27292 => 16423,
    27293 => 16421,
    27294 => 16418,
    27295 => 16415,
    27296 => 16413,
    27297 => 16410,
    27298 => 16407,
    27299 => 16404,
    27300 => 16402,
    27301 => 16399,
    27302 => 16396,
    27303 => 16393,
    27304 => 16391,
    27305 => 16388,
    27306 => 16385,
    27307 => 16383,
    27308 => 16380,
    27309 => 16377,
    27310 => 16374,
    27311 => 16372,
    27312 => 16369,
    27313 => 16366,
    27314 => 16364,
    27315 => 16361,
    27316 => 16358,
    27317 => 16355,
    27318 => 16353,
    27319 => 16350,
    27320 => 16347,
    27321 => 16344,
    27322 => 16342,
    27323 => 16339,
    27324 => 16336,
    27325 => 16334,
    27326 => 16331,
    27327 => 16328,
    27328 => 16325,
    27329 => 16323,
    27330 => 16320,
    27331 => 16317,
    27332 => 16315,
    27333 => 16312,
    27334 => 16309,
    27335 => 16306,
    27336 => 16304,
    27337 => 16301,
    27338 => 16298,
    27339 => 16295,
    27340 => 16293,
    27341 => 16290,
    27342 => 16287,
    27343 => 16285,
    27344 => 16282,
    27345 => 16279,
    27346 => 16276,
    27347 => 16274,
    27348 => 16271,
    27349 => 16268,
    27350 => 16265,
    27351 => 16263,
    27352 => 16260,
    27353 => 16257,
    27354 => 16255,
    27355 => 16252,
    27356 => 16249,
    27357 => 16246,
    27358 => 16244,
    27359 => 16241,
    27360 => 16238,
    27361 => 16235,
    27362 => 16233,
    27363 => 16230,
    27364 => 16227,
    27365 => 16225,
    27366 => 16222,
    27367 => 16219,
    27368 => 16216,
    27369 => 16214,
    27370 => 16211,
    27371 => 16208,
    27372 => 16205,
    27373 => 16203,
    27374 => 16200,
    27375 => 16197,
    27376 => 16195,
    27377 => 16192,
    27378 => 16189,
    27379 => 16186,
    27380 => 16184,
    27381 => 16181,
    27382 => 16178,
    27383 => 16175,
    27384 => 16173,
    27385 => 16170,
    27386 => 16167,
    27387 => 16164,
    27388 => 16162,
    27389 => 16159,
    27390 => 16156,
    27391 => 16154,
    27392 => 16151,
    27393 => 16148,
    27394 => 16145,
    27395 => 16143,
    27396 => 16140,
    27397 => 16137,
    27398 => 16134,
    27399 => 16132,
    27400 => 16129,
    27401 => 16126,
    27402 => 16123,
    27403 => 16121,
    27404 => 16118,
    27405 => 16115,
    27406 => 16113,
    27407 => 16110,
    27408 => 16107,
    27409 => 16104,
    27410 => 16102,
    27411 => 16099,
    27412 => 16096,
    27413 => 16093,
    27414 => 16091,
    27415 => 16088,
    27416 => 16085,
    27417 => 16082,
    27418 => 16080,
    27419 => 16077,
    27420 => 16074,
    27421 => 16071,
    27422 => 16069,
    27423 => 16066,
    27424 => 16063,
    27425 => 16061,
    27426 => 16058,
    27427 => 16055,
    27428 => 16052,
    27429 => 16050,
    27430 => 16047,
    27431 => 16044,
    27432 => 16041,
    27433 => 16039,
    27434 => 16036,
    27435 => 16033,
    27436 => 16030,
    27437 => 16028,
    27438 => 16025,
    27439 => 16022,
    27440 => 16019,
    27441 => 16017,
    27442 => 16014,
    27443 => 16011,
    27444 => 16008,
    27445 => 16006,
    27446 => 16003,
    27447 => 16000,
    27448 => 15997,
    27449 => 15995,
    27450 => 15992,
    27451 => 15989,
    27452 => 15987,
    27453 => 15984,
    27454 => 15981,
    27455 => 15978,
    27456 => 15976,
    27457 => 15973,
    27458 => 15970,
    27459 => 15967,
    27460 => 15965,
    27461 => 15962,
    27462 => 15959,
    27463 => 15956,
    27464 => 15954,
    27465 => 15951,
    27466 => 15948,
    27467 => 15945,
    27468 => 15943,
    27469 => 15940,
    27470 => 15937,
    27471 => 15934,
    27472 => 15932,
    27473 => 15929,
    27474 => 15926,
    27475 => 15923,
    27476 => 15921,
    27477 => 15918,
    27478 => 15915,
    27479 => 15912,
    27480 => 15910,
    27481 => 15907,
    27482 => 15904,
    27483 => 15901,
    27484 => 15899,
    27485 => 15896,
    27486 => 15893,
    27487 => 15890,
    27488 => 15888,
    27489 => 15885,
    27490 => 15882,
    27491 => 15879,
    27492 => 15877,
    27493 => 15874,
    27494 => 15871,
    27495 => 15868,
    27496 => 15866,
    27497 => 15863,
    27498 => 15860,
    27499 => 15857,
    27500 => 15855,
    27501 => 15852,
    27502 => 15849,
    27503 => 15846,
    27504 => 15844,
    27505 => 15841,
    27506 => 15838,
    27507 => 15835,
    27508 => 15833,
    27509 => 15830,
    27510 => 15827,
    27511 => 15824,
    27512 => 15822,
    27513 => 15819,
    27514 => 15816,
    27515 => 15813,
    27516 => 15811,
    27517 => 15808,
    27518 => 15805,
    27519 => 15802,
    27520 => 15800,
    27521 => 15797,
    27522 => 15794,
    27523 => 15791,
    27524 => 15789,
    27525 => 15786,
    27526 => 15783,
    27527 => 15780,
    27528 => 15778,
    27529 => 15775,
    27530 => 15772,
    27531 => 15769,
    27532 => 15767,
    27533 => 15764,
    27534 => 15761,
    27535 => 15758,
    27536 => 15756,
    27537 => 15753,
    27538 => 15750,
    27539 => 15747,
    27540 => 15745,
    27541 => 15742,
    27542 => 15739,
    27543 => 15736,
    27544 => 15734,
    27545 => 15731,
    27546 => 15728,
    27547 => 15725,
    27548 => 15723,
    27549 => 15720,
    27550 => 15717,
    27551 => 15714,
    27552 => 15712,
    27553 => 15709,
    27554 => 15706,
    27555 => 15703,
    27556 => 15701,
    27557 => 15698,
    27558 => 15695,
    27559 => 15692,
    27560 => 15690,
    27561 => 15687,
    27562 => 15684,
    27563 => 15681,
    27564 => 15678,
    27565 => 15676,
    27566 => 15673,
    27567 => 15670,
    27568 => 15667,
    27569 => 15665,
    27570 => 15662,
    27571 => 15659,
    27572 => 15656,
    27573 => 15654,
    27574 => 15651,
    27575 => 15648,
    27576 => 15645,
    27577 => 15643,
    27578 => 15640,
    27579 => 15637,
    27580 => 15634,
    27581 => 15632,
    27582 => 15629,
    27583 => 15626,
    27584 => 15623,
    27585 => 15621,
    27586 => 15618,
    27587 => 15615,
    27588 => 15612,
    27589 => 15609,
    27590 => 15607,
    27591 => 15604,
    27592 => 15601,
    27593 => 15598,
    27594 => 15596,
    27595 => 15593,
    27596 => 15590,
    27597 => 15587,
    27598 => 15585,
    27599 => 15582,
    27600 => 15579,
    27601 => 15576,
    27602 => 15574,
    27603 => 15571,
    27604 => 15568,
    27605 => 15565,
    27606 => 15562,
    27607 => 15560,
    27608 => 15557,
    27609 => 15554,
    27610 => 15551,
    27611 => 15549,
    27612 => 15546,
    27613 => 15543,
    27614 => 15540,
    27615 => 15538,
    27616 => 15535,
    27617 => 15532,
    27618 => 15529,
    27619 => 15527,
    27620 => 15524,
    27621 => 15521,
    27622 => 15518,
    27623 => 15515,
    27624 => 15513,
    27625 => 15510,
    27626 => 15507,
    27627 => 15504,
    27628 => 15502,
    27629 => 15499,
    27630 => 15496,
    27631 => 15493,
    27632 => 15491,
    27633 => 15488,
    27634 => 15485,
    27635 => 15482,
    27636 => 15479,
    27637 => 15477,
    27638 => 15474,
    27639 => 15471,
    27640 => 15468,
    27641 => 15466,
    27642 => 15463,
    27643 => 15460,
    27644 => 15457,
    27645 => 15455,
    27646 => 15452,
    27647 => 15449,
    27648 => 15446,
    27649 => 15443,
    27650 => 15441,
    27651 => 15438,
    27652 => 15435,
    27653 => 15432,
    27654 => 15430,
    27655 => 15427,
    27656 => 15424,
    27657 => 15421,
    27658 => 15419,
    27659 => 15416,
    27660 => 15413,
    27661 => 15410,
    27662 => 15407,
    27663 => 15405,
    27664 => 15402,
    27665 => 15399,
    27666 => 15396,
    27667 => 15394,
    27668 => 15391,
    27669 => 15388,
    27670 => 15385,
    27671 => 15382,
    27672 => 15380,
    27673 => 15377,
    27674 => 15374,
    27675 => 15371,
    27676 => 15369,
    27677 => 15366,
    27678 => 15363,
    27679 => 15360,
    27680 => 15358,
    27681 => 15355,
    27682 => 15352,
    27683 => 15349,
    27684 => 15346,
    27685 => 15344,
    27686 => 15341,
    27687 => 15338,
    27688 => 15335,
    27689 => 15333,
    27690 => 15330,
    27691 => 15327,
    27692 => 15324,
    27693 => 15321,
    27694 => 15319,
    27695 => 15316,
    27696 => 15313,
    27697 => 15310,
    27698 => 15308,
    27699 => 15305,
    27700 => 15302,
    27701 => 15299,
    27702 => 15296,
    27703 => 15294,
    27704 => 15291,
    27705 => 15288,
    27706 => 15285,
    27707 => 15283,
    27708 => 15280,
    27709 => 15277,
    27710 => 15274,
    27711 => 15271,
    27712 => 15269,
    27713 => 15266,
    27714 => 15263,
    27715 => 15260,
    27716 => 15258,
    27717 => 15255,
    27718 => 15252,
    27719 => 15249,
    27720 => 15246,
    27721 => 15244,
    27722 => 15241,
    27723 => 15238,
    27724 => 15235,
    27725 => 15233,
    27726 => 15230,
    27727 => 15227,
    27728 => 15224,
    27729 => 15221,
    27730 => 15219,
    27731 => 15216,
    27732 => 15213,
    27733 => 15210,
    27734 => 15207,
    27735 => 15205,
    27736 => 15202,
    27737 => 15199,
    27738 => 15196,
    27739 => 15194,
    27740 => 15191,
    27741 => 15188,
    27742 => 15185,
    27743 => 15182,
    27744 => 15180,
    27745 => 15177,
    27746 => 15174,
    27747 => 15171,
    27748 => 15168,
    27749 => 15166,
    27750 => 15163,
    27751 => 15160,
    27752 => 15157,
    27753 => 15155,
    27754 => 15152,
    27755 => 15149,
    27756 => 15146,
    27757 => 15143,
    27758 => 15141,
    27759 => 15138,
    27760 => 15135,
    27761 => 15132,
    27762 => 15129,
    27763 => 15127,
    27764 => 15124,
    27765 => 15121,
    27766 => 15118,
    27767 => 15116,
    27768 => 15113,
    27769 => 15110,
    27770 => 15107,
    27771 => 15104,
    27772 => 15102,
    27773 => 15099,
    27774 => 15096,
    27775 => 15093,
    27776 => 15090,
    27777 => 15088,
    27778 => 15085,
    27779 => 15082,
    27780 => 15079,
    27781 => 15077,
    27782 => 15074,
    27783 => 15071,
    27784 => 15068,
    27785 => 15065,
    27786 => 15063,
    27787 => 15060,
    27788 => 15057,
    27789 => 15054,
    27790 => 15051,
    27791 => 15049,
    27792 => 15046,
    27793 => 15043,
    27794 => 15040,
    27795 => 15037,
    27796 => 15035,
    27797 => 15032,
    27798 => 15029,
    27799 => 15026,
    27800 => 15024,
    27801 => 15021,
    27802 => 15018,
    27803 => 15015,
    27804 => 15012,
    27805 => 15010,
    27806 => 15007,
    27807 => 15004,
    27808 => 15001,
    27809 => 14998,
    27810 => 14996,
    27811 => 14993,
    27812 => 14990,
    27813 => 14987,
    27814 => 14984,
    27815 => 14982,
    27816 => 14979,
    27817 => 14976,
    27818 => 14973,
    27819 => 14970,
    27820 => 14968,
    27821 => 14965,
    27822 => 14962,
    27823 => 14959,
    27824 => 14956,
    27825 => 14954,
    27826 => 14951,
    27827 => 14948,
    27828 => 14945,
    27829 => 14942,
    27830 => 14940,
    27831 => 14937,
    27832 => 14934,
    27833 => 14931,
    27834 => 14929,
    27835 => 14926,
    27836 => 14923,
    27837 => 14920,
    27838 => 14917,
    27839 => 14915,
    27840 => 14912,
    27841 => 14909,
    27842 => 14906,
    27843 => 14903,
    27844 => 14901,
    27845 => 14898,
    27846 => 14895,
    27847 => 14892,
    27848 => 14889,
    27849 => 14887,
    27850 => 14884,
    27851 => 14881,
    27852 => 14878,
    27853 => 14875,
    27854 => 14873,
    27855 => 14870,
    27856 => 14867,
    27857 => 14864,
    27858 => 14861,
    27859 => 14859,
    27860 => 14856,
    27861 => 14853,
    27862 => 14850,
    27863 => 14847,
    27864 => 14845,
    27865 => 14842,
    27866 => 14839,
    27867 => 14836,
    27868 => 14833,
    27869 => 14831,
    27870 => 14828,
    27871 => 14825,
    27872 => 14822,
    27873 => 14819,
    27874 => 14817,
    27875 => 14814,
    27876 => 14811,
    27877 => 14808,
    27878 => 14805,
    27879 => 14803,
    27880 => 14800,
    27881 => 14797,
    27882 => 14794,
    27883 => 14791,
    27884 => 14789,
    27885 => 14786,
    27886 => 14783,
    27887 => 14780,
    27888 => 14777,
    27889 => 14774,
    27890 => 14772,
    27891 => 14769,
    27892 => 14766,
    27893 => 14763,
    27894 => 14760,
    27895 => 14758,
    27896 => 14755,
    27897 => 14752,
    27898 => 14749,
    27899 => 14746,
    27900 => 14744,
    27901 => 14741,
    27902 => 14738,
    27903 => 14735,
    27904 => 14732,
    27905 => 14730,
    27906 => 14727,
    27907 => 14724,
    27908 => 14721,
    27909 => 14718,
    27910 => 14716,
    27911 => 14713,
    27912 => 14710,
    27913 => 14707,
    27914 => 14704,
    27915 => 14702,
    27916 => 14699,
    27917 => 14696,
    27918 => 14693,
    27919 => 14690,
    27920 => 14688,
    27921 => 14685,
    27922 => 14682,
    27923 => 14679,
    27924 => 14676,
    27925 => 14673,
    27926 => 14671,
    27927 => 14668,
    27928 => 14665,
    27929 => 14662,
    27930 => 14659,
    27931 => 14657,
    27932 => 14654,
    27933 => 14651,
    27934 => 14648,
    27935 => 14645,
    27936 => 14643,
    27937 => 14640,
    27938 => 14637,
    27939 => 14634,
    27940 => 14631,
    27941 => 14628,
    27942 => 14626,
    27943 => 14623,
    27944 => 14620,
    27945 => 14617,
    27946 => 14614,
    27947 => 14612,
    27948 => 14609,
    27949 => 14606,
    27950 => 14603,
    27951 => 14600,
    27952 => 14598,
    27953 => 14595,
    27954 => 14592,
    27955 => 14589,
    27956 => 14586,
    27957 => 14584,
    27958 => 14581,
    27959 => 14578,
    27960 => 14575,
    27961 => 14572,
    27962 => 14569,
    27963 => 14567,
    27964 => 14564,
    27965 => 14561,
    27966 => 14558,
    27967 => 14555,
    27968 => 14553,
    27969 => 14550,
    27970 => 14547,
    27971 => 14544,
    27972 => 14541,
    27973 => 14538,
    27974 => 14536,
    27975 => 14533,
    27976 => 14530,
    27977 => 14527,
    27978 => 14524,
    27979 => 14522,
    27980 => 14519,
    27981 => 14516,
    27982 => 14513,
    27983 => 14510,
    27984 => 14507,
    27985 => 14505,
    27986 => 14502,
    27987 => 14499,
    27988 => 14496,
    27989 => 14493,
    27990 => 14491,
    27991 => 14488,
    27992 => 14485,
    27993 => 14482,
    27994 => 14479,
    27995 => 14477,
    27996 => 14474,
    27997 => 14471,
    27998 => 14468,
    27999 => 14465,
    28000 => 14462,
    28001 => 14460,
    28002 => 14457,
    28003 => 14454,
    28004 => 14451,
    28005 => 14448,
    28006 => 14445,
    28007 => 14443,
    28008 => 14440,
    28009 => 14437,
    28010 => 14434,
    28011 => 14431,
    28012 => 14429,
    28013 => 14426,
    28014 => 14423,
    28015 => 14420,
    28016 => 14417,
    28017 => 14414,
    28018 => 14412,
    28019 => 14409,
    28020 => 14406,
    28021 => 14403,
    28022 => 14400,
    28023 => 14398,
    28024 => 14395,
    28025 => 14392,
    28026 => 14389,
    28027 => 14386,
    28028 => 14383,
    28029 => 14381,
    28030 => 14378,
    28031 => 14375,
    28032 => 14372,
    28033 => 14369,
    28034 => 14366,
    28035 => 14364,
    28036 => 14361,
    28037 => 14358,
    28038 => 14355,
    28039 => 14352,
    28040 => 14350,
    28041 => 14347,
    28042 => 14344,
    28043 => 14341,
    28044 => 14338,
    28045 => 14335,
    28046 => 14333,
    28047 => 14330,
    28048 => 14327,
    28049 => 14324,
    28050 => 14321,
    28051 => 14318,
    28052 => 14316,
    28053 => 14313,
    28054 => 14310,
    28055 => 14307,
    28056 => 14304,
    28057 => 14302,
    28058 => 14299,
    28059 => 14296,
    28060 => 14293,
    28061 => 14290,
    28062 => 14287,
    28063 => 14285,
    28064 => 14282,
    28065 => 14279,
    28066 => 14276,
    28067 => 14273,
    28068 => 14270,
    28069 => 14268,
    28070 => 14265,
    28071 => 14262,
    28072 => 14259,
    28073 => 14256,
    28074 => 14253,
    28075 => 14251,
    28076 => 14248,
    28077 => 14245,
    28078 => 14242,
    28079 => 14239,
    28080 => 14236,
    28081 => 14234,
    28082 => 14231,
    28083 => 14228,
    28084 => 14225,
    28085 => 14222,
    28086 => 14219,
    28087 => 14217,
    28088 => 14214,
    28089 => 14211,
    28090 => 14208,
    28091 => 14205,
    28092 => 14203,
    28093 => 14200,
    28094 => 14197,
    28095 => 14194,
    28096 => 14191,
    28097 => 14188,
    28098 => 14186,
    28099 => 14183,
    28100 => 14180,
    28101 => 14177,
    28102 => 14174,
    28103 => 14171,
    28104 => 14169,
    28105 => 14166,
    28106 => 14163,
    28107 => 14160,
    28108 => 14157,
    28109 => 14154,
    28110 => 14152,
    28111 => 14149,
    28112 => 14146,
    28113 => 14143,
    28114 => 14140,
    28115 => 14137,
    28116 => 14135,
    28117 => 14132,
    28118 => 14129,
    28119 => 14126,
    28120 => 14123,
    28121 => 14120,
    28122 => 14118,
    28123 => 14115,
    28124 => 14112,
    28125 => 14109,
    28126 => 14106,
    28127 => 14103,
    28128 => 14101,
    28129 => 14098,
    28130 => 14095,
    28131 => 14092,
    28132 => 14089,
    28133 => 14086,
    28134 => 14083,
    28135 => 14081,
    28136 => 14078,
    28137 => 14075,
    28138 => 14072,
    28139 => 14069,
    28140 => 14066,
    28141 => 14064,
    28142 => 14061,
    28143 => 14058,
    28144 => 14055,
    28145 => 14052,
    28146 => 14049,
    28147 => 14047,
    28148 => 14044,
    28149 => 14041,
    28150 => 14038,
    28151 => 14035,
    28152 => 14032,
    28153 => 14030,
    28154 => 14027,
    28155 => 14024,
    28156 => 14021,
    28157 => 14018,
    28158 => 14015,
    28159 => 14013,
    28160 => 14010,
    28161 => 14007,
    28162 => 14004,
    28163 => 14001,
    28164 => 13998,
    28165 => 13995,
    28166 => 13993,
    28167 => 13990,
    28168 => 13987,
    28169 => 13984,
    28170 => 13981,
    28171 => 13978,
    28172 => 13976,
    28173 => 13973,
    28174 => 13970,
    28175 => 13967,
    28176 => 13964,
    28177 => 13961,
    28178 => 13959,
    28179 => 13956,
    28180 => 13953,
    28181 => 13950,
    28182 => 13947,
    28183 => 13944,
    28184 => 13942,
    28185 => 13939,
    28186 => 13936,
    28187 => 13933,
    28188 => 13930,
    28189 => 13927,
    28190 => 13924,
    28191 => 13922,
    28192 => 13919,
    28193 => 13916,
    28194 => 13913,
    28195 => 13910,
    28196 => 13907,
    28197 => 13905,
    28198 => 13902,
    28199 => 13899,
    28200 => 13896,
    28201 => 13893,
    28202 => 13890,
    28203 => 13887,
    28204 => 13885,
    28205 => 13882,
    28206 => 13879,
    28207 => 13876,
    28208 => 13873,
    28209 => 13870,
    28210 => 13868,
    28211 => 13865,
    28212 => 13862,
    28213 => 13859,
    28214 => 13856,
    28215 => 13853,
    28216 => 13850,
    28217 => 13848,
    28218 => 13845,
    28219 => 13842,
    28220 => 13839,
    28221 => 13836,
    28222 => 13833,
    28223 => 13831,
    28224 => 13828,
    28225 => 13825,
    28226 => 13822,
    28227 => 13819,
    28228 => 13816,
    28229 => 13813,
    28230 => 13811,
    28231 => 13808,
    28232 => 13805,
    28233 => 13802,
    28234 => 13799,
    28235 => 13796,
    28236 => 13793,
    28237 => 13791,
    28238 => 13788,
    28239 => 13785,
    28240 => 13782,
    28241 => 13779,
    28242 => 13776,
    28243 => 13774,
    28244 => 13771,
    28245 => 13768,
    28246 => 13765,
    28247 => 13762,
    28248 => 13759,
    28249 => 13756,
    28250 => 13754,
    28251 => 13751,
    28252 => 13748,
    28253 => 13745,
    28254 => 13742,
    28255 => 13739,
    28256 => 13736,
    28257 => 13734,
    28258 => 13731,
    28259 => 13728,
    28260 => 13725,
    28261 => 13722,
    28262 => 13719,
    28263 => 13717,
    28264 => 13714,
    28265 => 13711,
    28266 => 13708,
    28267 => 13705,
    28268 => 13702,
    28269 => 13699,
    28270 => 13697,
    28271 => 13694,
    28272 => 13691,
    28273 => 13688,
    28274 => 13685,
    28275 => 13682,
    28276 => 13679,
    28277 => 13677,
    28278 => 13674,
    28279 => 13671,
    28280 => 13668,
    28281 => 13665,
    28282 => 13662,
    28283 => 13659,
    28284 => 13657,
    28285 => 13654,
    28286 => 13651,
    28287 => 13648,
    28288 => 13645,
    28289 => 13642,
    28290 => 13639,
    28291 => 13637,
    28292 => 13634,
    28293 => 13631,
    28294 => 13628,
    28295 => 13625,
    28296 => 13622,
    28297 => 13619,
    28298 => 13617,
    28299 => 13614,
    28300 => 13611,
    28301 => 13608,
    28302 => 13605,
    28303 => 13602,
    28304 => 13599,
    28305 => 13597,
    28306 => 13594,
    28307 => 13591,
    28308 => 13588,
    28309 => 13585,
    28310 => 13582,
    28311 => 13579,
    28312 => 13577,
    28313 => 13574,
    28314 => 13571,
    28315 => 13568,
    28316 => 13565,
    28317 => 13562,
    28318 => 13559,
    28319 => 13557,
    28320 => 13554,
    28321 => 13551,
    28322 => 13548,
    28323 => 13545,
    28324 => 13542,
    28325 => 13539,
    28326 => 13537,
    28327 => 13534,
    28328 => 13531,
    28329 => 13528,
    28330 => 13525,
    28331 => 13522,
    28332 => 13519,
    28333 => 13516,
    28334 => 13514,
    28335 => 13511,
    28336 => 13508,
    28337 => 13505,
    28338 => 13502,
    28339 => 13499,
    28340 => 13496,
    28341 => 13494,
    28342 => 13491,
    28343 => 13488,
    28344 => 13485,
    28345 => 13482,
    28346 => 13479,
    28347 => 13476,
    28348 => 13474,
    28349 => 13471,
    28350 => 13468,
    28351 => 13465,
    28352 => 13462,
    28353 => 13459,
    28354 => 13456,
    28355 => 13454,
    28356 => 13451,
    28357 => 13448,
    28358 => 13445,
    28359 => 13442,
    28360 => 13439,
    28361 => 13436,
    28362 => 13433,
    28363 => 13431,
    28364 => 13428,
    28365 => 13425,
    28366 => 13422,
    28367 => 13419,
    28368 => 13416,
    28369 => 13413,
    28370 => 13411,
    28371 => 13408,
    28372 => 13405,
    28373 => 13402,
    28374 => 13399,
    28375 => 13396,
    28376 => 13393,
    28377 => 13390,
    28378 => 13388,
    28379 => 13385,
    28380 => 13382,
    28381 => 13379,
    28382 => 13376,
    28383 => 13373,
    28384 => 13370,
    28385 => 13368,
    28386 => 13365,
    28387 => 13362,
    28388 => 13359,
    28389 => 13356,
    28390 => 13353,
    28391 => 13350,
    28392 => 13347,
    28393 => 13345,
    28394 => 13342,
    28395 => 13339,
    28396 => 13336,
    28397 => 13333,
    28398 => 13330,
    28399 => 13327,
    28400 => 13324,
    28401 => 13322,
    28402 => 13319,
    28403 => 13316,
    28404 => 13313,
    28405 => 13310,
    28406 => 13307,
    28407 => 13304,
    28408 => 13302,
    28409 => 13299,
    28410 => 13296,
    28411 => 13293,
    28412 => 13290,
    28413 => 13287,
    28414 => 13284,
    28415 => 13281,
    28416 => 13279,
    28417 => 13276,
    28418 => 13273,
    28419 => 13270,
    28420 => 13267,
    28421 => 13264,
    28422 => 13261,
    28423 => 13258,
    28424 => 13256,
    28425 => 13253,
    28426 => 13250,
    28427 => 13247,
    28428 => 13244,
    28429 => 13241,
    28430 => 13238,
    28431 => 13235,
    28432 => 13233,
    28433 => 13230,
    28434 => 13227,
    28435 => 13224,
    28436 => 13221,
    28437 => 13218,
    28438 => 13215,
    28439 => 13212,
    28440 => 13210,
    28441 => 13207,
    28442 => 13204,
    28443 => 13201,
    28444 => 13198,
    28445 => 13195,
    28446 => 13192,
    28447 => 13189,
    28448 => 13187,
    28449 => 13184,
    28450 => 13181,
    28451 => 13178,
    28452 => 13175,
    28453 => 13172,
    28454 => 13169,
    28455 => 13166,
    28456 => 13164,
    28457 => 13161,
    28458 => 13158,
    28459 => 13155,
    28460 => 13152,
    28461 => 13149,
    28462 => 13146,
    28463 => 13143,
    28464 => 13141,
    28465 => 13138,
    28466 => 13135,
    28467 => 13132,
    28468 => 13129,
    28469 => 13126,
    28470 => 13123,
    28471 => 13120,
    28472 => 13118,
    28473 => 13115,
    28474 => 13112,
    28475 => 13109,
    28476 => 13106,
    28477 => 13103,
    28478 => 13100,
    28479 => 13097,
    28480 => 13094,
    28481 => 13092,
    28482 => 13089,
    28483 => 13086,
    28484 => 13083,
    28485 => 13080,
    28486 => 13077,
    28487 => 13074,
    28488 => 13071,
    28489 => 13069,
    28490 => 13066,
    28491 => 13063,
    28492 => 13060,
    28493 => 13057,
    28494 => 13054,
    28495 => 13051,
    28496 => 13048,
    28497 => 13046,
    28498 => 13043,
    28499 => 13040,
    28500 => 13037,
    28501 => 13034,
    28502 => 13031,
    28503 => 13028,
    28504 => 13025,
    28505 => 13022,
    28506 => 13020,
    28507 => 13017,
    28508 => 13014,
    28509 => 13011,
    28510 => 13008,
    28511 => 13005,
    28512 => 13002,
    28513 => 12999,
    28514 => 12997,
    28515 => 12994,
    28516 => 12991,
    28517 => 12988,
    28518 => 12985,
    28519 => 12982,
    28520 => 12979,
    28521 => 12976,
    28522 => 12973,
    28523 => 12971,
    28524 => 12968,
    28525 => 12965,
    28526 => 12962,
    28527 => 12959,
    28528 => 12956,
    28529 => 12953,
    28530 => 12950,
    28531 => 12947,
    28532 => 12945,
    28533 => 12942,
    28534 => 12939,
    28535 => 12936,
    28536 => 12933,
    28537 => 12930,
    28538 => 12927,
    28539 => 12924,
    28540 => 12921,
    28541 => 12919,
    28542 => 12916,
    28543 => 12913,
    28544 => 12910,
    28545 => 12907,
    28546 => 12904,
    28547 => 12901,
    28548 => 12898,
    28549 => 12895,
    28550 => 12893,
    28551 => 12890,
    28552 => 12887,
    28553 => 12884,
    28554 => 12881,
    28555 => 12878,
    28556 => 12875,
    28557 => 12872,
    28558 => 12870,
    28559 => 12867,
    28560 => 12864,
    28561 => 12861,
    28562 => 12858,
    28563 => 12855,
    28564 => 12852,
    28565 => 12849,
    28566 => 12846,
    28567 => 12843,
    28568 => 12841,
    28569 => 12838,
    28570 => 12835,
    28571 => 12832,
    28572 => 12829,
    28573 => 12826,
    28574 => 12823,
    28575 => 12820,
    28576 => 12817,
    28577 => 12815,
    28578 => 12812,
    28579 => 12809,
    28580 => 12806,
    28581 => 12803,
    28582 => 12800,
    28583 => 12797,
    28584 => 12794,
    28585 => 12791,
    28586 => 12789,
    28587 => 12786,
    28588 => 12783,
    28589 => 12780,
    28590 => 12777,
    28591 => 12774,
    28592 => 12771,
    28593 => 12768,
    28594 => 12765,
    28595 => 12763,
    28596 => 12760,
    28597 => 12757,
    28598 => 12754,
    28599 => 12751,
    28600 => 12748,
    28601 => 12745,
    28602 => 12742,
    28603 => 12739,
    28604 => 12736,
    28605 => 12734,
    28606 => 12731,
    28607 => 12728,
    28608 => 12725,
    28609 => 12722,
    28610 => 12719,
    28611 => 12716,
    28612 => 12713,
    28613 => 12710,
    28614 => 12708,
    28615 => 12705,
    28616 => 12702,
    28617 => 12699,
    28618 => 12696,
    28619 => 12693,
    28620 => 12690,
    28621 => 12687,
    28622 => 12684,
    28623 => 12681,
    28624 => 12679,
    28625 => 12676,
    28626 => 12673,
    28627 => 12670,
    28628 => 12667,
    28629 => 12664,
    28630 => 12661,
    28631 => 12658,
    28632 => 12655,
    28633 => 12652,
    28634 => 12650,
    28635 => 12647,
    28636 => 12644,
    28637 => 12641,
    28638 => 12638,
    28639 => 12635,
    28640 => 12632,
    28641 => 12629,
    28642 => 12626,
    28643 => 12624,
    28644 => 12621,
    28645 => 12618,
    28646 => 12615,
    28647 => 12612,
    28648 => 12609,
    28649 => 12606,
    28650 => 12603,
    28651 => 12600,
    28652 => 12597,
    28653 => 12595,
    28654 => 12592,
    28655 => 12589,
    28656 => 12586,
    28657 => 12583,
    28658 => 12580,
    28659 => 12577,
    28660 => 12574,
    28661 => 12571,
    28662 => 12568,
    28663 => 12566,
    28664 => 12563,
    28665 => 12560,
    28666 => 12557,
    28667 => 12554,
    28668 => 12551,
    28669 => 12548,
    28670 => 12545,
    28671 => 12542,
    28672 => 12539,
    28673 => 12536,
    28674 => 12534,
    28675 => 12531,
    28676 => 12528,
    28677 => 12525,
    28678 => 12522,
    28679 => 12519,
    28680 => 12516,
    28681 => 12513,
    28682 => 12510,
    28683 => 12507,
    28684 => 12505,
    28685 => 12502,
    28686 => 12499,
    28687 => 12496,
    28688 => 12493,
    28689 => 12490,
    28690 => 12487,
    28691 => 12484,
    28692 => 12481,
    28693 => 12478,
    28694 => 12476,
    28695 => 12473,
    28696 => 12470,
    28697 => 12467,
    28698 => 12464,
    28699 => 12461,
    28700 => 12458,
    28701 => 12455,
    28702 => 12452,
    28703 => 12449,
    28704 => 12446,
    28705 => 12444,
    28706 => 12441,
    28707 => 12438,
    28708 => 12435,
    28709 => 12432,
    28710 => 12429,
    28711 => 12426,
    28712 => 12423,
    28713 => 12420,
    28714 => 12417,
    28715 => 12414,
    28716 => 12412,
    28717 => 12409,
    28718 => 12406,
    28719 => 12403,
    28720 => 12400,
    28721 => 12397,
    28722 => 12394,
    28723 => 12391,
    28724 => 12388,
    28725 => 12385,
    28726 => 12382,
    28727 => 12380,
    28728 => 12377,
    28729 => 12374,
    28730 => 12371,
    28731 => 12368,
    28732 => 12365,
    28733 => 12362,
    28734 => 12359,
    28735 => 12356,
    28736 => 12353,
    28737 => 12350,
    28738 => 12348,
    28739 => 12345,
    28740 => 12342,
    28741 => 12339,
    28742 => 12336,
    28743 => 12333,
    28744 => 12330,
    28745 => 12327,
    28746 => 12324,
    28747 => 12321,
    28748 => 12318,
    28749 => 12316,
    28750 => 12313,
    28751 => 12310,
    28752 => 12307,
    28753 => 12304,
    28754 => 12301,
    28755 => 12298,
    28756 => 12295,
    28757 => 12292,
    28758 => 12289,
    28759 => 12286,
    28760 => 12284,
    28761 => 12281,
    28762 => 12278,
    28763 => 12275,
    28764 => 12272,
    28765 => 12269,
    28766 => 12266,
    28767 => 12263,
    28768 => 12260,
    28769 => 12257,
    28770 => 12254,
    28771 => 12251,
    28772 => 12249,
    28773 => 12246,
    28774 => 12243,
    28775 => 12240,
    28776 => 12237,
    28777 => 12234,
    28778 => 12231,
    28779 => 12228,
    28780 => 12225,
    28781 => 12222,
    28782 => 12219,
    28783 => 12217,
    28784 => 12214,
    28785 => 12211,
    28786 => 12208,
    28787 => 12205,
    28788 => 12202,
    28789 => 12199,
    28790 => 12196,
    28791 => 12193,
    28792 => 12190,
    28793 => 12187,
    28794 => 12184,
    28795 => 12182,
    28796 => 12179,
    28797 => 12176,
    28798 => 12173,
    28799 => 12170,
    28800 => 12167,
    28801 => 12164,
    28802 => 12161,
    28803 => 12158,
    28804 => 12155,
    28805 => 12152,
    28806 => 12149,
    28807 => 12147,
    28808 => 12144,
    28809 => 12141,
    28810 => 12138,
    28811 => 12135,
    28812 => 12132,
    28813 => 12129,
    28814 => 12126,
    28815 => 12123,
    28816 => 12120,
    28817 => 12117,
    28818 => 12114,
    28819 => 12112,
    28820 => 12109,
    28821 => 12106,
    28822 => 12103,
    28823 => 12100,
    28824 => 12097,
    28825 => 12094,
    28826 => 12091,
    28827 => 12088,
    28828 => 12085,
    28829 => 12082,
    28830 => 12079,
    28831 => 12076,
    28832 => 12074,
    28833 => 12071,
    28834 => 12068,
    28835 => 12065,
    28836 => 12062,
    28837 => 12059,
    28838 => 12056,
    28839 => 12053,
    28840 => 12050,
    28841 => 12047,
    28842 => 12044,
    28843 => 12041,
    28844 => 12038,
    28845 => 12036,
    28846 => 12033,
    28847 => 12030,
    28848 => 12027,
    28849 => 12024,
    28850 => 12021,
    28851 => 12018,
    28852 => 12015,
    28853 => 12012,
    28854 => 12009,
    28855 => 12006,
    28856 => 12003,
    28857 => 12001,
    28858 => 11998,
    28859 => 11995,
    28860 => 11992,
    28861 => 11989,
    28862 => 11986,
    28863 => 11983,
    28864 => 11980,
    28865 => 11977,
    28866 => 11974,
    28867 => 11971,
    28868 => 11968,
    28869 => 11965,
    28870 => 11962,
    28871 => 11960,
    28872 => 11957,
    28873 => 11954,
    28874 => 11951,
    28875 => 11948,
    28876 => 11945,
    28877 => 11942,
    28878 => 11939,
    28879 => 11936,
    28880 => 11933,
    28881 => 11930,
    28882 => 11927,
    28883 => 11924,
    28884 => 11922,
    28885 => 11919,
    28886 => 11916,
    28887 => 11913,
    28888 => 11910,
    28889 => 11907,
    28890 => 11904,
    28891 => 11901,
    28892 => 11898,
    28893 => 11895,
    28894 => 11892,
    28895 => 11889,
    28896 => 11886,
    28897 => 11883,
    28898 => 11881,
    28899 => 11878,
    28900 => 11875,
    28901 => 11872,
    28902 => 11869,
    28903 => 11866,
    28904 => 11863,
    28905 => 11860,
    28906 => 11857,
    28907 => 11854,
    28908 => 11851,
    28909 => 11848,
    28910 => 11845,
    28911 => 11842,
    28912 => 11840,
    28913 => 11837,
    28914 => 11834,
    28915 => 11831,
    28916 => 11828,
    28917 => 11825,
    28918 => 11822,
    28919 => 11819,
    28920 => 11816,
    28921 => 11813,
    28922 => 11810,
    28923 => 11807,
    28924 => 11804,
    28925 => 11801,
    28926 => 11799,
    28927 => 11796,
    28928 => 11793,
    28929 => 11790,
    28930 => 11787,
    28931 => 11784,
    28932 => 11781,
    28933 => 11778,
    28934 => 11775,
    28935 => 11772,
    28936 => 11769,
    28937 => 11766,
    28938 => 11763,
    28939 => 11760,
    28940 => 11758,
    28941 => 11755,
    28942 => 11752,
    28943 => 11749,
    28944 => 11746,
    28945 => 11743,
    28946 => 11740,
    28947 => 11737,
    28948 => 11734,
    28949 => 11731,
    28950 => 11728,
    28951 => 11725,
    28952 => 11722,
    28953 => 11719,
    28954 => 11716,
    28955 => 11714,
    28956 => 11711,
    28957 => 11708,
    28958 => 11705,
    28959 => 11702,
    28960 => 11699,
    28961 => 11696,
    28962 => 11693,
    28963 => 11690,
    28964 => 11687,
    28965 => 11684,
    28966 => 11681,
    28967 => 11678,
    28968 => 11675,
    28969 => 11672,
    28970 => 11669,
    28971 => 11667,
    28972 => 11664,
    28973 => 11661,
    28974 => 11658,
    28975 => 11655,
    28976 => 11652,
    28977 => 11649,
    28978 => 11646,
    28979 => 11643,
    28980 => 11640,
    28981 => 11637,
    28982 => 11634,
    28983 => 11631,
    28984 => 11628,
    28985 => 11625,
    28986 => 11623,
    28987 => 11620,
    28988 => 11617,
    28989 => 11614,
    28990 => 11611,
    28991 => 11608,
    28992 => 11605,
    28993 => 11602,
    28994 => 11599,
    28995 => 11596,
    28996 => 11593,
    28997 => 11590,
    28998 => 11587,
    28999 => 11584,
    29000 => 11581,
    29001 => 11578,
    29002 => 11575,
    29003 => 11573,
    29004 => 11570,
    29005 => 11567,
    29006 => 11564,
    29007 => 11561,
    29008 => 11558,
    29009 => 11555,
    29010 => 11552,
    29011 => 11549,
    29012 => 11546,
    29013 => 11543,
    29014 => 11540,
    29015 => 11537,
    29016 => 11534,
    29017 => 11531,
    29018 => 11528,
    29019 => 11526,
    29020 => 11523,
    29021 => 11520,
    29022 => 11517,
    29023 => 11514,
    29024 => 11511,
    29025 => 11508,
    29026 => 11505,
    29027 => 11502,
    29028 => 11499,
    29029 => 11496,
    29030 => 11493,
    29031 => 11490,
    29032 => 11487,
    29033 => 11484,
    29034 => 11481,
    29035 => 11478,
    29036 => 11476,
    29037 => 11473,
    29038 => 11470,
    29039 => 11467,
    29040 => 11464,
    29041 => 11461,
    29042 => 11458,
    29043 => 11455,
    29044 => 11452,
    29045 => 11449,
    29046 => 11446,
    29047 => 11443,
    29048 => 11440,
    29049 => 11437,
    29050 => 11434,
    29051 => 11431,
    29052 => 11428,
    29053 => 11425,
    29054 => 11423,
    29055 => 11420,
    29056 => 11417,
    29057 => 11414,
    29058 => 11411,
    29059 => 11408,
    29060 => 11405,
    29061 => 11402,
    29062 => 11399,
    29063 => 11396,
    29064 => 11393,
    29065 => 11390,
    29066 => 11387,
    29067 => 11384,
    29068 => 11381,
    29069 => 11378,
    29070 => 11375,
    29071 => 11372,
    29072 => 11370,
    29073 => 11367,
    29074 => 11364,
    29075 => 11361,
    29076 => 11358,
    29077 => 11355,
    29078 => 11352,
    29079 => 11349,
    29080 => 11346,
    29081 => 11343,
    29082 => 11340,
    29083 => 11337,
    29084 => 11334,
    29085 => 11331,
    29086 => 11328,
    29087 => 11325,
    29088 => 11322,
    29089 => 11319,
    29090 => 11316,
    29091 => 11314,
    29092 => 11311,
    29093 => 11308,
    29094 => 11305,
    29095 => 11302,
    29096 => 11299,
    29097 => 11296,
    29098 => 11293,
    29099 => 11290,
    29100 => 11287,
    29101 => 11284,
    29102 => 11281,
    29103 => 11278,
    29104 => 11275,
    29105 => 11272,
    29106 => 11269,
    29107 => 11266,
    29108 => 11263,
    29109 => 11260,
    29110 => 11257,
    29111 => 11255,
    29112 => 11252,
    29113 => 11249,
    29114 => 11246,
    29115 => 11243,
    29116 => 11240,
    29117 => 11237,
    29118 => 11234,
    29119 => 11231,
    29120 => 11228,
    29121 => 11225,
    29122 => 11222,
    29123 => 11219,
    29124 => 11216,
    29125 => 11213,
    29126 => 11210,
    29127 => 11207,
    29128 => 11204,
    29129 => 11201,
    29130 => 11198,
    29131 => 11195,
    29132 => 11193,
    29133 => 11190,
    29134 => 11187,
    29135 => 11184,
    29136 => 11181,
    29137 => 11178,
    29138 => 11175,
    29139 => 11172,
    29140 => 11169,
    29141 => 11166,
    29142 => 11163,
    29143 => 11160,
    29144 => 11157,
    29145 => 11154,
    29146 => 11151,
    29147 => 11148,
    29148 => 11145,
    29149 => 11142,
    29150 => 11139,
    29151 => 11136,
    29152 => 11133,
    29153 => 11131,
    29154 => 11128,
    29155 => 11125,
    29156 => 11122,
    29157 => 11119,
    29158 => 11116,
    29159 => 11113,
    29160 => 11110,
    29161 => 11107,
    29162 => 11104,
    29163 => 11101,
    29164 => 11098,
    29165 => 11095,
    29166 => 11092,
    29167 => 11089,
    29168 => 11086,
    29169 => 11083,
    29170 => 11080,
    29171 => 11077,
    29172 => 11074,
    29173 => 11071,
    29174 => 11068,
    29175 => 11065,
    29176 => 11063,
    29177 => 11060,
    29178 => 11057,
    29179 => 11054,
    29180 => 11051,
    29181 => 11048,
    29182 => 11045,
    29183 => 11042,
    29184 => 11039,
    29185 => 11036,
    29186 => 11033,
    29187 => 11030,
    29188 => 11027,
    29189 => 11024,
    29190 => 11021,
    29191 => 11018,
    29192 => 11015,
    29193 => 11012,
    29194 => 11009,
    29195 => 11006,
    29196 => 11003,
    29197 => 11000,
    29198 => 10997,
    29199 => 10994,
    29200 => 10992,
    29201 => 10989,
    29202 => 10986,
    29203 => 10983,
    29204 => 10980,
    29205 => 10977,
    29206 => 10974,
    29207 => 10971,
    29208 => 10968,
    29209 => 10965,
    29210 => 10962,
    29211 => 10959,
    29212 => 10956,
    29213 => 10953,
    29214 => 10950,
    29215 => 10947,
    29216 => 10944,
    29217 => 10941,
    29218 => 10938,
    29219 => 10935,
    29220 => 10932,
    29221 => 10929,
    29222 => 10926,
    29223 => 10923,
    29224 => 10920,
    29225 => 10918,
    29226 => 10915,
    29227 => 10912,
    29228 => 10909,
    29229 => 10906,
    29230 => 10903,
    29231 => 10900,
    29232 => 10897,
    29233 => 10894,
    29234 => 10891,
    29235 => 10888,
    29236 => 10885,
    29237 => 10882,
    29238 => 10879,
    29239 => 10876,
    29240 => 10873,
    29241 => 10870,
    29242 => 10867,
    29243 => 10864,
    29244 => 10861,
    29245 => 10858,
    29246 => 10855,
    29247 => 10852,
    29248 => 10849,
    29249 => 10846,
    29250 => 10843,
    29251 => 10840,
    29252 => 10838,
    29253 => 10835,
    29254 => 10832,
    29255 => 10829,
    29256 => 10826,
    29257 => 10823,
    29258 => 10820,
    29259 => 10817,
    29260 => 10814,
    29261 => 10811,
    29262 => 10808,
    29263 => 10805,
    29264 => 10802,
    29265 => 10799,
    29266 => 10796,
    29267 => 10793,
    29268 => 10790,
    29269 => 10787,
    29270 => 10784,
    29271 => 10781,
    29272 => 10778,
    29273 => 10775,
    29274 => 10772,
    29275 => 10769,
    29276 => 10766,
    29277 => 10763,
    29278 => 10760,
    29279 => 10757,
    29280 => 10754,
    29281 => 10751,
    29282 => 10749,
    29283 => 10746,
    29284 => 10743,
    29285 => 10740,
    29286 => 10737,
    29287 => 10734,
    29288 => 10731,
    29289 => 10728,
    29290 => 10725,
    29291 => 10722,
    29292 => 10719,
    29293 => 10716,
    29294 => 10713,
    29295 => 10710,
    29296 => 10707,
    29297 => 10704,
    29298 => 10701,
    29299 => 10698,
    29300 => 10695,
    29301 => 10692,
    29302 => 10689,
    29303 => 10686,
    29304 => 10683,
    29305 => 10680,
    29306 => 10677,
    29307 => 10674,
    29308 => 10671,
    29309 => 10668,
    29310 => 10665,
    29311 => 10662,
    29312 => 10659,
    29313 => 10656,
    29314 => 10654,
    29315 => 10651,
    29316 => 10648,
    29317 => 10645,
    29318 => 10642,
    29319 => 10639,
    29320 => 10636,
    29321 => 10633,
    29322 => 10630,
    29323 => 10627,
    29324 => 10624,
    29325 => 10621,
    29326 => 10618,
    29327 => 10615,
    29328 => 10612,
    29329 => 10609,
    29330 => 10606,
    29331 => 10603,
    29332 => 10600,
    29333 => 10597,
    29334 => 10594,
    29335 => 10591,
    29336 => 10588,
    29337 => 10585,
    29338 => 10582,
    29339 => 10579,
    29340 => 10576,
    29341 => 10573,
    29342 => 10570,
    29343 => 10567,
    29344 => 10564,
    29345 => 10561,
    29346 => 10558,
    29347 => 10555,
    29348 => 10552,
    29349 => 10549,
    29350 => 10546,
    29351 => 10544,
    29352 => 10541,
    29353 => 10538,
    29354 => 10535,
    29355 => 10532,
    29356 => 10529,
    29357 => 10526,
    29358 => 10523,
    29359 => 10520,
    29360 => 10517,
    29361 => 10514,
    29362 => 10511,
    29363 => 10508,
    29364 => 10505,
    29365 => 10502,
    29366 => 10499,
    29367 => 10496,
    29368 => 10493,
    29369 => 10490,
    29370 => 10487,
    29371 => 10484,
    29372 => 10481,
    29373 => 10478,
    29374 => 10475,
    29375 => 10472,
    29376 => 10469,
    29377 => 10466,
    29378 => 10463,
    29379 => 10460,
    29380 => 10457,
    29381 => 10454,
    29382 => 10451,
    29383 => 10448,
    29384 => 10445,
    29385 => 10442,
    29386 => 10439,
    29387 => 10436,
    29388 => 10433,
    29389 => 10430,
    29390 => 10427,
    29391 => 10424,
    29392 => 10421,
    29393 => 10419,
    29394 => 10416,
    29395 => 10413,
    29396 => 10410,
    29397 => 10407,
    29398 => 10404,
    29399 => 10401,
    29400 => 10398,
    29401 => 10395,
    29402 => 10392,
    29403 => 10389,
    29404 => 10386,
    29405 => 10383,
    29406 => 10380,
    29407 => 10377,
    29408 => 10374,
    29409 => 10371,
    29410 => 10368,
    29411 => 10365,
    29412 => 10362,
    29413 => 10359,
    29414 => 10356,
    29415 => 10353,
    29416 => 10350,
    29417 => 10347,
    29418 => 10344,
    29419 => 10341,
    29420 => 10338,
    29421 => 10335,
    29422 => 10332,
    29423 => 10329,
    29424 => 10326,
    29425 => 10323,
    29426 => 10320,
    29427 => 10317,
    29428 => 10314,
    29429 => 10311,
    29430 => 10308,
    29431 => 10305,
    29432 => 10302,
    29433 => 10299,
    29434 => 10296,
    29435 => 10293,
    29436 => 10290,
    29437 => 10287,
    29438 => 10284,
    29439 => 10281,
    29440 => 10278,
    29441 => 10275,
    29442 => 10272,
    29443 => 10269,
    29444 => 10266,
    29445 => 10263,
    29446 => 10261,
    29447 => 10258,
    29448 => 10255,
    29449 => 10252,
    29450 => 10249,
    29451 => 10246,
    29452 => 10243,
    29453 => 10240,
    29454 => 10237,
    29455 => 10234,
    29456 => 10231,
    29457 => 10228,
    29458 => 10225,
    29459 => 10222,
    29460 => 10219,
    29461 => 10216,
    29462 => 10213,
    29463 => 10210,
    29464 => 10207,
    29465 => 10204,
    29466 => 10201,
    29467 => 10198,
    29468 => 10195,
    29469 => 10192,
    29470 => 10189,
    29471 => 10186,
    29472 => 10183,
    29473 => 10180,
    29474 => 10177,
    29475 => 10174,
    29476 => 10171,
    29477 => 10168,
    29478 => 10165,
    29479 => 10162,
    29480 => 10159,
    29481 => 10156,
    29482 => 10153,
    29483 => 10150,
    29484 => 10147,
    29485 => 10144,
    29486 => 10141,
    29487 => 10138,
    29488 => 10135,
    29489 => 10132,
    29490 => 10129,
    29491 => 10126,
    29492 => 10123,
    29493 => 10120,
    29494 => 10117,
    29495 => 10114,
    29496 => 10111,
    29497 => 10108,
    29498 => 10105,
    29499 => 10102,
    29500 => 10099,
    29501 => 10096,
    29502 => 10093,
    29503 => 10090,
    29504 => 10087,
    29505 => 10084,
    29506 => 10081,
    29507 => 10078,
    29508 => 10075,
    29509 => 10072,
    29510 => 10069,
    29511 => 10066,
    29512 => 10063,
    29513 => 10060,
    29514 => 10057,
    29515 => 10054,
    29516 => 10051,
    29517 => 10048,
    29518 => 10045,
    29519 => 10042,
    29520 => 10039,
    29521 => 10036,
    29522 => 10033,
    29523 => 10031,
    29524 => 10028,
    29525 => 10025,
    29526 => 10022,
    29527 => 10019,
    29528 => 10016,
    29529 => 10013,
    29530 => 10010,
    29531 => 10007,
    29532 => 10004,
    29533 => 10001,
    29534 => 9998,
    29535 => 9995,
    29536 => 9992,
    29537 => 9989,
    29538 => 9986,
    29539 => 9983,
    29540 => 9980,
    29541 => 9977,
    29542 => 9974,
    29543 => 9971,
    29544 => 9968,
    29545 => 9965,
    29546 => 9962,
    29547 => 9959,
    29548 => 9956,
    29549 => 9953,
    29550 => 9950,
    29551 => 9947,
    29552 => 9944,
    29553 => 9941,
    29554 => 9938,
    29555 => 9935,
    29556 => 9932,
    29557 => 9929,
    29558 => 9926,
    29559 => 9923,
    29560 => 9920,
    29561 => 9917,
    29562 => 9914,
    29563 => 9911,
    29564 => 9908,
    29565 => 9905,
    29566 => 9902,
    29567 => 9899,
    29568 => 9896,
    29569 => 9893,
    29570 => 9890,
    29571 => 9887,
    29572 => 9884,
    29573 => 9881,
    29574 => 9878,
    29575 => 9875,
    29576 => 9872,
    29577 => 9869,
    29578 => 9866,
    29579 => 9863,
    29580 => 9860,
    29581 => 9857,
    29582 => 9854,
    29583 => 9851,
    29584 => 9848,
    29585 => 9845,
    29586 => 9842,
    29587 => 9839,
    29588 => 9836,
    29589 => 9833,
    29590 => 9830,
    29591 => 9827,
    29592 => 9824,
    29593 => 9821,
    29594 => 9818,
    29595 => 9815,
    29596 => 9812,
    29597 => 9809,
    29598 => 9806,
    29599 => 9803,
    29600 => 9800,
    29601 => 9797,
    29602 => 9794,
    29603 => 9791,
    29604 => 9788,
    29605 => 9785,
    29606 => 9782,
    29607 => 9779,
    29608 => 9776,
    29609 => 9773,
    29610 => 9770,
    29611 => 9767,
    29612 => 9764,
    29613 => 9761,
    29614 => 9758,
    29615 => 9755,
    29616 => 9752,
    29617 => 9749,
    29618 => 9746,
    29619 => 9743,
    29620 => 9740,
    29621 => 9737,
    29622 => 9734,
    29623 => 9731,
    29624 => 9728,
    29625 => 9725,
    29626 => 9722,
    29627 => 9719,
    29628 => 9716,
    29629 => 9713,
    29630 => 9710,
    29631 => 9707,
    29632 => 9704,
    29633 => 9701,
    29634 => 9698,
    29635 => 9695,
    29636 => 9692,
    29637 => 9689,
    29638 => 9686,
    29639 => 9683,
    29640 => 9680,
    29641 => 9677,
    29642 => 9674,
    29643 => 9671,
    29644 => 9668,
    29645 => 9665,
    29646 => 9662,
    29647 => 9659,
    29648 => 9656,
    29649 => 9653,
    29650 => 9650,
    29651 => 9647,
    29652 => 9644,
    29653 => 9641,
    29654 => 9638,
    29655 => 9635,
    29656 => 9632,
    29657 => 9629,
    29658 => 9626,
    29659 => 9623,
    29660 => 9620,
    29661 => 9617,
    29662 => 9614,
    29663 => 9611,
    29664 => 9608,
    29665 => 9605,
    29666 => 9602,
    29667 => 9599,
    29668 => 9596,
    29669 => 9593,
    29670 => 9590,
    29671 => 9587,
    29672 => 9584,
    29673 => 9581,
    29674 => 9578,
    29675 => 9575,
    29676 => 9572,
    29677 => 9569,
    29678 => 9566,
    29679 => 9563,
    29680 => 9560,
    29681 => 9557,
    29682 => 9554,
    29683 => 9551,
    29684 => 9548,
    29685 => 9545,
    29686 => 9542,
    29687 => 9539,
    29688 => 9536,
    29689 => 9533,
    29690 => 9530,
    29691 => 9527,
    29692 => 9524,
    29693 => 9521,
    29694 => 9518,
    29695 => 9515,
    29696 => 9512,
    29697 => 9509,
    29698 => 9506,
    29699 => 9503,
    29700 => 9500,
    29701 => 9497,
    29702 => 9494,
    29703 => 9491,
    29704 => 9488,
    29705 => 9485,
    29706 => 9482,
    29707 => 9479,
    29708 => 9476,
    29709 => 9473,
    29710 => 9470,
    29711 => 9467,
    29712 => 9464,
    29713 => 9461,
    29714 => 9458,
    29715 => 9455,
    29716 => 9452,
    29717 => 9449,
    29718 => 9446,
    29719 => 9443,
    29720 => 9440,
    29721 => 9437,
    29722 => 9434,
    29723 => 9431,
    29724 => 9428,
    29725 => 9425,
    29726 => 9422,
    29727 => 9419,
    29728 => 9416,
    29729 => 9413,
    29730 => 9409,
    29731 => 9406,
    29732 => 9403,
    29733 => 9400,
    29734 => 9397,
    29735 => 9394,
    29736 => 9391,
    29737 => 9388,
    29738 => 9385,
    29739 => 9382,
    29740 => 9379,
    29741 => 9376,
    29742 => 9373,
    29743 => 9370,
    29744 => 9367,
    29745 => 9364,
    29746 => 9361,
    29747 => 9358,
    29748 => 9355,
    29749 => 9352,
    29750 => 9349,
    29751 => 9346,
    29752 => 9343,
    29753 => 9340,
    29754 => 9337,
    29755 => 9334,
    29756 => 9331,
    29757 => 9328,
    29758 => 9325,
    29759 => 9322,
    29760 => 9319,
    29761 => 9316,
    29762 => 9313,
    29763 => 9310,
    29764 => 9307,
    29765 => 9304,
    29766 => 9301,
    29767 => 9298,
    29768 => 9295,
    29769 => 9292,
    29770 => 9289,
    29771 => 9286,
    29772 => 9283,
    29773 => 9280,
    29774 => 9277,
    29775 => 9274,
    29776 => 9271,
    29777 => 9268,
    29778 => 9265,
    29779 => 9262,
    29780 => 9259,
    29781 => 9256,
    29782 => 9253,
    29783 => 9250,
    29784 => 9247,
    29785 => 9244,
    29786 => 9241,
    29787 => 9238,
    29788 => 9235,
    29789 => 9232,
    29790 => 9229,
    29791 => 9226,
    29792 => 9223,
    29793 => 9220,
    29794 => 9217,
    29795 => 9214,
    29796 => 9211,
    29797 => 9208,
    29798 => 9205,
    29799 => 9202,
    29800 => 9199,
    29801 => 9196,
    29802 => 9193,
    29803 => 9190,
    29804 => 9187,
    29805 => 9184,
    29806 => 9181,
    29807 => 9178,
    29808 => 9175,
    29809 => 9172,
    29810 => 9168,
    29811 => 9165,
    29812 => 9162,
    29813 => 9159,
    29814 => 9156,
    29815 => 9153,
    29816 => 9150,
    29817 => 9147,
    29818 => 9144,
    29819 => 9141,
    29820 => 9138,
    29821 => 9135,
    29822 => 9132,
    29823 => 9129,
    29824 => 9126,
    29825 => 9123,
    29826 => 9120,
    29827 => 9117,
    29828 => 9114,
    29829 => 9111,
    29830 => 9108,
    29831 => 9105,
    29832 => 9102,
    29833 => 9099,
    29834 => 9096,
    29835 => 9093,
    29836 => 9090,
    29837 => 9087,
    29838 => 9084,
    29839 => 9081,
    29840 => 9078,
    29841 => 9075,
    29842 => 9072,
    29843 => 9069,
    29844 => 9066,
    29845 => 9063,
    29846 => 9060,
    29847 => 9057,
    29848 => 9054,
    29849 => 9051,
    29850 => 9048,
    29851 => 9045,
    29852 => 9042,
    29853 => 9039,
    29854 => 9036,
    29855 => 9033,
    29856 => 9030,
    29857 => 9027,
    29858 => 9024,
    29859 => 9021,
    29860 => 9018,
    29861 => 9015,
    29862 => 9012,
    29863 => 9009,
    29864 => 9006,
    29865 => 9002,
    29866 => 8999,
    29867 => 8996,
    29868 => 8993,
    29869 => 8990,
    29870 => 8987,
    29871 => 8984,
    29872 => 8981,
    29873 => 8978,
    29874 => 8975,
    29875 => 8972,
    29876 => 8969,
    29877 => 8966,
    29878 => 8963,
    29879 => 8960,
    29880 => 8957,
    29881 => 8954,
    29882 => 8951,
    29883 => 8948,
    29884 => 8945,
    29885 => 8942,
    29886 => 8939,
    29887 => 8936,
    29888 => 8933,
    29889 => 8930,
    29890 => 8927,
    29891 => 8924,
    29892 => 8921,
    29893 => 8918,
    29894 => 8915,
    29895 => 8912,
    29896 => 8909,
    29897 => 8906,
    29898 => 8903,
    29899 => 8900,
    29900 => 8897,
    29901 => 8894,
    29902 => 8891,
    29903 => 8888,
    29904 => 8885,
    29905 => 8882,
    29906 => 8879,
    29907 => 8876,
    29908 => 8873,
    29909 => 8869,
    29910 => 8866,
    29911 => 8863,
    29912 => 8860,
    29913 => 8857,
    29914 => 8854,
    29915 => 8851,
    29916 => 8848,
    29917 => 8845,
    29918 => 8842,
    29919 => 8839,
    29920 => 8836,
    29921 => 8833,
    29922 => 8830,
    29923 => 8827,
    29924 => 8824,
    29925 => 8821,
    29926 => 8818,
    29927 => 8815,
    29928 => 8812,
    29929 => 8809,
    29930 => 8806,
    29931 => 8803,
    29932 => 8800,
    29933 => 8797,
    29934 => 8794,
    29935 => 8791,
    29936 => 8788,
    29937 => 8785,
    29938 => 8782,
    29939 => 8779,
    29940 => 8776,
    29941 => 8773,
    29942 => 8770,
    29943 => 8767,
    29944 => 8764,
    29945 => 8761,
    29946 => 8758,
    29947 => 8755,
    29948 => 8751,
    29949 => 8748,
    29950 => 8745,
    29951 => 8742,
    29952 => 8739,
    29953 => 8736,
    29954 => 8733,
    29955 => 8730,
    29956 => 8727,
    29957 => 8724,
    29958 => 8721,
    29959 => 8718,
    29960 => 8715,
    29961 => 8712,
    29962 => 8709,
    29963 => 8706,
    29964 => 8703,
    29965 => 8700,
    29966 => 8697,
    29967 => 8694,
    29968 => 8691,
    29969 => 8688,
    29970 => 8685,
    29971 => 8682,
    29972 => 8679,
    29973 => 8676,
    29974 => 8673,
    29975 => 8670,
    29976 => 8667,
    29977 => 8664,
    29978 => 8661,
    29979 => 8658,
    29980 => 8655,
    29981 => 8652,
    29982 => 8649,
    29983 => 8645,
    29984 => 8642,
    29985 => 8639,
    29986 => 8636,
    29987 => 8633,
    29988 => 8630,
    29989 => 8627,
    29990 => 8624,
    29991 => 8621,
    29992 => 8618,
    29993 => 8615,
    29994 => 8612,
    29995 => 8609,
    29996 => 8606,
    29997 => 8603,
    29998 => 8600,
    29999 => 8597,
    30000 => 8594,
    30001 => 8591,
    30002 => 8588,
    30003 => 8585,
    30004 => 8582,
    30005 => 8579,
    30006 => 8576,
    30007 => 8573,
    30008 => 8570,
    30009 => 8567,
    30010 => 8564,
    30011 => 8561,
    30012 => 8558,
    30013 => 8555,
    30014 => 8552,
    30015 => 8548,
    30016 => 8545,
    30017 => 8542,
    30018 => 8539,
    30019 => 8536,
    30020 => 8533,
    30021 => 8530,
    30022 => 8527,
    30023 => 8524,
    30024 => 8521,
    30025 => 8518,
    30026 => 8515,
    30027 => 8512,
    30028 => 8509,
    30029 => 8506,
    30030 => 8503,
    30031 => 8500,
    30032 => 8497,
    30033 => 8494,
    30034 => 8491,
    30035 => 8488,
    30036 => 8485,
    30037 => 8482,
    30038 => 8479,
    30039 => 8476,
    30040 => 8473,
    30041 => 8470,
    30042 => 8467,
    30043 => 8464,
    30044 => 8460,
    30045 => 8457,
    30046 => 8454,
    30047 => 8451,
    30048 => 8448,
    30049 => 8445,
    30050 => 8442,
    30051 => 8439,
    30052 => 8436,
    30053 => 8433,
    30054 => 8430,
    30055 => 8427,
    30056 => 8424,
    30057 => 8421,
    30058 => 8418,
    30059 => 8415,
    30060 => 8412,
    30061 => 8409,
    30062 => 8406,
    30063 => 8403,
    30064 => 8400,
    30065 => 8397,
    30066 => 8394,
    30067 => 8391,
    30068 => 8388,
    30069 => 8385,
    30070 => 8382,
    30071 => 8379,
    30072 => 8375,
    30073 => 8372,
    30074 => 8369,
    30075 => 8366,
    30076 => 8363,
    30077 => 8360,
    30078 => 8357,
    30079 => 8354,
    30080 => 8351,
    30081 => 8348,
    30082 => 8345,
    30083 => 8342,
    30084 => 8339,
    30085 => 8336,
    30086 => 8333,
    30087 => 8330,
    30088 => 8327,
    30089 => 8324,
    30090 => 8321,
    30091 => 8318,
    30092 => 8315,
    30093 => 8312,
    30094 => 8309,
    30095 => 8306,
    30096 => 8303,
    30097 => 8300,
    30098 => 8296,
    30099 => 8293,
    30100 => 8290,
    30101 => 8287,
    30102 => 8284,
    30103 => 8281,
    30104 => 8278,
    30105 => 8275,
    30106 => 8272,
    30107 => 8269,
    30108 => 8266,
    30109 => 8263,
    30110 => 8260,
    30111 => 8257,
    30112 => 8254,
    30113 => 8251,
    30114 => 8248,
    30115 => 8245,
    30116 => 8242,
    30117 => 8239,
    30118 => 8236,
    30119 => 8233,
    30120 => 8230,
    30121 => 8227,
    30122 => 8224,
    30123 => 8220,
    30124 => 8217,
    30125 => 8214,
    30126 => 8211,
    30127 => 8208,
    30128 => 8205,
    30129 => 8202,
    30130 => 8199,
    30131 => 8196,
    30132 => 8193,
    30133 => 8190,
    30134 => 8187,
    30135 => 8184,
    30136 => 8181,
    30137 => 8178,
    30138 => 8175,
    30139 => 8172,
    30140 => 8169,
    30141 => 8166,
    30142 => 8163,
    30143 => 8160,
    30144 => 8157,
    30145 => 8154,
    30146 => 8151,
    30147 => 8147,
    30148 => 8144,
    30149 => 8141,
    30150 => 8138,
    30151 => 8135,
    30152 => 8132,
    30153 => 8129,
    30154 => 8126,
    30155 => 8123,
    30156 => 8120,
    30157 => 8117,
    30158 => 8114,
    30159 => 8111,
    30160 => 8108,
    30161 => 8105,
    30162 => 8102,
    30163 => 8099,
    30164 => 8096,
    30165 => 8093,
    30166 => 8090,
    30167 => 8087,
    30168 => 8084,
    30169 => 8081,
    30170 => 8077,
    30171 => 8074,
    30172 => 8071,
    30173 => 8068,
    30174 => 8065,
    30175 => 8062,
    30176 => 8059,
    30177 => 8056,
    30178 => 8053,
    30179 => 8050,
    30180 => 8047,
    30181 => 8044,
    30182 => 8041,
    30183 => 8038,
    30184 => 8035,
    30185 => 8032,
    30186 => 8029,
    30187 => 8026,
    30188 => 8023,
    30189 => 8020,
    30190 => 8017,
    30191 => 8014,
    30192 => 8010,
    30193 => 8007,
    30194 => 8004,
    30195 => 8001,
    30196 => 7998,
    30197 => 7995,
    30198 => 7992,
    30199 => 7989,
    30200 => 7986,
    30201 => 7983,
    30202 => 7980,
    30203 => 7977,
    30204 => 7974,
    30205 => 7971,
    30206 => 7968,
    30207 => 7965,
    30208 => 7962,
    30209 => 7959,
    30210 => 7956,
    30211 => 7953,
    30212 => 7950,
    30213 => 7946,
    30214 => 7943,
    30215 => 7940,
    30216 => 7937,
    30217 => 7934,
    30218 => 7931,
    30219 => 7928,
    30220 => 7925,
    30221 => 7922,
    30222 => 7919,
    30223 => 7916,
    30224 => 7913,
    30225 => 7910,
    30226 => 7907,
    30227 => 7904,
    30228 => 7901,
    30229 => 7898,
    30230 => 7895,
    30231 => 7892,
    30232 => 7889,
    30233 => 7886,
    30234 => 7882,
    30235 => 7879,
    30236 => 7876,
    30237 => 7873,
    30238 => 7870,
    30239 => 7867,
    30240 => 7864,
    30241 => 7861,
    30242 => 7858,
    30243 => 7855,
    30244 => 7852,
    30245 => 7849,
    30246 => 7846,
    30247 => 7843,
    30248 => 7840,
    30249 => 7837,
    30250 => 7834,
    30251 => 7831,
    30252 => 7828,
    30253 => 7825,
    30254 => 7821,
    30255 => 7818,
    30256 => 7815,
    30257 => 7812,
    30258 => 7809,
    30259 => 7806,
    30260 => 7803,
    30261 => 7800,
    30262 => 7797,
    30263 => 7794,
    30264 => 7791,
    30265 => 7788,
    30266 => 7785,
    30267 => 7782,
    30268 => 7779,
    30269 => 7776,
    30270 => 7773,
    30271 => 7770,
    30272 => 7767,
    30273 => 7764,
    30274 => 7760,
    30275 => 7757,
    30276 => 7754,
    30277 => 7751,
    30278 => 7748,
    30279 => 7745,
    30280 => 7742,
    30281 => 7739,
    30282 => 7736,
    30283 => 7733,
    30284 => 7730,
    30285 => 7727,
    30286 => 7724,
    30287 => 7721,
    30288 => 7718,
    30289 => 7715,
    30290 => 7712,
    30291 => 7709,
    30292 => 7705,
    30293 => 7702,
    30294 => 7699,
    30295 => 7696,
    30296 => 7693,
    30297 => 7690,
    30298 => 7687,
    30299 => 7684,
    30300 => 7681,
    30301 => 7678,
    30302 => 7675,
    30303 => 7672,
    30304 => 7669,
    30305 => 7666,
    30306 => 7663,
    30307 => 7660,
    30308 => 7657,
    30309 => 7654,
    30310 => 7651,
    30311 => 7647,
    30312 => 7644,
    30313 => 7641,
    30314 => 7638,
    30315 => 7635,
    30316 => 7632,
    30317 => 7629,
    30318 => 7626,
    30319 => 7623,
    30320 => 7620,
    30321 => 7617,
    30322 => 7614,
    30323 => 7611,
    30324 => 7608,
    30325 => 7605,
    30326 => 7602,
    30327 => 7599,
    30328 => 7596,
    30329 => 7592,
    30330 => 7589,
    30331 => 7586,
    30332 => 7583,
    30333 => 7580,
    30334 => 7577,
    30335 => 7574,
    30336 => 7571,
    30337 => 7568,
    30338 => 7565,
    30339 => 7562,
    30340 => 7559,
    30341 => 7556,
    30342 => 7553,
    30343 => 7550,
    30344 => 7547,
    30345 => 7544,
    30346 => 7541,
    30347 => 7537,
    30348 => 7534,
    30349 => 7531,
    30350 => 7528,
    30351 => 7525,
    30352 => 7522,
    30353 => 7519,
    30354 => 7516,
    30355 => 7513,
    30356 => 7510,
    30357 => 7507,
    30358 => 7504,
    30359 => 7501,
    30360 => 7498,
    30361 => 7495,
    30362 => 7492,
    30363 => 7489,
    30364 => 7485,
    30365 => 7482,
    30366 => 7479,
    30367 => 7476,
    30368 => 7473,
    30369 => 7470,
    30370 => 7467,
    30371 => 7464,
    30372 => 7461,
    30373 => 7458,
    30374 => 7455,
    30375 => 7452,
    30376 => 7449,
    30377 => 7446,
    30378 => 7443,
    30379 => 7440,
    30380 => 7437,
    30381 => 7433,
    30382 => 7430,
    30383 => 7427,
    30384 => 7424,
    30385 => 7421,
    30386 => 7418,
    30387 => 7415,
    30388 => 7412,
    30389 => 7409,
    30390 => 7406,
    30391 => 7403,
    30392 => 7400,
    30393 => 7397,
    30394 => 7394,
    30395 => 7391,
    30396 => 7388,
    30397 => 7385,
    30398 => 7381,
    30399 => 7378,
    30400 => 7375,
    30401 => 7372,
    30402 => 7369,
    30403 => 7366,
    30404 => 7363,
    30405 => 7360,
    30406 => 7357,
    30407 => 7354,
    30408 => 7351,
    30409 => 7348,
    30410 => 7345,
    30411 => 7342,
    30412 => 7339,
    30413 => 7336,
    30414 => 7332,
    30415 => 7329,
    30416 => 7326,
    30417 => 7323,
    30418 => 7320,
    30419 => 7317,
    30420 => 7314,
    30421 => 7311,
    30422 => 7308,
    30423 => 7305,
    30424 => 7302,
    30425 => 7299,
    30426 => 7296,
    30427 => 7293,
    30428 => 7290,
    30429 => 7287,
    30430 => 7283,
    30431 => 7280,
    30432 => 7277,
    30433 => 7274,
    30434 => 7271,
    30435 => 7268,
    30436 => 7265,
    30437 => 7262,
    30438 => 7259,
    30439 => 7256,
    30440 => 7253,
    30441 => 7250,
    30442 => 7247,
    30443 => 7244,
    30444 => 7241,
    30445 => 7238,
    30446 => 7234,
    30447 => 7231,
    30448 => 7228,
    30449 => 7225,
    30450 => 7222,
    30451 => 7219,
    30452 => 7216,
    30453 => 7213,
    30454 => 7210,
    30455 => 7207,
    30456 => 7204,
    30457 => 7201,
    30458 => 7198,
    30459 => 7195,
    30460 => 7192,
    30461 => 7188,
    30462 => 7185,
    30463 => 7182,
    30464 => 7179,
    30465 => 7176,
    30466 => 7173,
    30467 => 7170,
    30468 => 7167,
    30469 => 7164,
    30470 => 7161,
    30471 => 7158,
    30472 => 7155,
    30473 => 7152,
    30474 => 7149,
    30475 => 7146,
    30476 => 7143,
    30477 => 7139,
    30478 => 7136,
    30479 => 7133,
    30480 => 7130,
    30481 => 7127,
    30482 => 7124,
    30483 => 7121,
    30484 => 7118,
    30485 => 7115,
    30486 => 7112,
    30487 => 7109,
    30488 => 7106,
    30489 => 7103,
    30490 => 7100,
    30491 => 7097,
    30492 => 7093,
    30493 => 7090,
    30494 => 7087,
    30495 => 7084,
    30496 => 7081,
    30497 => 7078,
    30498 => 7075,
    30499 => 7072,
    30500 => 7069,
    30501 => 7066,
    30502 => 7063,
    30503 => 7060,
    30504 => 7057,
    30505 => 7054,
    30506 => 7050,
    30507 => 7047,
    30508 => 7044,
    30509 => 7041,
    30510 => 7038,
    30511 => 7035,
    30512 => 7032,
    30513 => 7029,
    30514 => 7026,
    30515 => 7023,
    30516 => 7020,
    30517 => 7017,
    30518 => 7014,
    30519 => 7011,
    30520 => 7008,
    30521 => 7004,
    30522 => 7001,
    30523 => 6998,
    30524 => 6995,
    30525 => 6992,
    30526 => 6989,
    30527 => 6986,
    30528 => 6983,
    30529 => 6980,
    30530 => 6977,
    30531 => 6974,
    30532 => 6971,
    30533 => 6968,
    30534 => 6965,
    30535 => 6961,
    30536 => 6958,
    30537 => 6955,
    30538 => 6952,
    30539 => 6949,
    30540 => 6946,
    30541 => 6943,
    30542 => 6940,
    30543 => 6937,
    30544 => 6934,
    30545 => 6931,
    30546 => 6928,
    30547 => 6925,
    30548 => 6922,
    30549 => 6919,
    30550 => 6915,
    30551 => 6912,
    30552 => 6909,
    30553 => 6906,
    30554 => 6903,
    30555 => 6900,
    30556 => 6897,
    30557 => 6894,
    30558 => 6891,
    30559 => 6888,
    30560 => 6885,
    30561 => 6882,
    30562 => 6879,
    30563 => 6876,
    30564 => 6872,
    30565 => 6869,
    30566 => 6866,
    30567 => 6863,
    30568 => 6860,
    30569 => 6857,
    30570 => 6854,
    30571 => 6851,
    30572 => 6848,
    30573 => 6845,
    30574 => 6842,
    30575 => 6839,
    30576 => 6836,
    30577 => 6833,
    30578 => 6829,
    30579 => 6826,
    30580 => 6823,
    30581 => 6820,
    30582 => 6817,
    30583 => 6814,
    30584 => 6811,
    30585 => 6808,
    30586 => 6805,
    30587 => 6802,
    30588 => 6799,
    30589 => 6796,
    30590 => 6793,
    30591 => 6789,
    30592 => 6786,
    30593 => 6783,
    30594 => 6780,
    30595 => 6777,
    30596 => 6774,
    30597 => 6771,
    30598 => 6768,
    30599 => 6765,
    30600 => 6762,
    30601 => 6759,
    30602 => 6756,
    30603 => 6753,
    30604 => 6750,
    30605 => 6746,
    30606 => 6743,
    30607 => 6740,
    30608 => 6737,
    30609 => 6734,
    30610 => 6731,
    30611 => 6728,
    30612 => 6725,
    30613 => 6722,
    30614 => 6719,
    30615 => 6716,
    30616 => 6713,
    30617 => 6710,
    30618 => 6706,
    30619 => 6703,
    30620 => 6700,
    30621 => 6697,
    30622 => 6694,
    30623 => 6691,
    30624 => 6688,
    30625 => 6685,
    30626 => 6682,
    30627 => 6679,
    30628 => 6676,
    30629 => 6673,
    30630 => 6670,
    30631 => 6667,
    30632 => 6663,
    30633 => 6660,
    30634 => 6657,
    30635 => 6654,
    30636 => 6651,
    30637 => 6648,
    30638 => 6645,
    30639 => 6642,
    30640 => 6639,
    30641 => 6636,
    30642 => 6633,
    30643 => 6630,
    30644 => 6627,
    30645 => 6623,
    30646 => 6620,
    30647 => 6617,
    30648 => 6614,
    30649 => 6611,
    30650 => 6608,
    30651 => 6605,
    30652 => 6602,
    30653 => 6599,
    30654 => 6596,
    30655 => 6593,
    30656 => 6590,
    30657 => 6587,
    30658 => 6583,
    30659 => 6580,
    30660 => 6577,
    30661 => 6574,
    30662 => 6571,
    30663 => 6568,
    30664 => 6565,
    30665 => 6562,
    30666 => 6559,
    30667 => 6556,
    30668 => 6553,
    30669 => 6550,
    30670 => 6547,
    30671 => 6543,
    30672 => 6540,
    30673 => 6537,
    30674 => 6534,
    30675 => 6531,
    30676 => 6528,
    30677 => 6525,
    30678 => 6522,
    30679 => 6519,
    30680 => 6516,
    30681 => 6513,
    30682 => 6510,
    30683 => 6506,
    30684 => 6503,
    30685 => 6500,
    30686 => 6497,
    30687 => 6494,
    30688 => 6491,
    30689 => 6488,
    30690 => 6485,
    30691 => 6482,
    30692 => 6479,
    30693 => 6476,
    30694 => 6473,
    30695 => 6470,
    30696 => 6466,
    30697 => 6463,
    30698 => 6460,
    30699 => 6457,
    30700 => 6454,
    30701 => 6451,
    30702 => 6448,
    30703 => 6445,
    30704 => 6442,
    30705 => 6439,
    30706 => 6436,
    30707 => 6433,
    30708 => 6429,
    30709 => 6426,
    30710 => 6423,
    30711 => 6420,
    30712 => 6417,
    30713 => 6414,
    30714 => 6411,
    30715 => 6408,
    30716 => 6405,
    30717 => 6402,
    30718 => 6399,
    30719 => 6396,
    30720 => 6393,
    30721 => 6389,
    30722 => 6386,
    30723 => 6383,
    30724 => 6380,
    30725 => 6377,
    30726 => 6374,
    30727 => 6371,
    30728 => 6368,
    30729 => 6365,
    30730 => 6362,
    30731 => 6359,
    30732 => 6356,
    30733 => 6352,
    30734 => 6349,
    30735 => 6346,
    30736 => 6343,
    30737 => 6340,
    30738 => 6337,
    30739 => 6334,
    30740 => 6331,
    30741 => 6328,
    30742 => 6325,
    30743 => 6322,
    30744 => 6319,
    30745 => 6315,
    30746 => 6312,
    30747 => 6309,
    30748 => 6306,
    30749 => 6303,
    30750 => 6300,
    30751 => 6297,
    30752 => 6294,
    30753 => 6291,
    30754 => 6288,
    30755 => 6285,
    30756 => 6282,
    30757 => 6278,
    30758 => 6275,
    30759 => 6272,
    30760 => 6269,
    30761 => 6266,
    30762 => 6263,
    30763 => 6260,
    30764 => 6257,
    30765 => 6254,
    30766 => 6251,
    30767 => 6248,
    30768 => 6245,
    30769 => 6241,
    30770 => 6238,
    30771 => 6235,
    30772 => 6232,
    30773 => 6229,
    30774 => 6226,
    30775 => 6223,
    30776 => 6220,
    30777 => 6217,
    30778 => 6214,
    30779 => 6211,
    30780 => 6208,
    30781 => 6204,
    30782 => 6201,
    30783 => 6198,
    30784 => 6195,
    30785 => 6192,
    30786 => 6189,
    30787 => 6186,
    30788 => 6183,
    30789 => 6180,
    30790 => 6177,
    30791 => 6174,
    30792 => 6171,
    30793 => 6167,
    30794 => 6164,
    30795 => 6161,
    30796 => 6158,
    30797 => 6155,
    30798 => 6152,
    30799 => 6149,
    30800 => 6146,
    30801 => 6143,
    30802 => 6140,
    30803 => 6137,
    30804 => 6134,
    30805 => 6130,
    30806 => 6127,
    30807 => 6124,
    30808 => 6121,
    30809 => 6118,
    30810 => 6115,
    30811 => 6112,
    30812 => 6109,
    30813 => 6106,
    30814 => 6103,
    30815 => 6100,
    30816 => 6096,
    30817 => 6093,
    30818 => 6090,
    30819 => 6087,
    30820 => 6084,
    30821 => 6081,
    30822 => 6078,
    30823 => 6075,
    30824 => 6072,
    30825 => 6069,
    30826 => 6066,
    30827 => 6063,
    30828 => 6059,
    30829 => 6056,
    30830 => 6053,
    30831 => 6050,
    30832 => 6047,
    30833 => 6044,
    30834 => 6041,
    30835 => 6038,
    30836 => 6035,
    30837 => 6032,
    30838 => 6029,
    30839 => 6025,
    30840 => 6022,
    30841 => 6019,
    30842 => 6016,
    30843 => 6013,
    30844 => 6010,
    30845 => 6007,
    30846 => 6004,
    30847 => 6001,
    30848 => 5998,
    30849 => 5995,
    30850 => 5991,
    30851 => 5988,
    30852 => 5985,
    30853 => 5982,
    30854 => 5979,
    30855 => 5976,
    30856 => 5973,
    30857 => 5970,
    30858 => 5967,
    30859 => 5964,
    30860 => 5961,
    30861 => 5958,
    30862 => 5954,
    30863 => 5951,
    30864 => 5948,
    30865 => 5945,
    30866 => 5942,
    30867 => 5939,
    30868 => 5936,
    30869 => 5933,
    30870 => 5930,
    30871 => 5927,
    30872 => 5924,
    30873 => 5920,
    30874 => 5917,
    30875 => 5914,
    30876 => 5911,
    30877 => 5908,
    30878 => 5905,
    30879 => 5902,
    30880 => 5899,
    30881 => 5896,
    30882 => 5893,
    30883 => 5890,
    30884 => 5886,
    30885 => 5883,
    30886 => 5880,
    30887 => 5877,
    30888 => 5874,
    30889 => 5871,
    30890 => 5868,
    30891 => 5865,
    30892 => 5862,
    30893 => 5859,
    30894 => 5856,
    30895 => 5852,
    30896 => 5849,
    30897 => 5846,
    30898 => 5843,
    30899 => 5840,
    30900 => 5837,
    30901 => 5834,
    30902 => 5831,
    30903 => 5828,
    30904 => 5825,
    30905 => 5822,
    30906 => 5818,
    30907 => 5815,
    30908 => 5812,
    30909 => 5809,
    30910 => 5806,
    30911 => 5803,
    30912 => 5800,
    30913 => 5797,
    30914 => 5794,
    30915 => 5791,
    30916 => 5788,
    30917 => 5784,
    30918 => 5781,
    30919 => 5778,
    30920 => 5775,
    30921 => 5772,
    30922 => 5769,
    30923 => 5766,
    30924 => 5763,
    30925 => 5760,
    30926 => 5757,
    30927 => 5754,
    30928 => 5750,
    30929 => 5747,
    30930 => 5744,
    30931 => 5741,
    30932 => 5738,
    30933 => 5735,
    30934 => 5732,
    30935 => 5729,
    30936 => 5726,
    30937 => 5723,
    30938 => 5719,
    30939 => 5716,
    30940 => 5713,
    30941 => 5710,
    30942 => 5707,
    30943 => 5704,
    30944 => 5701,
    30945 => 5698,
    30946 => 5695,
    30947 => 5692,
    30948 => 5689,
    30949 => 5685,
    30950 => 5682,
    30951 => 5679,
    30952 => 5676,
    30953 => 5673,
    30954 => 5670,
    30955 => 5667,
    30956 => 5664,
    30957 => 5661,
    30958 => 5658,
    30959 => 5655,
    30960 => 5651,
    30961 => 5648,
    30962 => 5645,
    30963 => 5642,
    30964 => 5639,
    30965 => 5636,
    30966 => 5633,
    30967 => 5630,
    30968 => 5627,
    30969 => 5624,
    30970 => 5620,
    30971 => 5617,
    30972 => 5614,
    30973 => 5611,
    30974 => 5608,
    30975 => 5605,
    30976 => 5602,
    30977 => 5599,
    30978 => 5596,
    30979 => 5593,
    30980 => 5590,
    30981 => 5586,
    30982 => 5583,
    30983 => 5580,
    30984 => 5577,
    30985 => 5574,
    30986 => 5571,
    30987 => 5568,
    30988 => 5565,
    30989 => 5562,
    30990 => 5559,
    30991 => 5555,
    30992 => 5552,
    30993 => 5549,
    30994 => 5546,
    30995 => 5543,
    30996 => 5540,
    30997 => 5537,
    30998 => 5534,
    30999 => 5531,
    31000 => 5528,
    31001 => 5525,
    31002 => 5521,
    31003 => 5518,
    31004 => 5515,
    31005 => 5512,
    31006 => 5509,
    31007 => 5506,
    31008 => 5503,
    31009 => 5500,
    31010 => 5497,
    31011 => 5494,
    31012 => 5490,
    31013 => 5487,
    31014 => 5484,
    31015 => 5481,
    31016 => 5478,
    31017 => 5475,
    31018 => 5472,
    31019 => 5469,
    31020 => 5466,
    31021 => 5463,
    31022 => 5459,
    31023 => 5456,
    31024 => 5453,
    31025 => 5450,
    31026 => 5447,
    31027 => 5444,
    31028 => 5441,
    31029 => 5438,
    31030 => 5435,
    31031 => 5432,
    31032 => 5428,
    31033 => 5425,
    31034 => 5422,
    31035 => 5419,
    31036 => 5416,
    31037 => 5413,
    31038 => 5410,
    31039 => 5407,
    31040 => 5404,
    31041 => 5401,
    31042 => 5398,
    31043 => 5394,
    31044 => 5391,
    31045 => 5388,
    31046 => 5385,
    31047 => 5382,
    31048 => 5379,
    31049 => 5376,
    31050 => 5373,
    31051 => 5370,
    31052 => 5367,
    31053 => 5363,
    31054 => 5360,
    31055 => 5357,
    31056 => 5354,
    31057 => 5351,
    31058 => 5348,
    31059 => 5345,
    31060 => 5342,
    31061 => 5339,
    31062 => 5336,
    31063 => 5332,
    31064 => 5329,
    31065 => 5326,
    31066 => 5323,
    31067 => 5320,
    31068 => 5317,
    31069 => 5314,
    31070 => 5311,
    31071 => 5308,
    31072 => 5305,
    31073 => 5301,
    31074 => 5298,
    31075 => 5295,
    31076 => 5292,
    31077 => 5289,
    31078 => 5286,
    31079 => 5283,
    31080 => 5280,
    31081 => 5277,
    31082 => 5274,
    31083 => 5270,
    31084 => 5267,
    31085 => 5264,
    31086 => 5261,
    31087 => 5258,
    31088 => 5255,
    31089 => 5252,
    31090 => 5249,
    31091 => 5246,
    31092 => 5243,
    31093 => 5239,
    31094 => 5236,
    31095 => 5233,
    31096 => 5230,
    31097 => 5227,
    31098 => 5224,
    31099 => 5221,
    31100 => 5218,
    31101 => 5215,
    31102 => 5212,
    31103 => 5208,
    31104 => 5205,
    31105 => 5202,
    31106 => 5199,
    31107 => 5196,
    31108 => 5193,
    31109 => 5190,
    31110 => 5187,
    31111 => 5184,
    31112 => 5180,
    31113 => 5177,
    31114 => 5174,
    31115 => 5171,
    31116 => 5168,
    31117 => 5165,
    31118 => 5162,
    31119 => 5159,
    31120 => 5156,
    31121 => 5153,
    31122 => 5149,
    31123 => 5146,
    31124 => 5143,
    31125 => 5140,
    31126 => 5137,
    31127 => 5134,
    31128 => 5131,
    31129 => 5128,
    31130 => 5125,
    31131 => 5122,
    31132 => 5118,
    31133 => 5115,
    31134 => 5112,
    31135 => 5109,
    31136 => 5106,
    31137 => 5103,
    31138 => 5100,
    31139 => 5097,
    31140 => 5094,
    31141 => 5091,
    31142 => 5087,
    31143 => 5084,
    31144 => 5081,
    31145 => 5078,
    31146 => 5075,
    31147 => 5072,
    31148 => 5069,
    31149 => 5066,
    31150 => 5063,
    31151 => 5059,
    31152 => 5056,
    31153 => 5053,
    31154 => 5050,
    31155 => 5047,
    31156 => 5044,
    31157 => 5041,
    31158 => 5038,
    31159 => 5035,
    31160 => 5032,
    31161 => 5028,
    31162 => 5025,
    31163 => 5022,
    31164 => 5019,
    31165 => 5016,
    31166 => 5013,
    31167 => 5010,
    31168 => 5007,
    31169 => 5004,
    31170 => 5000,
    31171 => 4997,
    31172 => 4994,
    31173 => 4991,
    31174 => 4988,
    31175 => 4985,
    31176 => 4982,
    31177 => 4979,
    31178 => 4976,
    31179 => 4973,
    31180 => 4969,
    31181 => 4966,
    31182 => 4963,
    31183 => 4960,
    31184 => 4957,
    31185 => 4954,
    31186 => 4951,
    31187 => 4948,
    31188 => 4945,
    31189 => 4941,
    31190 => 4938,
    31191 => 4935,
    31192 => 4932,
    31193 => 4929,
    31194 => 4926,
    31195 => 4923,
    31196 => 4920,
    31197 => 4917,
    31198 => 4914,
    31199 => 4910,
    31200 => 4907,
    31201 => 4904,
    31202 => 4901,
    31203 => 4898,
    31204 => 4895,
    31205 => 4892,
    31206 => 4889,
    31207 => 4886,
    31208 => 4882,
    31209 => 4879,
    31210 => 4876,
    31211 => 4873,
    31212 => 4870,
    31213 => 4867,
    31214 => 4864,
    31215 => 4861,
    31216 => 4858,
    31217 => 4855,
    31218 => 4851,
    31219 => 4848,
    31220 => 4845,
    31221 => 4842,
    31222 => 4839,
    31223 => 4836,
    31224 => 4833,
    31225 => 4830,
    31226 => 4827,
    31227 => 4823,
    31228 => 4820,
    31229 => 4817,
    31230 => 4814,
    31231 => 4811,
    31232 => 4808,
    31233 => 4805,
    31234 => 4802,
    31235 => 4799,
    31236 => 4795,
    31237 => 4792,
    31238 => 4789,
    31239 => 4786,
    31240 => 4783,
    31241 => 4780,
    31242 => 4777,
    31243 => 4774,
    31244 => 4771,
    31245 => 4768,
    31246 => 4764,
    31247 => 4761,
    31248 => 4758,
    31249 => 4755,
    31250 => 4752,
    31251 => 4749,
    31252 => 4746,
    31253 => 4743,
    31254 => 4740,
    31255 => 4736,
    31256 => 4733,
    31257 => 4730,
    31258 => 4727,
    31259 => 4724,
    31260 => 4721,
    31261 => 4718,
    31262 => 4715,
    31263 => 4712,
    31264 => 4708,
    31265 => 4705,
    31266 => 4702,
    31267 => 4699,
    31268 => 4696,
    31269 => 4693,
    31270 => 4690,
    31271 => 4687,
    31272 => 4684,
    31273 => 4680,
    31274 => 4677,
    31275 => 4674,
    31276 => 4671,
    31277 => 4668,
    31278 => 4665,
    31279 => 4662,
    31280 => 4659,
    31281 => 4656,
    31282 => 4652,
    31283 => 4649,
    31284 => 4646,
    31285 => 4643,
    31286 => 4640,
    31287 => 4637,
    31288 => 4634,
    31289 => 4631,
    31290 => 4628,
    31291 => 4624,
    31292 => 4621,
    31293 => 4618,
    31294 => 4615,
    31295 => 4612,
    31296 => 4609,
    31297 => 4606,
    31298 => 4603,
    31299 => 4600,
    31300 => 4597,
    31301 => 4593,
    31302 => 4590,
    31303 => 4587,
    31304 => 4584,
    31305 => 4581,
    31306 => 4578,
    31307 => 4575,
    31308 => 4572,
    31309 => 4569,
    31310 => 4565,
    31311 => 4562,
    31312 => 4559,
    31313 => 4556,
    31314 => 4553,
    31315 => 4550,
    31316 => 4547,
    31317 => 4544,
    31318 => 4541,
    31319 => 4537,
    31320 => 4534,
    31321 => 4531,
    31322 => 4528,
    31323 => 4525,
    31324 => 4522,
    31325 => 4519,
    31326 => 4516,
    31327 => 4513,
    31328 => 4509,
    31329 => 4506,
    31330 => 4503,
    31331 => 4500,
    31332 => 4497,
    31333 => 4494,
    31334 => 4491,
    31335 => 4488,
    31336 => 4485,
    31337 => 4481,
    31338 => 4478,
    31339 => 4475,
    31340 => 4472,
    31341 => 4469,
    31342 => 4466,
    31343 => 4463,
    31344 => 4460,
    31345 => 4456,
    31346 => 4453,
    31347 => 4450,
    31348 => 4447,
    31349 => 4444,
    31350 => 4441,
    31351 => 4438,
    31352 => 4435,
    31353 => 4432,
    31354 => 4428,
    31355 => 4425,
    31356 => 4422,
    31357 => 4419,
    31358 => 4416,
    31359 => 4413,
    31360 => 4410,
    31361 => 4407,
    31362 => 4404,
    31363 => 4400,
    31364 => 4397,
    31365 => 4394,
    31366 => 4391,
    31367 => 4388,
    31368 => 4385,
    31369 => 4382,
    31370 => 4379,
    31371 => 4376,
    31372 => 4372,
    31373 => 4369,
    31374 => 4366,
    31375 => 4363,
    31376 => 4360,
    31377 => 4357,
    31378 => 4354,
    31379 => 4351,
    31380 => 4348,
    31381 => 4344,
    31382 => 4341,
    31383 => 4338,
    31384 => 4335,
    31385 => 4332,
    31386 => 4329,
    31387 => 4326,
    31388 => 4323,
    31389 => 4320,
    31390 => 4316,
    31391 => 4313,
    31392 => 4310,
    31393 => 4307,
    31394 => 4304,
    31395 => 4301,
    31396 => 4298,
    31397 => 4295,
    31398 => 4291,
    31399 => 4288,
    31400 => 4285,
    31401 => 4282,
    31402 => 4279,
    31403 => 4276,
    31404 => 4273,
    31405 => 4270,
    31406 => 4267,
    31407 => 4263,
    31408 => 4260,
    31409 => 4257,
    31410 => 4254,
    31411 => 4251,
    31412 => 4248,
    31413 => 4245,
    31414 => 4242,
    31415 => 4239,
    31416 => 4235,
    31417 => 4232,
    31418 => 4229,
    31419 => 4226,
    31420 => 4223,
    31421 => 4220,
    31422 => 4217,
    31423 => 4214,
    31424 => 4210,
    31425 => 4207,
    31426 => 4204,
    31427 => 4201,
    31428 => 4198,
    31429 => 4195,
    31430 => 4192,
    31431 => 4189,
    31432 => 4186,
    31433 => 4182,
    31434 => 4179,
    31435 => 4176,
    31436 => 4173,
    31437 => 4170,
    31438 => 4167,
    31439 => 4164,
    31440 => 4161,
    31441 => 4158,
    31442 => 4154,
    31443 => 4151,
    31444 => 4148,
    31445 => 4145,
    31446 => 4142,
    31447 => 4139,
    31448 => 4136,
    31449 => 4133,
    31450 => 4129,
    31451 => 4126,
    31452 => 4123,
    31453 => 4120,
    31454 => 4117,
    31455 => 4114,
    31456 => 4111,
    31457 => 4108,
    31458 => 4105,
    31459 => 4101,
    31460 => 4098,
    31461 => 4095,
    31462 => 4092,
    31463 => 4089,
    31464 => 4086,
    31465 => 4083,
    31466 => 4080,
    31467 => 4076,
    31468 => 4073,
    31469 => 4070,
    31470 => 4067,
    31471 => 4064,
    31472 => 4061,
    31473 => 4058,
    31474 => 4055,
    31475 => 4052,
    31476 => 4048,
    31477 => 4045,
    31478 => 4042,
    31479 => 4039,
    31480 => 4036,
    31481 => 4033,
    31482 => 4030,
    31483 => 4027,
    31484 => 4024,
    31485 => 4020,
    31486 => 4017,
    31487 => 4014,
    31488 => 4011,
    31489 => 4008,
    31490 => 4005,
    31491 => 4002,
    31492 => 3999,
    31493 => 3995,
    31494 => 3992,
    31495 => 3989,
    31496 => 3986,
    31497 => 3983,
    31498 => 3980,
    31499 => 3977,
    31500 => 3974,
    31501 => 3970,
    31502 => 3967,
    31503 => 3964,
    31504 => 3961,
    31505 => 3958,
    31506 => 3955,
    31507 => 3952,
    31508 => 3949,
    31509 => 3946,
    31510 => 3942,
    31511 => 3939,
    31512 => 3936,
    31513 => 3933,
    31514 => 3930,
    31515 => 3927,
    31516 => 3924,
    31517 => 3921,
    31518 => 3917,
    31519 => 3914,
    31520 => 3911,
    31521 => 3908,
    31522 => 3905,
    31523 => 3902,
    31524 => 3899,
    31525 => 3896,
    31526 => 3893,
    31527 => 3889,
    31528 => 3886,
    31529 => 3883,
    31530 => 3880,
    31531 => 3877,
    31532 => 3874,
    31533 => 3871,
    31534 => 3868,
    31535 => 3864,
    31536 => 3861,
    31537 => 3858,
    31538 => 3855,
    31539 => 3852,
    31540 => 3849,
    31541 => 3846,
    31542 => 3843,
    31543 => 3839,
    31544 => 3836,
    31545 => 3833,
    31546 => 3830,
    31547 => 3827,
    31548 => 3824,
    31549 => 3821,
    31550 => 3818,
    31551 => 3815,
    31552 => 3811,
    31553 => 3808,
    31554 => 3805,
    31555 => 3802,
    31556 => 3799,
    31557 => 3796,
    31558 => 3793,
    31559 => 3790,
    31560 => 3786,
    31561 => 3783,
    31562 => 3780,
    31563 => 3777,
    31564 => 3774,
    31565 => 3771,
    31566 => 3768,
    31567 => 3765,
    31568 => 3761,
    31569 => 3758,
    31570 => 3755,
    31571 => 3752,
    31572 => 3749,
    31573 => 3746,
    31574 => 3743,
    31575 => 3740,
    31576 => 3737,
    31577 => 3733,
    31578 => 3730,
    31579 => 3727,
    31580 => 3724,
    31581 => 3721,
    31582 => 3718,
    31583 => 3715,
    31584 => 3712,
    31585 => 3708,
    31586 => 3705,
    31587 => 3702,
    31588 => 3699,
    31589 => 3696,
    31590 => 3693,
    31591 => 3690,
    31592 => 3687,
    31593 => 3683,
    31594 => 3680,
    31595 => 3677,
    31596 => 3674,
    31597 => 3671,
    31598 => 3668,
    31599 => 3665,
    31600 => 3662,
    31601 => 3658,
    31602 => 3655,
    31603 => 3652,
    31604 => 3649,
    31605 => 3646,
    31606 => 3643,
    31607 => 3640,
    31608 => 3637,
    31609 => 3634,
    31610 => 3630,
    31611 => 3627,
    31612 => 3624,
    31613 => 3621,
    31614 => 3618,
    31615 => 3615,
    31616 => 3612,
    31617 => 3609,
    31618 => 3605,
    31619 => 3602,
    31620 => 3599,
    31621 => 3596,
    31622 => 3593,
    31623 => 3590,
    31624 => 3587,
    31625 => 3584,
    31626 => 3580,
    31627 => 3577,
    31628 => 3574,
    31629 => 3571,
    31630 => 3568,
    31631 => 3565,
    31632 => 3562,
    31633 => 3559,
    31634 => 3555,
    31635 => 3552,
    31636 => 3549,
    31637 => 3546,
    31638 => 3543,
    31639 => 3540,
    31640 => 3537,
    31641 => 3534,
    31642 => 3530,
    31643 => 3527,
    31644 => 3524,
    31645 => 3521,
    31646 => 3518,
    31647 => 3515,
    31648 => 3512,
    31649 => 3509,
    31650 => 3505,
    31651 => 3502,
    31652 => 3499,
    31653 => 3496,
    31654 => 3493,
    31655 => 3490,
    31656 => 3487,
    31657 => 3484,
    31658 => 3480,
    31659 => 3477,
    31660 => 3474,
    31661 => 3471,
    31662 => 3468,
    31663 => 3465,
    31664 => 3462,
    31665 => 3459,
    31666 => 3455,
    31667 => 3452,
    31668 => 3449,
    31669 => 3446,
    31670 => 3443,
    31671 => 3440,
    31672 => 3437,
    31673 => 3434,
    31674 => 3430,
    31675 => 3427,
    31676 => 3424,
    31677 => 3421,
    31678 => 3418,
    31679 => 3415,
    31680 => 3412,
    31681 => 3409,
    31682 => 3406,
    31683 => 3402,
    31684 => 3399,
    31685 => 3396,
    31686 => 3393,
    31687 => 3390,
    31688 => 3387,
    31689 => 3384,
    31690 => 3381,
    31691 => 3377,
    31692 => 3374,
    31693 => 3371,
    31694 => 3368,
    31695 => 3365,
    31696 => 3362,
    31697 => 3359,
    31698 => 3356,
    31699 => 3352,
    31700 => 3349,
    31701 => 3346,
    31702 => 3343,
    31703 => 3340,
    31704 => 3337,
    31705 => 3334,
    31706 => 3331,
    31707 => 3327,
    31708 => 3324,
    31709 => 3321,
    31710 => 3318,
    31711 => 3315,
    31712 => 3312,
    31713 => 3309,
    31714 => 3306,
    31715 => 3302,
    31716 => 3299,
    31717 => 3296,
    31718 => 3293,
    31719 => 3290,
    31720 => 3287,
    31721 => 3284,
    31722 => 3281,
    31723 => 3277,
    31724 => 3274,
    31725 => 3271,
    31726 => 3268,
    31727 => 3265,
    31728 => 3262,
    31729 => 3259,
    31730 => 3255,
    31731 => 3252,
    31732 => 3249,
    31733 => 3246,
    31734 => 3243,
    31735 => 3240,
    31736 => 3237,
    31737 => 3234,
    31738 => 3230,
    31739 => 3227,
    31740 => 3224,
    31741 => 3221,
    31742 => 3218,
    31743 => 3215,
    31744 => 3212,
    31745 => 3209,
    31746 => 3205,
    31747 => 3202,
    31748 => 3199,
    31749 => 3196,
    31750 => 3193,
    31751 => 3190,
    31752 => 3187,
    31753 => 3184,
    31754 => 3180,
    31755 => 3177,
    31756 => 3174,
    31757 => 3171,
    31758 => 3168,
    31759 => 3165,
    31760 => 3162,
    31761 => 3159,
    31762 => 3155,
    31763 => 3152,
    31764 => 3149,
    31765 => 3146,
    31766 => 3143,
    31767 => 3140,
    31768 => 3137,
    31769 => 3134,
    31770 => 3130,
    31771 => 3127,
    31772 => 3124,
    31773 => 3121,
    31774 => 3118,
    31775 => 3115,
    31776 => 3112,
    31777 => 3109,
    31778 => 3105,
    31779 => 3102,
    31780 => 3099,
    31781 => 3096,
    31782 => 3093,
    31783 => 3090,
    31784 => 3087,
    31785 => 3084,
    31786 => 3080,
    31787 => 3077,
    31788 => 3074,
    31789 => 3071,
    31790 => 3068,
    31791 => 3065,
    31792 => 3062,
    31793 => 3059,
    31794 => 3055,
    31795 => 3052,
    31796 => 3049,
    31797 => 3046,
    31798 => 3043,
    31799 => 3040,
    31800 => 3037,
    31801 => 3033,
    31802 => 3030,
    31803 => 3027,
    31804 => 3024,
    31805 => 3021,
    31806 => 3018,
    31807 => 3015,
    31808 => 3012,
    31809 => 3008,
    31810 => 3005,
    31811 => 3002,
    31812 => 2999,
    31813 => 2996,
    31814 => 2993,
    31815 => 2990,
    31816 => 2987,
    31817 => 2983,
    31818 => 2980,
    31819 => 2977,
    31820 => 2974,
    31821 => 2971,
    31822 => 2968,
    31823 => 2965,
    31824 => 2962,
    31825 => 2958,
    31826 => 2955,
    31827 => 2952,
    31828 => 2949,
    31829 => 2946,
    31830 => 2943,
    31831 => 2940,
    31832 => 2936,
    31833 => 2933,
    31834 => 2930,
    31835 => 2927,
    31836 => 2924,
    31837 => 2921,
    31838 => 2918,
    31839 => 2915,
    31840 => 2911,
    31841 => 2908,
    31842 => 2905,
    31843 => 2902,
    31844 => 2899,
    31845 => 2896,
    31846 => 2893,
    31847 => 2890,
    31848 => 2886,
    31849 => 2883,
    31850 => 2880,
    31851 => 2877,
    31852 => 2874,
    31853 => 2871,
    31854 => 2868,
    31855 => 2865,
    31856 => 2861,
    31857 => 2858,
    31858 => 2855,
    31859 => 2852,
    31860 => 2849,
    31861 => 2846,
    31862 => 2843,
    31863 => 2839,
    31864 => 2836,
    31865 => 2833,
    31866 => 2830,
    31867 => 2827,
    31868 => 2824,
    31869 => 2821,
    31870 => 2818,
    31871 => 2814,
    31872 => 2811,
    31873 => 2808,
    31874 => 2805,
    31875 => 2802,
    31876 => 2799,
    31877 => 2796,
    31878 => 2793,
    31879 => 2789,
    31880 => 2786,
    31881 => 2783,
    31882 => 2780,
    31883 => 2777,
    31884 => 2774,
    31885 => 2771,
    31886 => 2767,
    31887 => 2764,
    31888 => 2761,
    31889 => 2758,
    31890 => 2755,
    31891 => 2752,
    31892 => 2749,
    31893 => 2746,
    31894 => 2742,
    31895 => 2739,
    31896 => 2736,
    31897 => 2733,
    31898 => 2730,
    31899 => 2727,
    31900 => 2724,
    31901 => 2721,
    31902 => 2717,
    31903 => 2714,
    31904 => 2711,
    31905 => 2708,
    31906 => 2705,
    31907 => 2702,
    31908 => 2699,
    31909 => 2695,
    31910 => 2692,
    31911 => 2689,
    31912 => 2686,
    31913 => 2683,
    31914 => 2680,
    31915 => 2677,
    31916 => 2674,
    31917 => 2670,
    31918 => 2667,
    31919 => 2664,
    31920 => 2661,
    31921 => 2658,
    31922 => 2655,
    31923 => 2652,
    31924 => 2649,
    31925 => 2645,
    31926 => 2642,
    31927 => 2639,
    31928 => 2636,
    31929 => 2633,
    31930 => 2630,
    31931 => 2627,
    31932 => 2623,
    31933 => 2620,
    31934 => 2617,
    31935 => 2614,
    31936 => 2611,
    31937 => 2608,
    31938 => 2605,
    31939 => 2602,
    31940 => 2598,
    31941 => 2595,
    31942 => 2592,
    31943 => 2589,
    31944 => 2586,
    31945 => 2583,
    31946 => 2580,
    31947 => 2577,
    31948 => 2573,
    31949 => 2570,
    31950 => 2567,
    31951 => 2564,
    31952 => 2561,
    31953 => 2558,
    31954 => 2555,
    31955 => 2551,
    31956 => 2548,
    31957 => 2545,
    31958 => 2542,
    31959 => 2539,
    31960 => 2536,
    31961 => 2533,
    31962 => 2530,
    31963 => 2526,
    31964 => 2523,
    31965 => 2520,
    31966 => 2517,
    31967 => 2514,
    31968 => 2511,
    31969 => 2508,
    31970 => 2504,
    31971 => 2501,
    31972 => 2498,
    31973 => 2495,
    31974 => 2492,
    31975 => 2489,
    31976 => 2486,
    31977 => 2483,
    31978 => 2479,
    31979 => 2476,
    31980 => 2473,
    31981 => 2470,
    31982 => 2467,
    31983 => 2464,
    31984 => 2461,
    31985 => 2457,
    31986 => 2454,
    31987 => 2451,
    31988 => 2448,
    31989 => 2445,
    31990 => 2442,
    31991 => 2439,
    31992 => 2436,
    31993 => 2432,
    31994 => 2429,
    31995 => 2426,
    31996 => 2423,
    31997 => 2420,
    31998 => 2417,
    31999 => 2414,
    32000 => 2410,
    32001 => 2407,
    32002 => 2404,
    32003 => 2401,
    32004 => 2398,
    32005 => 2395,
    32006 => 2392,
    32007 => 2389,
    32008 => 2385,
    32009 => 2382,
    32010 => 2379,
    32011 => 2376,
    32012 => 2373,
    32013 => 2370,
    32014 => 2367,
    32015 => 2363,
    32016 => 2360,
    32017 => 2357,
    32018 => 2354,
    32019 => 2351,
    32020 => 2348,
    32021 => 2345,
    32022 => 2342,
    32023 => 2338,
    32024 => 2335,
    32025 => 2332,
    32026 => 2329,
    32027 => 2326,
    32028 => 2323,
    32029 => 2320,
    32030 => 2316,
    32031 => 2313,
    32032 => 2310,
    32033 => 2307,
    32034 => 2304,
    32035 => 2301,
    32036 => 2298,
    32037 => 2295,
    32038 => 2291,
    32039 => 2288,
    32040 => 2285,
    32041 => 2282,
    32042 => 2279,
    32043 => 2276,
    32044 => 2273,
    32045 => 2269,
    32046 => 2266,
    32047 => 2263,
    32048 => 2260,
    32049 => 2257,
    32050 => 2254,
    32051 => 2251,
    32052 => 2248,
    32053 => 2244,
    32054 => 2241,
    32055 => 2238,
    32056 => 2235,
    32057 => 2232,
    32058 => 2229,
    32059 => 2226,
    32060 => 2222,
    32061 => 2219,
    32062 => 2216,
    32063 => 2213,
    32064 => 2210,
    32065 => 2207,
    32066 => 2204,
    32067 => 2201,
    32068 => 2197,
    32069 => 2194,
    32070 => 2191,
    32071 => 2188,
    32072 => 2185,
    32073 => 2182,
    32074 => 2179,
    32075 => 2175,
    32076 => 2172,
    32077 => 2169,
    32078 => 2166,
    32079 => 2163,
    32080 => 2160,
    32081 => 2157,
    32082 => 2154,
    32083 => 2150,
    32084 => 2147,
    32085 => 2144,
    32086 => 2141,
    32087 => 2138,
    32088 => 2135,
    32089 => 2132,
    32090 => 2128,
    32091 => 2125,
    32092 => 2122,
    32093 => 2119,
    32094 => 2116,
    32095 => 2113,
    32096 => 2110,
    32097 => 2106,
    32098 => 2103,
    32099 => 2100,
    32100 => 2097,
    32101 => 2094,
    32102 => 2091,
    32103 => 2088,
    32104 => 2085,
    32105 => 2081,
    32106 => 2078,
    32107 => 2075,
    32108 => 2072,
    32109 => 2069,
    32110 => 2066,
    32111 => 2063,
    32112 => 2059,
    32113 => 2056,
    32114 => 2053,
    32115 => 2050,
    32116 => 2047,
    32117 => 2044,
    32118 => 2041,
    32119 => 2038,
    32120 => 2034,
    32121 => 2031,
    32122 => 2028,
    32123 => 2025,
    32124 => 2022,
    32125 => 2019,
    32126 => 2016,
    32127 => 2012,
    32128 => 2009,
    32129 => 2006,
    32130 => 2003,
    32131 => 2000,
    32132 => 1997,
    32133 => 1994,
    32134 => 1990,
    32135 => 1987,
    32136 => 1984,
    32137 => 1981,
    32138 => 1978,
    32139 => 1975,
    32140 => 1972,
    32141 => 1969,
    32142 => 1965,
    32143 => 1962,
    32144 => 1959,
    32145 => 1956,
    32146 => 1953,
    32147 => 1950,
    32148 => 1947,
    32149 => 1943,
    32150 => 1940,
    32151 => 1937,
    32152 => 1934,
    32153 => 1931,
    32154 => 1928,
    32155 => 1925,
    32156 => 1921,
    32157 => 1918,
    32158 => 1915,
    32159 => 1912,
    32160 => 1909,
    32161 => 1906,
    32162 => 1903,
    32163 => 1900,
    32164 => 1896,
    32165 => 1893,
    32166 => 1890,
    32167 => 1887,
    32168 => 1884,
    32169 => 1881,
    32170 => 1878,
    32171 => 1874,
    32172 => 1871,
    32173 => 1868,
    32174 => 1865,
    32175 => 1862,
    32176 => 1859,
    32177 => 1856,
    32178 => 1852,
    32179 => 1849,
    32180 => 1846,
    32181 => 1843,
    32182 => 1840,
    32183 => 1837,
    32184 => 1834,
    32185 => 1831,
    32186 => 1827,
    32187 => 1824,
    32188 => 1821,
    32189 => 1818,
    32190 => 1815,
    32191 => 1812,
    32192 => 1809,
    32193 => 1805,
    32194 => 1802,
    32195 => 1799,
    32196 => 1796,
    32197 => 1793,
    32198 => 1790,
    32199 => 1787,
    32200 => 1783,
    32201 => 1780,
    32202 => 1777,
    32203 => 1774,
    32204 => 1771,
    32205 => 1768,
    32206 => 1765,
    32207 => 1762,
    32208 => 1758,
    32209 => 1755,
    32210 => 1752,
    32211 => 1749,
    32212 => 1746,
    32213 => 1743,
    32214 => 1740,
    32215 => 1736,
    32216 => 1733,
    32217 => 1730,
    32218 => 1727,
    32219 => 1724,
    32220 => 1721,
    32221 => 1718,
    32222 => 1714,
    32223 => 1711,
    32224 => 1708,
    32225 => 1705,
    32226 => 1702,
    32227 => 1699,
    32228 => 1696,
    32229 => 1693,
    32230 => 1689,
    32231 => 1686,
    32232 => 1683,
    32233 => 1680,
    32234 => 1677,
    32235 => 1674,
    32236 => 1671,
    32237 => 1667,
    32238 => 1664,
    32239 => 1661,
    32240 => 1658,
    32241 => 1655,
    32242 => 1652,
    32243 => 1649,
    32244 => 1645,
    32245 => 1642,
    32246 => 1639,
    32247 => 1636,
    32248 => 1633,
    32249 => 1630,
    32250 => 1627,
    32251 => 1623,
    32252 => 1620,
    32253 => 1617,
    32254 => 1614,
    32255 => 1611,
    32256 => 1608,
    32257 => 1605,
    32258 => 1602,
    32259 => 1598,
    32260 => 1595,
    32261 => 1592,
    32262 => 1589,
    32263 => 1586,
    32264 => 1583,
    32265 => 1580,
    32266 => 1576,
    32267 => 1573,
    32268 => 1570,
    32269 => 1567,
    32270 => 1564,
    32271 => 1561,
    32272 => 1558,
    32273 => 1554,
    32274 => 1551,
    32275 => 1548,
    32276 => 1545,
    32277 => 1542,
    32278 => 1539,
    32279 => 1536,
    32280 => 1532,
    32281 => 1529,
    32282 => 1526,
    32283 => 1523,
    32284 => 1520,
    32285 => 1517,
    32286 => 1514,
    32287 => 1511,
    32288 => 1507,
    32289 => 1504,
    32290 => 1501,
    32291 => 1498,
    32292 => 1495,
    32293 => 1492,
    32294 => 1489,
    32295 => 1485,
    32296 => 1482,
    32297 => 1479,
    32298 => 1476,
    32299 => 1473,
    32300 => 1470,
    32301 => 1467,
    32302 => 1463,
    32303 => 1460,
    32304 => 1457,
    32305 => 1454,
    32306 => 1451,
    32307 => 1448,
    32308 => 1445,
    32309 => 1441,
    32310 => 1438,
    32311 => 1435,
    32312 => 1432,
    32313 => 1429,
    32314 => 1426,
    32315 => 1423,
    32316 => 1420,
    32317 => 1416,
    32318 => 1413,
    32319 => 1410,
    32320 => 1407,
    32321 => 1404,
    32322 => 1401,
    32323 => 1398,
    32324 => 1394,
    32325 => 1391,
    32326 => 1388,
    32327 => 1385,
    32328 => 1382,
    32329 => 1379,
    32330 => 1376,
    32331 => 1372,
    32332 => 1369,
    32333 => 1366,
    32334 => 1363,
    32335 => 1360,
    32336 => 1357,
    32337 => 1354,
    32338 => 1350,
    32339 => 1347,
    32340 => 1344,
    32341 => 1341,
    32342 => 1338,
    32343 => 1335,
    32344 => 1332,
    32345 => 1328,
    32346 => 1325,
    32347 => 1322,
    32348 => 1319,
    32349 => 1316,
    32350 => 1313,
    32351 => 1310,
    32352 => 1307,
    32353 => 1303,
    32354 => 1300,
    32355 => 1297,
    32356 => 1294,
    32357 => 1291,
    32358 => 1288,
    32359 => 1285,
    32360 => 1281,
    32361 => 1278,
    32362 => 1275,
    32363 => 1272,
    32364 => 1269,
    32365 => 1266,
    32366 => 1263,
    32367 => 1259,
    32368 => 1256,
    32369 => 1253,
    32370 => 1250,
    32371 => 1247,
    32372 => 1244,
    32373 => 1241,
    32374 => 1237,
    32375 => 1234,
    32376 => 1231,
    32377 => 1228,
    32378 => 1225,
    32379 => 1222,
    32380 => 1219,
    32381 => 1215,
    32382 => 1212,
    32383 => 1209,
    32384 => 1206,
    32385 => 1203,
    32386 => 1200,
    32387 => 1197,
    32388 => 1194,
    32389 => 1190,
    32390 => 1187,
    32391 => 1184,
    32392 => 1181,
    32393 => 1178,
    32394 => 1175,
    32395 => 1172,
    32396 => 1168,
    32397 => 1165,
    32398 => 1162,
    32399 => 1159,
    32400 => 1156,
    32401 => 1153,
    32402 => 1150,
    32403 => 1146,
    32404 => 1143,
    32405 => 1140,
    32406 => 1137,
    32407 => 1134,
    32408 => 1131,
    32409 => 1128,
    32410 => 1124,
    32411 => 1121,
    32412 => 1118,
    32413 => 1115,
    32414 => 1112,
    32415 => 1109,
    32416 => 1106,
    32417 => 1102,
    32418 => 1099,
    32419 => 1096,
    32420 => 1093,
    32421 => 1090,
    32422 => 1087,
    32423 => 1084,
    32424 => 1080,
    32425 => 1077,
    32426 => 1074,
    32427 => 1071,
    32428 => 1068,
    32429 => 1065,
    32430 => 1062,
    32431 => 1059,
    32432 => 1055,
    32433 => 1052,
    32434 => 1049,
    32435 => 1046,
    32436 => 1043,
    32437 => 1040,
    32438 => 1037,
    32439 => 1033,
    32440 => 1030,
    32441 => 1027,
    32442 => 1024,
    32443 => 1021,
    32444 => 1018,
    32445 => 1015,
    32446 => 1011,
    32447 => 1008,
    32448 => 1005,
    32449 => 1002,
    32450 => 999,
    32451 => 996,
    32452 => 993,
    32453 => 989,
    32454 => 986,
    32455 => 983,
    32456 => 980,
    32457 => 977,
    32458 => 974,
    32459 => 971,
    32460 => 967,
    32461 => 964,
    32462 => 961,
    32463 => 958,
    32464 => 955,
    32465 => 952,
    32466 => 949,
    32467 => 945,
    32468 => 942,
    32469 => 939,
    32470 => 936,
    32471 => 933,
    32472 => 930,
    32473 => 927,
    32474 => 923,
    32475 => 920,
    32476 => 917,
    32477 => 914,
    32478 => 911,
    32479 => 908,
    32480 => 905,
    32481 => 901,
    32482 => 898,
    32483 => 895,
    32484 => 892,
    32485 => 889,
    32486 => 886,
    32487 => 883,
    32488 => 880,
    32489 => 876,
    32490 => 873,
    32491 => 870,
    32492 => 867,
    32493 => 864,
    32494 => 861,
    32495 => 858,
    32496 => 854,
    32497 => 851,
    32498 => 848,
    32499 => 845,
    32500 => 842,
    32501 => 839,
    32502 => 836,
    32503 => 832,
    32504 => 829,
    32505 => 826,
    32506 => 823,
    32507 => 820,
    32508 => 817,
    32509 => 814,
    32510 => 810,
    32511 => 807,
    32512 => 804,
    32513 => 801,
    32514 => 798,
    32515 => 795,
    32516 => 792,
    32517 => 788,
    32518 => 785,
    32519 => 782,
    32520 => 779,
    32521 => 776,
    32522 => 773,
    32523 => 770,
    32524 => 766,
    32525 => 763,
    32526 => 760,
    32527 => 757,
    32528 => 754,
    32529 => 751,
    32530 => 748,
    32531 => 744,
    32532 => 741,
    32533 => 738,
    32534 => 735,
    32535 => 732,
    32536 => 729,
    32537 => 726,
    32538 => 722,
    32539 => 719,
    32540 => 716,
    32541 => 713,
    32542 => 710,
    32543 => 707,
    32544 => 704,
    32545 => 701,
    32546 => 697,
    32547 => 694,
    32548 => 691,
    32549 => 688,
    32550 => 685,
    32551 => 682,
    32552 => 679,
    32553 => 675,
    32554 => 672,
    32555 => 669,
    32556 => 666,
    32557 => 663,
    32558 => 660,
    32559 => 657,
    32560 => 653,
    32561 => 650,
    32562 => 647,
    32563 => 644,
    32564 => 641,
    32565 => 638,
    32566 => 635,
    32567 => 631,
    32568 => 628,
    32569 => 625,
    32570 => 622,
    32571 => 619,
    32572 => 616,
    32573 => 613,
    32574 => 609,
    32575 => 606,
    32576 => 603,
    32577 => 600,
    32578 => 597,
    32579 => 594,
    32580 => 591,
    32581 => 587,
    32582 => 584,
    32583 => 581,
    32584 => 578,
    32585 => 575,
    32586 => 572,
    32587 => 569,
    32588 => 565,
    32589 => 562,
    32590 => 559,
    32591 => 556,
    32592 => 553,
    32593 => 550,
    32594 => 547,
    32595 => 543,
    32596 => 540,
    32597 => 537,
    32598 => 534,
    32599 => 531,
    32600 => 528,
    32601 => 525,
    32602 => 521,
    32603 => 518,
    32604 => 515,
    32605 => 512,
    32606 => 509,
    32607 => 506,
    32608 => 503,
    32609 => 499,
    32610 => 496,
    32611 => 493,
    32612 => 490,
    32613 => 487,
    32614 => 484,
    32615 => 481,
    32616 => 477,
    32617 => 474,
    32618 => 471,
    32619 => 468,
    32620 => 465,
    32621 => 462,
    32622 => 459,
    32623 => 456,
    32624 => 452,
    32625 => 449,
    32626 => 446,
    32627 => 443,
    32628 => 440,
    32629 => 437,
    32630 => 434,
    32631 => 430,
    32632 => 427,
    32633 => 424,
    32634 => 421,
    32635 => 418,
    32636 => 415,
    32637 => 412,
    32638 => 408,
    32639 => 405,
    32640 => 402,
    32641 => 399,
    32642 => 396,
    32643 => 393,
    32644 => 390,
    32645 => 386,
    32646 => 383,
    32647 => 380,
    32648 => 377,
    32649 => 374,
    32650 => 371,
    32651 => 368,
    32652 => 364,
    32653 => 361,
    32654 => 358,
    32655 => 355,
    32656 => 352,
    32657 => 349,
    32658 => 346,
    32659 => 342,
    32660 => 339,
    32661 => 336,
    32662 => 333,
    32663 => 330,
    32664 => 327,
    32665 => 324,
    32666 => 320,
    32667 => 317,
    32668 => 314,
    32669 => 311,
    32670 => 308,
    32671 => 305,
    32672 => 302,
    32673 => 298,
    32674 => 295,
    32675 => 292,
    32676 => 289,
    32677 => 286,
    32678 => 283,
    32679 => 280,
    32680 => 276,
    32681 => 273,
    32682 => 270,
    32683 => 267,
    32684 => 264,
    32685 => 261,
    32686 => 258,
    32687 => 254,
    32688 => 251,
    32689 => 248,
    32690 => 245,
    32691 => 242,
    32692 => 239,
    32693 => 236,
    32694 => 232,
    32695 => 229,
    32696 => 226,
    32697 => 223,
    32698 => 220,
    32699 => 217,
    32700 => 214,
    32701 => 210,
    32702 => 207,
    32703 => 204,
    32704 => 201,
    32705 => 198,
    32706 => 195,
    32707 => 192,
    32708 => 188,
    32709 => 185,
    32710 => 182,
    32711 => 179,
    32712 => 176,
    32713 => 173,
    32714 => 170,
    32715 => 166,
    32716 => 163,
    32717 => 160,
    32718 => 157,
    32719 => 154,
    32720 => 151,
    32721 => 148,
    32722 => 145,
    32723 => 141,
    32724 => 138,
    32725 => 135,
    32726 => 132,
    32727 => 129,
    32728 => 126,
    32729 => 123,
    32730 => 119,
    32731 => 116,
    32732 => 113,
    32733 => 110,
    32734 => 107,
    32735 => 104,
    32736 => 101,
    32737 => 97,
    32738 => 94,
    32739 => 91,
    32740 => 88,
    32741 => 85,
    32742 => 82,
    32743 => 79,
    32744 => 75,
    32745 => 72,
    32746 => 69,
    32747 => 66,
    32748 => 63,
    32749 => 60,
    32750 => 57,
    32751 => 53,
    32752 => 50,
    32753 => 47,
    32754 => 44,
    32755 => 41,
    32756 => 38,
    32757 => 35,
    32758 => 31,
    32759 => 28,
    32760 => 25,
    32761 => 22,
    32762 => 19,
    32763 => 16,
    32764 => 13,
    32765 => 9,
    32766 => 6,
    32767 => 3,
    32768 => 0,
    32769 => -3,
    32770 => -6,
    32771 => -9,
    32772 => -13,
    32773 => -16,
    32774 => -19,
    32775 => -22,
    32776 => -25,
    32777 => -28,
    32778 => -31,
    32779 => -35,
    32780 => -38,
    32781 => -41,
    32782 => -44,
    32783 => -47,
    32784 => -50,
    32785 => -53,
    32786 => -57,
    32787 => -60,
    32788 => -63,
    32789 => -66,
    32790 => -69,
    32791 => -72,
    32792 => -75,
    32793 => -79,
    32794 => -82,
    32795 => -85,
    32796 => -88,
    32797 => -91,
    32798 => -94,
    32799 => -97,
    32800 => -101,
    32801 => -104,
    32802 => -107,
    32803 => -110,
    32804 => -113,
    32805 => -116,
    32806 => -119,
    32807 => -123,
    32808 => -126,
    32809 => -129,
    32810 => -132,
    32811 => -135,
    32812 => -138,
    32813 => -141,
    32814 => -145,
    32815 => -148,
    32816 => -151,
    32817 => -154,
    32818 => -157,
    32819 => -160,
    32820 => -163,
    32821 => -166,
    32822 => -170,
    32823 => -173,
    32824 => -176,
    32825 => -179,
    32826 => -182,
    32827 => -185,
    32828 => -188,
    32829 => -192,
    32830 => -195,
    32831 => -198,
    32832 => -201,
    32833 => -204,
    32834 => -207,
    32835 => -210,
    32836 => -214,
    32837 => -217,
    32838 => -220,
    32839 => -223,
    32840 => -226,
    32841 => -229,
    32842 => -232,
    32843 => -236,
    32844 => -239,
    32845 => -242,
    32846 => -245,
    32847 => -248,
    32848 => -251,
    32849 => -254,
    32850 => -258,
    32851 => -261,
    32852 => -264,
    32853 => -267,
    32854 => -270,
    32855 => -273,
    32856 => -276,
    32857 => -280,
    32858 => -283,
    32859 => -286,
    32860 => -289,
    32861 => -292,
    32862 => -295,
    32863 => -298,
    32864 => -302,
    32865 => -305,
    32866 => -308,
    32867 => -311,
    32868 => -314,
    32869 => -317,
    32870 => -320,
    32871 => -324,
    32872 => -327,
    32873 => -330,
    32874 => -333,
    32875 => -336,
    32876 => -339,
    32877 => -342,
    32878 => -346,
    32879 => -349,
    32880 => -352,
    32881 => -355,
    32882 => -358,
    32883 => -361,
    32884 => -364,
    32885 => -368,
    32886 => -371,
    32887 => -374,
    32888 => -377,
    32889 => -380,
    32890 => -383,
    32891 => -386,
    32892 => -390,
    32893 => -393,
    32894 => -396,
    32895 => -399,
    32896 => -402,
    32897 => -405,
    32898 => -408,
    32899 => -412,
    32900 => -415,
    32901 => -418,
    32902 => -421,
    32903 => -424,
    32904 => -427,
    32905 => -430,
    32906 => -434,
    32907 => -437,
    32908 => -440,
    32909 => -443,
    32910 => -446,
    32911 => -449,
    32912 => -452,
    32913 => -456,
    32914 => -459,
    32915 => -462,
    32916 => -465,
    32917 => -468,
    32918 => -471,
    32919 => -474,
    32920 => -477,
    32921 => -481,
    32922 => -484,
    32923 => -487,
    32924 => -490,
    32925 => -493,
    32926 => -496,
    32927 => -499,
    32928 => -503,
    32929 => -506,
    32930 => -509,
    32931 => -512,
    32932 => -515,
    32933 => -518,
    32934 => -521,
    32935 => -525,
    32936 => -528,
    32937 => -531,
    32938 => -534,
    32939 => -537,
    32940 => -540,
    32941 => -543,
    32942 => -547,
    32943 => -550,
    32944 => -553,
    32945 => -556,
    32946 => -559,
    32947 => -562,
    32948 => -565,
    32949 => -569,
    32950 => -572,
    32951 => -575,
    32952 => -578,
    32953 => -581,
    32954 => -584,
    32955 => -587,
    32956 => -591,
    32957 => -594,
    32958 => -597,
    32959 => -600,
    32960 => -603,
    32961 => -606,
    32962 => -609,
    32963 => -613,
    32964 => -616,
    32965 => -619,
    32966 => -622,
    32967 => -625,
    32968 => -628,
    32969 => -631,
    32970 => -635,
    32971 => -638,
    32972 => -641,
    32973 => -644,
    32974 => -647,
    32975 => -650,
    32976 => -653,
    32977 => -657,
    32978 => -660,
    32979 => -663,
    32980 => -666,
    32981 => -669,
    32982 => -672,
    32983 => -675,
    32984 => -679,
    32985 => -682,
    32986 => -685,
    32987 => -688,
    32988 => -691,
    32989 => -694,
    32990 => -697,
    32991 => -701,
    32992 => -704,
    32993 => -707,
    32994 => -710,
    32995 => -713,
    32996 => -716,
    32997 => -719,
    32998 => -722,
    32999 => -726,
    33000 => -729,
    33001 => -732,
    33002 => -735,
    33003 => -738,
    33004 => -741,
    33005 => -744,
    33006 => -748,
    33007 => -751,
    33008 => -754,
    33009 => -757,
    33010 => -760,
    33011 => -763,
    33012 => -766,
    33013 => -770,
    33014 => -773,
    33015 => -776,
    33016 => -779,
    33017 => -782,
    33018 => -785,
    33019 => -788,
    33020 => -792,
    33021 => -795,
    33022 => -798,
    33023 => -801,
    33024 => -804,
    33025 => -807,
    33026 => -810,
    33027 => -814,
    33028 => -817,
    33029 => -820,
    33030 => -823,
    33031 => -826,
    33032 => -829,
    33033 => -832,
    33034 => -836,
    33035 => -839,
    33036 => -842,
    33037 => -845,
    33038 => -848,
    33039 => -851,
    33040 => -854,
    33041 => -858,
    33042 => -861,
    33043 => -864,
    33044 => -867,
    33045 => -870,
    33046 => -873,
    33047 => -876,
    33048 => -880,
    33049 => -883,
    33050 => -886,
    33051 => -889,
    33052 => -892,
    33053 => -895,
    33054 => -898,
    33055 => -901,
    33056 => -905,
    33057 => -908,
    33058 => -911,
    33059 => -914,
    33060 => -917,
    33061 => -920,
    33062 => -923,
    33063 => -927,
    33064 => -930,
    33065 => -933,
    33066 => -936,
    33067 => -939,
    33068 => -942,
    33069 => -945,
    33070 => -949,
    33071 => -952,
    33072 => -955,
    33073 => -958,
    33074 => -961,
    33075 => -964,
    33076 => -967,
    33077 => -971,
    33078 => -974,
    33079 => -977,
    33080 => -980,
    33081 => -983,
    33082 => -986,
    33083 => -989,
    33084 => -993,
    33085 => -996,
    33086 => -999,
    33087 => -1002,
    33088 => -1005,
    33089 => -1008,
    33090 => -1011,
    33091 => -1015,
    33092 => -1018,
    33093 => -1021,
    33094 => -1024,
    33095 => -1027,
    33096 => -1030,
    33097 => -1033,
    33098 => -1037,
    33099 => -1040,
    33100 => -1043,
    33101 => -1046,
    33102 => -1049,
    33103 => -1052,
    33104 => -1055,
    33105 => -1059,
    33106 => -1062,
    33107 => -1065,
    33108 => -1068,
    33109 => -1071,
    33110 => -1074,
    33111 => -1077,
    33112 => -1080,
    33113 => -1084,
    33114 => -1087,
    33115 => -1090,
    33116 => -1093,
    33117 => -1096,
    33118 => -1099,
    33119 => -1102,
    33120 => -1106,
    33121 => -1109,
    33122 => -1112,
    33123 => -1115,
    33124 => -1118,
    33125 => -1121,
    33126 => -1124,
    33127 => -1128,
    33128 => -1131,
    33129 => -1134,
    33130 => -1137,
    33131 => -1140,
    33132 => -1143,
    33133 => -1146,
    33134 => -1150,
    33135 => -1153,
    33136 => -1156,
    33137 => -1159,
    33138 => -1162,
    33139 => -1165,
    33140 => -1168,
    33141 => -1172,
    33142 => -1175,
    33143 => -1178,
    33144 => -1181,
    33145 => -1184,
    33146 => -1187,
    33147 => -1190,
    33148 => -1194,
    33149 => -1197,
    33150 => -1200,
    33151 => -1203,
    33152 => -1206,
    33153 => -1209,
    33154 => -1212,
    33155 => -1215,
    33156 => -1219,
    33157 => -1222,
    33158 => -1225,
    33159 => -1228,
    33160 => -1231,
    33161 => -1234,
    33162 => -1237,
    33163 => -1241,
    33164 => -1244,
    33165 => -1247,
    33166 => -1250,
    33167 => -1253,
    33168 => -1256,
    33169 => -1259,
    33170 => -1263,
    33171 => -1266,
    33172 => -1269,
    33173 => -1272,
    33174 => -1275,
    33175 => -1278,
    33176 => -1281,
    33177 => -1285,
    33178 => -1288,
    33179 => -1291,
    33180 => -1294,
    33181 => -1297,
    33182 => -1300,
    33183 => -1303,
    33184 => -1307,
    33185 => -1310,
    33186 => -1313,
    33187 => -1316,
    33188 => -1319,
    33189 => -1322,
    33190 => -1325,
    33191 => -1328,
    33192 => -1332,
    33193 => -1335,
    33194 => -1338,
    33195 => -1341,
    33196 => -1344,
    33197 => -1347,
    33198 => -1350,
    33199 => -1354,
    33200 => -1357,
    33201 => -1360,
    33202 => -1363,
    33203 => -1366,
    33204 => -1369,
    33205 => -1372,
    33206 => -1376,
    33207 => -1379,
    33208 => -1382,
    33209 => -1385,
    33210 => -1388,
    33211 => -1391,
    33212 => -1394,
    33213 => -1398,
    33214 => -1401,
    33215 => -1404,
    33216 => -1407,
    33217 => -1410,
    33218 => -1413,
    33219 => -1416,
    33220 => -1420,
    33221 => -1423,
    33222 => -1426,
    33223 => -1429,
    33224 => -1432,
    33225 => -1435,
    33226 => -1438,
    33227 => -1441,
    33228 => -1445,
    33229 => -1448,
    33230 => -1451,
    33231 => -1454,
    33232 => -1457,
    33233 => -1460,
    33234 => -1463,
    33235 => -1467,
    33236 => -1470,
    33237 => -1473,
    33238 => -1476,
    33239 => -1479,
    33240 => -1482,
    33241 => -1485,
    33242 => -1489,
    33243 => -1492,
    33244 => -1495,
    33245 => -1498,
    33246 => -1501,
    33247 => -1504,
    33248 => -1507,
    33249 => -1511,
    33250 => -1514,
    33251 => -1517,
    33252 => -1520,
    33253 => -1523,
    33254 => -1526,
    33255 => -1529,
    33256 => -1532,
    33257 => -1536,
    33258 => -1539,
    33259 => -1542,
    33260 => -1545,
    33261 => -1548,
    33262 => -1551,
    33263 => -1554,
    33264 => -1558,
    33265 => -1561,
    33266 => -1564,
    33267 => -1567,
    33268 => -1570,
    33269 => -1573,
    33270 => -1576,
    33271 => -1580,
    33272 => -1583,
    33273 => -1586,
    33274 => -1589,
    33275 => -1592,
    33276 => -1595,
    33277 => -1598,
    33278 => -1602,
    33279 => -1605,
    33280 => -1608,
    33281 => -1611,
    33282 => -1614,
    33283 => -1617,
    33284 => -1620,
    33285 => -1623,
    33286 => -1627,
    33287 => -1630,
    33288 => -1633,
    33289 => -1636,
    33290 => -1639,
    33291 => -1642,
    33292 => -1645,
    33293 => -1649,
    33294 => -1652,
    33295 => -1655,
    33296 => -1658,
    33297 => -1661,
    33298 => -1664,
    33299 => -1667,
    33300 => -1671,
    33301 => -1674,
    33302 => -1677,
    33303 => -1680,
    33304 => -1683,
    33305 => -1686,
    33306 => -1689,
    33307 => -1693,
    33308 => -1696,
    33309 => -1699,
    33310 => -1702,
    33311 => -1705,
    33312 => -1708,
    33313 => -1711,
    33314 => -1714,
    33315 => -1718,
    33316 => -1721,
    33317 => -1724,
    33318 => -1727,
    33319 => -1730,
    33320 => -1733,
    33321 => -1736,
    33322 => -1740,
    33323 => -1743,
    33324 => -1746,
    33325 => -1749,
    33326 => -1752,
    33327 => -1755,
    33328 => -1758,
    33329 => -1762,
    33330 => -1765,
    33331 => -1768,
    33332 => -1771,
    33333 => -1774,
    33334 => -1777,
    33335 => -1780,
    33336 => -1783,
    33337 => -1787,
    33338 => -1790,
    33339 => -1793,
    33340 => -1796,
    33341 => -1799,
    33342 => -1802,
    33343 => -1805,
    33344 => -1809,
    33345 => -1812,
    33346 => -1815,
    33347 => -1818,
    33348 => -1821,
    33349 => -1824,
    33350 => -1827,
    33351 => -1831,
    33352 => -1834,
    33353 => -1837,
    33354 => -1840,
    33355 => -1843,
    33356 => -1846,
    33357 => -1849,
    33358 => -1852,
    33359 => -1856,
    33360 => -1859,
    33361 => -1862,
    33362 => -1865,
    33363 => -1868,
    33364 => -1871,
    33365 => -1874,
    33366 => -1878,
    33367 => -1881,
    33368 => -1884,
    33369 => -1887,
    33370 => -1890,
    33371 => -1893,
    33372 => -1896,
    33373 => -1900,
    33374 => -1903,
    33375 => -1906,
    33376 => -1909,
    33377 => -1912,
    33378 => -1915,
    33379 => -1918,
    33380 => -1921,
    33381 => -1925,
    33382 => -1928,
    33383 => -1931,
    33384 => -1934,
    33385 => -1937,
    33386 => -1940,
    33387 => -1943,
    33388 => -1947,
    33389 => -1950,
    33390 => -1953,
    33391 => -1956,
    33392 => -1959,
    33393 => -1962,
    33394 => -1965,
    33395 => -1969,
    33396 => -1972,
    33397 => -1975,
    33398 => -1978,
    33399 => -1981,
    33400 => -1984,
    33401 => -1987,
    33402 => -1990,
    33403 => -1994,
    33404 => -1997,
    33405 => -2000,
    33406 => -2003,
    33407 => -2006,
    33408 => -2009,
    33409 => -2012,
    33410 => -2016,
    33411 => -2019,
    33412 => -2022,
    33413 => -2025,
    33414 => -2028,
    33415 => -2031,
    33416 => -2034,
    33417 => -2038,
    33418 => -2041,
    33419 => -2044,
    33420 => -2047,
    33421 => -2050,
    33422 => -2053,
    33423 => -2056,
    33424 => -2059,
    33425 => -2063,
    33426 => -2066,
    33427 => -2069,
    33428 => -2072,
    33429 => -2075,
    33430 => -2078,
    33431 => -2081,
    33432 => -2085,
    33433 => -2088,
    33434 => -2091,
    33435 => -2094,
    33436 => -2097,
    33437 => -2100,
    33438 => -2103,
    33439 => -2106,
    33440 => -2110,
    33441 => -2113,
    33442 => -2116,
    33443 => -2119,
    33444 => -2122,
    33445 => -2125,
    33446 => -2128,
    33447 => -2132,
    33448 => -2135,
    33449 => -2138,
    33450 => -2141,
    33451 => -2144,
    33452 => -2147,
    33453 => -2150,
    33454 => -2154,
    33455 => -2157,
    33456 => -2160,
    33457 => -2163,
    33458 => -2166,
    33459 => -2169,
    33460 => -2172,
    33461 => -2175,
    33462 => -2179,
    33463 => -2182,
    33464 => -2185,
    33465 => -2188,
    33466 => -2191,
    33467 => -2194,
    33468 => -2197,
    33469 => -2201,
    33470 => -2204,
    33471 => -2207,
    33472 => -2210,
    33473 => -2213,
    33474 => -2216,
    33475 => -2219,
    33476 => -2222,
    33477 => -2226,
    33478 => -2229,
    33479 => -2232,
    33480 => -2235,
    33481 => -2238,
    33482 => -2241,
    33483 => -2244,
    33484 => -2248,
    33485 => -2251,
    33486 => -2254,
    33487 => -2257,
    33488 => -2260,
    33489 => -2263,
    33490 => -2266,
    33491 => -2269,
    33492 => -2273,
    33493 => -2276,
    33494 => -2279,
    33495 => -2282,
    33496 => -2285,
    33497 => -2288,
    33498 => -2291,
    33499 => -2295,
    33500 => -2298,
    33501 => -2301,
    33502 => -2304,
    33503 => -2307,
    33504 => -2310,
    33505 => -2313,
    33506 => -2316,
    33507 => -2320,
    33508 => -2323,
    33509 => -2326,
    33510 => -2329,
    33511 => -2332,
    33512 => -2335,
    33513 => -2338,
    33514 => -2342,
    33515 => -2345,
    33516 => -2348,
    33517 => -2351,
    33518 => -2354,
    33519 => -2357,
    33520 => -2360,
    33521 => -2363,
    33522 => -2367,
    33523 => -2370,
    33524 => -2373,
    33525 => -2376,
    33526 => -2379,
    33527 => -2382,
    33528 => -2385,
    33529 => -2389,
    33530 => -2392,
    33531 => -2395,
    33532 => -2398,
    33533 => -2401,
    33534 => -2404,
    33535 => -2407,
    33536 => -2410,
    33537 => -2414,
    33538 => -2417,
    33539 => -2420,
    33540 => -2423,
    33541 => -2426,
    33542 => -2429,
    33543 => -2432,
    33544 => -2436,
    33545 => -2439,
    33546 => -2442,
    33547 => -2445,
    33548 => -2448,
    33549 => -2451,
    33550 => -2454,
    33551 => -2457,
    33552 => -2461,
    33553 => -2464,
    33554 => -2467,
    33555 => -2470,
    33556 => -2473,
    33557 => -2476,
    33558 => -2479,
    33559 => -2483,
    33560 => -2486,
    33561 => -2489,
    33562 => -2492,
    33563 => -2495,
    33564 => -2498,
    33565 => -2501,
    33566 => -2504,
    33567 => -2508,
    33568 => -2511,
    33569 => -2514,
    33570 => -2517,
    33571 => -2520,
    33572 => -2523,
    33573 => -2526,
    33574 => -2530,
    33575 => -2533,
    33576 => -2536,
    33577 => -2539,
    33578 => -2542,
    33579 => -2545,
    33580 => -2548,
    33581 => -2551,
    33582 => -2555,
    33583 => -2558,
    33584 => -2561,
    33585 => -2564,
    33586 => -2567,
    33587 => -2570,
    33588 => -2573,
    33589 => -2577,
    33590 => -2580,
    33591 => -2583,
    33592 => -2586,
    33593 => -2589,
    33594 => -2592,
    33595 => -2595,
    33596 => -2598,
    33597 => -2602,
    33598 => -2605,
    33599 => -2608,
    33600 => -2611,
    33601 => -2614,
    33602 => -2617,
    33603 => -2620,
    33604 => -2623,
    33605 => -2627,
    33606 => -2630,
    33607 => -2633,
    33608 => -2636,
    33609 => -2639,
    33610 => -2642,
    33611 => -2645,
    33612 => -2649,
    33613 => -2652,
    33614 => -2655,
    33615 => -2658,
    33616 => -2661,
    33617 => -2664,
    33618 => -2667,
    33619 => -2670,
    33620 => -2674,
    33621 => -2677,
    33622 => -2680,
    33623 => -2683,
    33624 => -2686,
    33625 => -2689,
    33626 => -2692,
    33627 => -2695,
    33628 => -2699,
    33629 => -2702,
    33630 => -2705,
    33631 => -2708,
    33632 => -2711,
    33633 => -2714,
    33634 => -2717,
    33635 => -2721,
    33636 => -2724,
    33637 => -2727,
    33638 => -2730,
    33639 => -2733,
    33640 => -2736,
    33641 => -2739,
    33642 => -2742,
    33643 => -2746,
    33644 => -2749,
    33645 => -2752,
    33646 => -2755,
    33647 => -2758,
    33648 => -2761,
    33649 => -2764,
    33650 => -2767,
    33651 => -2771,
    33652 => -2774,
    33653 => -2777,
    33654 => -2780,
    33655 => -2783,
    33656 => -2786,
    33657 => -2789,
    33658 => -2793,
    33659 => -2796,
    33660 => -2799,
    33661 => -2802,
    33662 => -2805,
    33663 => -2808,
    33664 => -2811,
    33665 => -2814,
    33666 => -2818,
    33667 => -2821,
    33668 => -2824,
    33669 => -2827,
    33670 => -2830,
    33671 => -2833,
    33672 => -2836,
    33673 => -2839,
    33674 => -2843,
    33675 => -2846,
    33676 => -2849,
    33677 => -2852,
    33678 => -2855,
    33679 => -2858,
    33680 => -2861,
    33681 => -2865,
    33682 => -2868,
    33683 => -2871,
    33684 => -2874,
    33685 => -2877,
    33686 => -2880,
    33687 => -2883,
    33688 => -2886,
    33689 => -2890,
    33690 => -2893,
    33691 => -2896,
    33692 => -2899,
    33693 => -2902,
    33694 => -2905,
    33695 => -2908,
    33696 => -2911,
    33697 => -2915,
    33698 => -2918,
    33699 => -2921,
    33700 => -2924,
    33701 => -2927,
    33702 => -2930,
    33703 => -2933,
    33704 => -2936,
    33705 => -2940,
    33706 => -2943,
    33707 => -2946,
    33708 => -2949,
    33709 => -2952,
    33710 => -2955,
    33711 => -2958,
    33712 => -2962,
    33713 => -2965,
    33714 => -2968,
    33715 => -2971,
    33716 => -2974,
    33717 => -2977,
    33718 => -2980,
    33719 => -2983,
    33720 => -2987,
    33721 => -2990,
    33722 => -2993,
    33723 => -2996,
    33724 => -2999,
    33725 => -3002,
    33726 => -3005,
    33727 => -3008,
    33728 => -3012,
    33729 => -3015,
    33730 => -3018,
    33731 => -3021,
    33732 => -3024,
    33733 => -3027,
    33734 => -3030,
    33735 => -3033,
    33736 => -3037,
    33737 => -3040,
    33738 => -3043,
    33739 => -3046,
    33740 => -3049,
    33741 => -3052,
    33742 => -3055,
    33743 => -3059,
    33744 => -3062,
    33745 => -3065,
    33746 => -3068,
    33747 => -3071,
    33748 => -3074,
    33749 => -3077,
    33750 => -3080,
    33751 => -3084,
    33752 => -3087,
    33753 => -3090,
    33754 => -3093,
    33755 => -3096,
    33756 => -3099,
    33757 => -3102,
    33758 => -3105,
    33759 => -3109,
    33760 => -3112,
    33761 => -3115,
    33762 => -3118,
    33763 => -3121,
    33764 => -3124,
    33765 => -3127,
    33766 => -3130,
    33767 => -3134,
    33768 => -3137,
    33769 => -3140,
    33770 => -3143,
    33771 => -3146,
    33772 => -3149,
    33773 => -3152,
    33774 => -3155,
    33775 => -3159,
    33776 => -3162,
    33777 => -3165,
    33778 => -3168,
    33779 => -3171,
    33780 => -3174,
    33781 => -3177,
    33782 => -3180,
    33783 => -3184,
    33784 => -3187,
    33785 => -3190,
    33786 => -3193,
    33787 => -3196,
    33788 => -3199,
    33789 => -3202,
    33790 => -3205,
    33791 => -3209,
    33792 => -3212,
    33793 => -3215,
    33794 => -3218,
    33795 => -3221,
    33796 => -3224,
    33797 => -3227,
    33798 => -3230,
    33799 => -3234,
    33800 => -3237,
    33801 => -3240,
    33802 => -3243,
    33803 => -3246,
    33804 => -3249,
    33805 => -3252,
    33806 => -3255,
    33807 => -3259,
    33808 => -3262,
    33809 => -3265,
    33810 => -3268,
    33811 => -3271,
    33812 => -3274,
    33813 => -3277,
    33814 => -3281,
    33815 => -3284,
    33816 => -3287,
    33817 => -3290,
    33818 => -3293,
    33819 => -3296,
    33820 => -3299,
    33821 => -3302,
    33822 => -3306,
    33823 => -3309,
    33824 => -3312,
    33825 => -3315,
    33826 => -3318,
    33827 => -3321,
    33828 => -3324,
    33829 => -3327,
    33830 => -3331,
    33831 => -3334,
    33832 => -3337,
    33833 => -3340,
    33834 => -3343,
    33835 => -3346,
    33836 => -3349,
    33837 => -3352,
    33838 => -3356,
    33839 => -3359,
    33840 => -3362,
    33841 => -3365,
    33842 => -3368,
    33843 => -3371,
    33844 => -3374,
    33845 => -3377,
    33846 => -3381,
    33847 => -3384,
    33848 => -3387,
    33849 => -3390,
    33850 => -3393,
    33851 => -3396,
    33852 => -3399,
    33853 => -3402,
    33854 => -3406,
    33855 => -3409,
    33856 => -3412,
    33857 => -3415,
    33858 => -3418,
    33859 => -3421,
    33860 => -3424,
    33861 => -3427,
    33862 => -3430,
    33863 => -3434,
    33864 => -3437,
    33865 => -3440,
    33866 => -3443,
    33867 => -3446,
    33868 => -3449,
    33869 => -3452,
    33870 => -3455,
    33871 => -3459,
    33872 => -3462,
    33873 => -3465,
    33874 => -3468,
    33875 => -3471,
    33876 => -3474,
    33877 => -3477,
    33878 => -3480,
    33879 => -3484,
    33880 => -3487,
    33881 => -3490,
    33882 => -3493,
    33883 => -3496,
    33884 => -3499,
    33885 => -3502,
    33886 => -3505,
    33887 => -3509,
    33888 => -3512,
    33889 => -3515,
    33890 => -3518,
    33891 => -3521,
    33892 => -3524,
    33893 => -3527,
    33894 => -3530,
    33895 => -3534,
    33896 => -3537,
    33897 => -3540,
    33898 => -3543,
    33899 => -3546,
    33900 => -3549,
    33901 => -3552,
    33902 => -3555,
    33903 => -3559,
    33904 => -3562,
    33905 => -3565,
    33906 => -3568,
    33907 => -3571,
    33908 => -3574,
    33909 => -3577,
    33910 => -3580,
    33911 => -3584,
    33912 => -3587,
    33913 => -3590,
    33914 => -3593,
    33915 => -3596,
    33916 => -3599,
    33917 => -3602,
    33918 => -3605,
    33919 => -3609,
    33920 => -3612,
    33921 => -3615,
    33922 => -3618,
    33923 => -3621,
    33924 => -3624,
    33925 => -3627,
    33926 => -3630,
    33927 => -3634,
    33928 => -3637,
    33929 => -3640,
    33930 => -3643,
    33931 => -3646,
    33932 => -3649,
    33933 => -3652,
    33934 => -3655,
    33935 => -3658,
    33936 => -3662,
    33937 => -3665,
    33938 => -3668,
    33939 => -3671,
    33940 => -3674,
    33941 => -3677,
    33942 => -3680,
    33943 => -3683,
    33944 => -3687,
    33945 => -3690,
    33946 => -3693,
    33947 => -3696,
    33948 => -3699,
    33949 => -3702,
    33950 => -3705,
    33951 => -3708,
    33952 => -3712,
    33953 => -3715,
    33954 => -3718,
    33955 => -3721,
    33956 => -3724,
    33957 => -3727,
    33958 => -3730,
    33959 => -3733,
    33960 => -3737,
    33961 => -3740,
    33962 => -3743,
    33963 => -3746,
    33964 => -3749,
    33965 => -3752,
    33966 => -3755,
    33967 => -3758,
    33968 => -3761,
    33969 => -3765,
    33970 => -3768,
    33971 => -3771,
    33972 => -3774,
    33973 => -3777,
    33974 => -3780,
    33975 => -3783,
    33976 => -3786,
    33977 => -3790,
    33978 => -3793,
    33979 => -3796,
    33980 => -3799,
    33981 => -3802,
    33982 => -3805,
    33983 => -3808,
    33984 => -3811,
    33985 => -3815,
    33986 => -3818,
    33987 => -3821,
    33988 => -3824,
    33989 => -3827,
    33990 => -3830,
    33991 => -3833,
    33992 => -3836,
    33993 => -3839,
    33994 => -3843,
    33995 => -3846,
    33996 => -3849,
    33997 => -3852,
    33998 => -3855,
    33999 => -3858,
    34000 => -3861,
    34001 => -3864,
    34002 => -3868,
    34003 => -3871,
    34004 => -3874,
    34005 => -3877,
    34006 => -3880,
    34007 => -3883,
    34008 => -3886,
    34009 => -3889,
    34010 => -3893,
    34011 => -3896,
    34012 => -3899,
    34013 => -3902,
    34014 => -3905,
    34015 => -3908,
    34016 => -3911,
    34017 => -3914,
    34018 => -3917,
    34019 => -3921,
    34020 => -3924,
    34021 => -3927,
    34022 => -3930,
    34023 => -3933,
    34024 => -3936,
    34025 => -3939,
    34026 => -3942,
    34027 => -3946,
    34028 => -3949,
    34029 => -3952,
    34030 => -3955,
    34031 => -3958,
    34032 => -3961,
    34033 => -3964,
    34034 => -3967,
    34035 => -3970,
    34036 => -3974,
    34037 => -3977,
    34038 => -3980,
    34039 => -3983,
    34040 => -3986,
    34041 => -3989,
    34042 => -3992,
    34043 => -3995,
    34044 => -3999,
    34045 => -4002,
    34046 => -4005,
    34047 => -4008,
    34048 => -4011,
    34049 => -4014,
    34050 => -4017,
    34051 => -4020,
    34052 => -4024,
    34053 => -4027,
    34054 => -4030,
    34055 => -4033,
    34056 => -4036,
    34057 => -4039,
    34058 => -4042,
    34059 => -4045,
    34060 => -4048,
    34061 => -4052,
    34062 => -4055,
    34063 => -4058,
    34064 => -4061,
    34065 => -4064,
    34066 => -4067,
    34067 => -4070,
    34068 => -4073,
    34069 => -4076,
    34070 => -4080,
    34071 => -4083,
    34072 => -4086,
    34073 => -4089,
    34074 => -4092,
    34075 => -4095,
    34076 => -4098,
    34077 => -4101,
    34078 => -4105,
    34079 => -4108,
    34080 => -4111,
    34081 => -4114,
    34082 => -4117,
    34083 => -4120,
    34084 => -4123,
    34085 => -4126,
    34086 => -4129,
    34087 => -4133,
    34088 => -4136,
    34089 => -4139,
    34090 => -4142,
    34091 => -4145,
    34092 => -4148,
    34093 => -4151,
    34094 => -4154,
    34095 => -4158,
    34096 => -4161,
    34097 => -4164,
    34098 => -4167,
    34099 => -4170,
    34100 => -4173,
    34101 => -4176,
    34102 => -4179,
    34103 => -4182,
    34104 => -4186,
    34105 => -4189,
    34106 => -4192,
    34107 => -4195,
    34108 => -4198,
    34109 => -4201,
    34110 => -4204,
    34111 => -4207,
    34112 => -4210,
    34113 => -4214,
    34114 => -4217,
    34115 => -4220,
    34116 => -4223,
    34117 => -4226,
    34118 => -4229,
    34119 => -4232,
    34120 => -4235,
    34121 => -4239,
    34122 => -4242,
    34123 => -4245,
    34124 => -4248,
    34125 => -4251,
    34126 => -4254,
    34127 => -4257,
    34128 => -4260,
    34129 => -4263,
    34130 => -4267,
    34131 => -4270,
    34132 => -4273,
    34133 => -4276,
    34134 => -4279,
    34135 => -4282,
    34136 => -4285,
    34137 => -4288,
    34138 => -4291,
    34139 => -4295,
    34140 => -4298,
    34141 => -4301,
    34142 => -4304,
    34143 => -4307,
    34144 => -4310,
    34145 => -4313,
    34146 => -4316,
    34147 => -4320,
    34148 => -4323,
    34149 => -4326,
    34150 => -4329,
    34151 => -4332,
    34152 => -4335,
    34153 => -4338,
    34154 => -4341,
    34155 => -4344,
    34156 => -4348,
    34157 => -4351,
    34158 => -4354,
    34159 => -4357,
    34160 => -4360,
    34161 => -4363,
    34162 => -4366,
    34163 => -4369,
    34164 => -4372,
    34165 => -4376,
    34166 => -4379,
    34167 => -4382,
    34168 => -4385,
    34169 => -4388,
    34170 => -4391,
    34171 => -4394,
    34172 => -4397,
    34173 => -4400,
    34174 => -4404,
    34175 => -4407,
    34176 => -4410,
    34177 => -4413,
    34178 => -4416,
    34179 => -4419,
    34180 => -4422,
    34181 => -4425,
    34182 => -4428,
    34183 => -4432,
    34184 => -4435,
    34185 => -4438,
    34186 => -4441,
    34187 => -4444,
    34188 => -4447,
    34189 => -4450,
    34190 => -4453,
    34191 => -4456,
    34192 => -4460,
    34193 => -4463,
    34194 => -4466,
    34195 => -4469,
    34196 => -4472,
    34197 => -4475,
    34198 => -4478,
    34199 => -4481,
    34200 => -4485,
    34201 => -4488,
    34202 => -4491,
    34203 => -4494,
    34204 => -4497,
    34205 => -4500,
    34206 => -4503,
    34207 => -4506,
    34208 => -4509,
    34209 => -4513,
    34210 => -4516,
    34211 => -4519,
    34212 => -4522,
    34213 => -4525,
    34214 => -4528,
    34215 => -4531,
    34216 => -4534,
    34217 => -4537,
    34218 => -4541,
    34219 => -4544,
    34220 => -4547,
    34221 => -4550,
    34222 => -4553,
    34223 => -4556,
    34224 => -4559,
    34225 => -4562,
    34226 => -4565,
    34227 => -4569,
    34228 => -4572,
    34229 => -4575,
    34230 => -4578,
    34231 => -4581,
    34232 => -4584,
    34233 => -4587,
    34234 => -4590,
    34235 => -4593,
    34236 => -4597,
    34237 => -4600,
    34238 => -4603,
    34239 => -4606,
    34240 => -4609,
    34241 => -4612,
    34242 => -4615,
    34243 => -4618,
    34244 => -4621,
    34245 => -4624,
    34246 => -4628,
    34247 => -4631,
    34248 => -4634,
    34249 => -4637,
    34250 => -4640,
    34251 => -4643,
    34252 => -4646,
    34253 => -4649,
    34254 => -4652,
    34255 => -4656,
    34256 => -4659,
    34257 => -4662,
    34258 => -4665,
    34259 => -4668,
    34260 => -4671,
    34261 => -4674,
    34262 => -4677,
    34263 => -4680,
    34264 => -4684,
    34265 => -4687,
    34266 => -4690,
    34267 => -4693,
    34268 => -4696,
    34269 => -4699,
    34270 => -4702,
    34271 => -4705,
    34272 => -4708,
    34273 => -4712,
    34274 => -4715,
    34275 => -4718,
    34276 => -4721,
    34277 => -4724,
    34278 => -4727,
    34279 => -4730,
    34280 => -4733,
    34281 => -4736,
    34282 => -4740,
    34283 => -4743,
    34284 => -4746,
    34285 => -4749,
    34286 => -4752,
    34287 => -4755,
    34288 => -4758,
    34289 => -4761,
    34290 => -4764,
    34291 => -4768,
    34292 => -4771,
    34293 => -4774,
    34294 => -4777,
    34295 => -4780,
    34296 => -4783,
    34297 => -4786,
    34298 => -4789,
    34299 => -4792,
    34300 => -4795,
    34301 => -4799,
    34302 => -4802,
    34303 => -4805,
    34304 => -4808,
    34305 => -4811,
    34306 => -4814,
    34307 => -4817,
    34308 => -4820,
    34309 => -4823,
    34310 => -4827,
    34311 => -4830,
    34312 => -4833,
    34313 => -4836,
    34314 => -4839,
    34315 => -4842,
    34316 => -4845,
    34317 => -4848,
    34318 => -4851,
    34319 => -4855,
    34320 => -4858,
    34321 => -4861,
    34322 => -4864,
    34323 => -4867,
    34324 => -4870,
    34325 => -4873,
    34326 => -4876,
    34327 => -4879,
    34328 => -4882,
    34329 => -4886,
    34330 => -4889,
    34331 => -4892,
    34332 => -4895,
    34333 => -4898,
    34334 => -4901,
    34335 => -4904,
    34336 => -4907,
    34337 => -4910,
    34338 => -4914,
    34339 => -4917,
    34340 => -4920,
    34341 => -4923,
    34342 => -4926,
    34343 => -4929,
    34344 => -4932,
    34345 => -4935,
    34346 => -4938,
    34347 => -4941,
    34348 => -4945,
    34349 => -4948,
    34350 => -4951,
    34351 => -4954,
    34352 => -4957,
    34353 => -4960,
    34354 => -4963,
    34355 => -4966,
    34356 => -4969,
    34357 => -4973,
    34358 => -4976,
    34359 => -4979,
    34360 => -4982,
    34361 => -4985,
    34362 => -4988,
    34363 => -4991,
    34364 => -4994,
    34365 => -4997,
    34366 => -5000,
    34367 => -5004,
    34368 => -5007,
    34369 => -5010,
    34370 => -5013,
    34371 => -5016,
    34372 => -5019,
    34373 => -5022,
    34374 => -5025,
    34375 => -5028,
    34376 => -5032,
    34377 => -5035,
    34378 => -5038,
    34379 => -5041,
    34380 => -5044,
    34381 => -5047,
    34382 => -5050,
    34383 => -5053,
    34384 => -5056,
    34385 => -5059,
    34386 => -5063,
    34387 => -5066,
    34388 => -5069,
    34389 => -5072,
    34390 => -5075,
    34391 => -5078,
    34392 => -5081,
    34393 => -5084,
    34394 => -5087,
    34395 => -5091,
    34396 => -5094,
    34397 => -5097,
    34398 => -5100,
    34399 => -5103,
    34400 => -5106,
    34401 => -5109,
    34402 => -5112,
    34403 => -5115,
    34404 => -5118,
    34405 => -5122,
    34406 => -5125,
    34407 => -5128,
    34408 => -5131,
    34409 => -5134,
    34410 => -5137,
    34411 => -5140,
    34412 => -5143,
    34413 => -5146,
    34414 => -5149,
    34415 => -5153,
    34416 => -5156,
    34417 => -5159,
    34418 => -5162,
    34419 => -5165,
    34420 => -5168,
    34421 => -5171,
    34422 => -5174,
    34423 => -5177,
    34424 => -5180,
    34425 => -5184,
    34426 => -5187,
    34427 => -5190,
    34428 => -5193,
    34429 => -5196,
    34430 => -5199,
    34431 => -5202,
    34432 => -5205,
    34433 => -5208,
    34434 => -5212,
    34435 => -5215,
    34436 => -5218,
    34437 => -5221,
    34438 => -5224,
    34439 => -5227,
    34440 => -5230,
    34441 => -5233,
    34442 => -5236,
    34443 => -5239,
    34444 => -5243,
    34445 => -5246,
    34446 => -5249,
    34447 => -5252,
    34448 => -5255,
    34449 => -5258,
    34450 => -5261,
    34451 => -5264,
    34452 => -5267,
    34453 => -5270,
    34454 => -5274,
    34455 => -5277,
    34456 => -5280,
    34457 => -5283,
    34458 => -5286,
    34459 => -5289,
    34460 => -5292,
    34461 => -5295,
    34462 => -5298,
    34463 => -5301,
    34464 => -5305,
    34465 => -5308,
    34466 => -5311,
    34467 => -5314,
    34468 => -5317,
    34469 => -5320,
    34470 => -5323,
    34471 => -5326,
    34472 => -5329,
    34473 => -5332,
    34474 => -5336,
    34475 => -5339,
    34476 => -5342,
    34477 => -5345,
    34478 => -5348,
    34479 => -5351,
    34480 => -5354,
    34481 => -5357,
    34482 => -5360,
    34483 => -5363,
    34484 => -5367,
    34485 => -5370,
    34486 => -5373,
    34487 => -5376,
    34488 => -5379,
    34489 => -5382,
    34490 => -5385,
    34491 => -5388,
    34492 => -5391,
    34493 => -5394,
    34494 => -5398,
    34495 => -5401,
    34496 => -5404,
    34497 => -5407,
    34498 => -5410,
    34499 => -5413,
    34500 => -5416,
    34501 => -5419,
    34502 => -5422,
    34503 => -5425,
    34504 => -5428,
    34505 => -5432,
    34506 => -5435,
    34507 => -5438,
    34508 => -5441,
    34509 => -5444,
    34510 => -5447,
    34511 => -5450,
    34512 => -5453,
    34513 => -5456,
    34514 => -5459,
    34515 => -5463,
    34516 => -5466,
    34517 => -5469,
    34518 => -5472,
    34519 => -5475,
    34520 => -5478,
    34521 => -5481,
    34522 => -5484,
    34523 => -5487,
    34524 => -5490,
    34525 => -5494,
    34526 => -5497,
    34527 => -5500,
    34528 => -5503,
    34529 => -5506,
    34530 => -5509,
    34531 => -5512,
    34532 => -5515,
    34533 => -5518,
    34534 => -5521,
    34535 => -5525,
    34536 => -5528,
    34537 => -5531,
    34538 => -5534,
    34539 => -5537,
    34540 => -5540,
    34541 => -5543,
    34542 => -5546,
    34543 => -5549,
    34544 => -5552,
    34545 => -5555,
    34546 => -5559,
    34547 => -5562,
    34548 => -5565,
    34549 => -5568,
    34550 => -5571,
    34551 => -5574,
    34552 => -5577,
    34553 => -5580,
    34554 => -5583,
    34555 => -5586,
    34556 => -5590,
    34557 => -5593,
    34558 => -5596,
    34559 => -5599,
    34560 => -5602,
    34561 => -5605,
    34562 => -5608,
    34563 => -5611,
    34564 => -5614,
    34565 => -5617,
    34566 => -5620,
    34567 => -5624,
    34568 => -5627,
    34569 => -5630,
    34570 => -5633,
    34571 => -5636,
    34572 => -5639,
    34573 => -5642,
    34574 => -5645,
    34575 => -5648,
    34576 => -5651,
    34577 => -5655,
    34578 => -5658,
    34579 => -5661,
    34580 => -5664,
    34581 => -5667,
    34582 => -5670,
    34583 => -5673,
    34584 => -5676,
    34585 => -5679,
    34586 => -5682,
    34587 => -5685,
    34588 => -5689,
    34589 => -5692,
    34590 => -5695,
    34591 => -5698,
    34592 => -5701,
    34593 => -5704,
    34594 => -5707,
    34595 => -5710,
    34596 => -5713,
    34597 => -5716,
    34598 => -5719,
    34599 => -5723,
    34600 => -5726,
    34601 => -5729,
    34602 => -5732,
    34603 => -5735,
    34604 => -5738,
    34605 => -5741,
    34606 => -5744,
    34607 => -5747,
    34608 => -5750,
    34609 => -5754,
    34610 => -5757,
    34611 => -5760,
    34612 => -5763,
    34613 => -5766,
    34614 => -5769,
    34615 => -5772,
    34616 => -5775,
    34617 => -5778,
    34618 => -5781,
    34619 => -5784,
    34620 => -5788,
    34621 => -5791,
    34622 => -5794,
    34623 => -5797,
    34624 => -5800,
    34625 => -5803,
    34626 => -5806,
    34627 => -5809,
    34628 => -5812,
    34629 => -5815,
    34630 => -5818,
    34631 => -5822,
    34632 => -5825,
    34633 => -5828,
    34634 => -5831,
    34635 => -5834,
    34636 => -5837,
    34637 => -5840,
    34638 => -5843,
    34639 => -5846,
    34640 => -5849,
    34641 => -5852,
    34642 => -5856,
    34643 => -5859,
    34644 => -5862,
    34645 => -5865,
    34646 => -5868,
    34647 => -5871,
    34648 => -5874,
    34649 => -5877,
    34650 => -5880,
    34651 => -5883,
    34652 => -5886,
    34653 => -5890,
    34654 => -5893,
    34655 => -5896,
    34656 => -5899,
    34657 => -5902,
    34658 => -5905,
    34659 => -5908,
    34660 => -5911,
    34661 => -5914,
    34662 => -5917,
    34663 => -5920,
    34664 => -5924,
    34665 => -5927,
    34666 => -5930,
    34667 => -5933,
    34668 => -5936,
    34669 => -5939,
    34670 => -5942,
    34671 => -5945,
    34672 => -5948,
    34673 => -5951,
    34674 => -5954,
    34675 => -5958,
    34676 => -5961,
    34677 => -5964,
    34678 => -5967,
    34679 => -5970,
    34680 => -5973,
    34681 => -5976,
    34682 => -5979,
    34683 => -5982,
    34684 => -5985,
    34685 => -5988,
    34686 => -5991,
    34687 => -5995,
    34688 => -5998,
    34689 => -6001,
    34690 => -6004,
    34691 => -6007,
    34692 => -6010,
    34693 => -6013,
    34694 => -6016,
    34695 => -6019,
    34696 => -6022,
    34697 => -6025,
    34698 => -6029,
    34699 => -6032,
    34700 => -6035,
    34701 => -6038,
    34702 => -6041,
    34703 => -6044,
    34704 => -6047,
    34705 => -6050,
    34706 => -6053,
    34707 => -6056,
    34708 => -6059,
    34709 => -6063,
    34710 => -6066,
    34711 => -6069,
    34712 => -6072,
    34713 => -6075,
    34714 => -6078,
    34715 => -6081,
    34716 => -6084,
    34717 => -6087,
    34718 => -6090,
    34719 => -6093,
    34720 => -6096,
    34721 => -6100,
    34722 => -6103,
    34723 => -6106,
    34724 => -6109,
    34725 => -6112,
    34726 => -6115,
    34727 => -6118,
    34728 => -6121,
    34729 => -6124,
    34730 => -6127,
    34731 => -6130,
    34732 => -6134,
    34733 => -6137,
    34734 => -6140,
    34735 => -6143,
    34736 => -6146,
    34737 => -6149,
    34738 => -6152,
    34739 => -6155,
    34740 => -6158,
    34741 => -6161,
    34742 => -6164,
    34743 => -6167,
    34744 => -6171,
    34745 => -6174,
    34746 => -6177,
    34747 => -6180,
    34748 => -6183,
    34749 => -6186,
    34750 => -6189,
    34751 => -6192,
    34752 => -6195,
    34753 => -6198,
    34754 => -6201,
    34755 => -6204,
    34756 => -6208,
    34757 => -6211,
    34758 => -6214,
    34759 => -6217,
    34760 => -6220,
    34761 => -6223,
    34762 => -6226,
    34763 => -6229,
    34764 => -6232,
    34765 => -6235,
    34766 => -6238,
    34767 => -6241,
    34768 => -6245,
    34769 => -6248,
    34770 => -6251,
    34771 => -6254,
    34772 => -6257,
    34773 => -6260,
    34774 => -6263,
    34775 => -6266,
    34776 => -6269,
    34777 => -6272,
    34778 => -6275,
    34779 => -6278,
    34780 => -6282,
    34781 => -6285,
    34782 => -6288,
    34783 => -6291,
    34784 => -6294,
    34785 => -6297,
    34786 => -6300,
    34787 => -6303,
    34788 => -6306,
    34789 => -6309,
    34790 => -6312,
    34791 => -6315,
    34792 => -6319,
    34793 => -6322,
    34794 => -6325,
    34795 => -6328,
    34796 => -6331,
    34797 => -6334,
    34798 => -6337,
    34799 => -6340,
    34800 => -6343,
    34801 => -6346,
    34802 => -6349,
    34803 => -6352,
    34804 => -6356,
    34805 => -6359,
    34806 => -6362,
    34807 => -6365,
    34808 => -6368,
    34809 => -6371,
    34810 => -6374,
    34811 => -6377,
    34812 => -6380,
    34813 => -6383,
    34814 => -6386,
    34815 => -6389,
    34816 => -6393,
    34817 => -6396,
    34818 => -6399,
    34819 => -6402,
    34820 => -6405,
    34821 => -6408,
    34822 => -6411,
    34823 => -6414,
    34824 => -6417,
    34825 => -6420,
    34826 => -6423,
    34827 => -6426,
    34828 => -6429,
    34829 => -6433,
    34830 => -6436,
    34831 => -6439,
    34832 => -6442,
    34833 => -6445,
    34834 => -6448,
    34835 => -6451,
    34836 => -6454,
    34837 => -6457,
    34838 => -6460,
    34839 => -6463,
    34840 => -6466,
    34841 => -6470,
    34842 => -6473,
    34843 => -6476,
    34844 => -6479,
    34845 => -6482,
    34846 => -6485,
    34847 => -6488,
    34848 => -6491,
    34849 => -6494,
    34850 => -6497,
    34851 => -6500,
    34852 => -6503,
    34853 => -6506,
    34854 => -6510,
    34855 => -6513,
    34856 => -6516,
    34857 => -6519,
    34858 => -6522,
    34859 => -6525,
    34860 => -6528,
    34861 => -6531,
    34862 => -6534,
    34863 => -6537,
    34864 => -6540,
    34865 => -6543,
    34866 => -6547,
    34867 => -6550,
    34868 => -6553,
    34869 => -6556,
    34870 => -6559,
    34871 => -6562,
    34872 => -6565,
    34873 => -6568,
    34874 => -6571,
    34875 => -6574,
    34876 => -6577,
    34877 => -6580,
    34878 => -6583,
    34879 => -6587,
    34880 => -6590,
    34881 => -6593,
    34882 => -6596,
    34883 => -6599,
    34884 => -6602,
    34885 => -6605,
    34886 => -6608,
    34887 => -6611,
    34888 => -6614,
    34889 => -6617,
    34890 => -6620,
    34891 => -6623,
    34892 => -6627,
    34893 => -6630,
    34894 => -6633,
    34895 => -6636,
    34896 => -6639,
    34897 => -6642,
    34898 => -6645,
    34899 => -6648,
    34900 => -6651,
    34901 => -6654,
    34902 => -6657,
    34903 => -6660,
    34904 => -6663,
    34905 => -6667,
    34906 => -6670,
    34907 => -6673,
    34908 => -6676,
    34909 => -6679,
    34910 => -6682,
    34911 => -6685,
    34912 => -6688,
    34913 => -6691,
    34914 => -6694,
    34915 => -6697,
    34916 => -6700,
    34917 => -6703,
    34918 => -6706,
    34919 => -6710,
    34920 => -6713,
    34921 => -6716,
    34922 => -6719,
    34923 => -6722,
    34924 => -6725,
    34925 => -6728,
    34926 => -6731,
    34927 => -6734,
    34928 => -6737,
    34929 => -6740,
    34930 => -6743,
    34931 => -6746,
    34932 => -6750,
    34933 => -6753,
    34934 => -6756,
    34935 => -6759,
    34936 => -6762,
    34937 => -6765,
    34938 => -6768,
    34939 => -6771,
    34940 => -6774,
    34941 => -6777,
    34942 => -6780,
    34943 => -6783,
    34944 => -6786,
    34945 => -6789,
    34946 => -6793,
    34947 => -6796,
    34948 => -6799,
    34949 => -6802,
    34950 => -6805,
    34951 => -6808,
    34952 => -6811,
    34953 => -6814,
    34954 => -6817,
    34955 => -6820,
    34956 => -6823,
    34957 => -6826,
    34958 => -6829,
    34959 => -6833,
    34960 => -6836,
    34961 => -6839,
    34962 => -6842,
    34963 => -6845,
    34964 => -6848,
    34965 => -6851,
    34966 => -6854,
    34967 => -6857,
    34968 => -6860,
    34969 => -6863,
    34970 => -6866,
    34971 => -6869,
    34972 => -6872,
    34973 => -6876,
    34974 => -6879,
    34975 => -6882,
    34976 => -6885,
    34977 => -6888,
    34978 => -6891,
    34979 => -6894,
    34980 => -6897,
    34981 => -6900,
    34982 => -6903,
    34983 => -6906,
    34984 => -6909,
    34985 => -6912,
    34986 => -6915,
    34987 => -6919,
    34988 => -6922,
    34989 => -6925,
    34990 => -6928,
    34991 => -6931,
    34992 => -6934,
    34993 => -6937,
    34994 => -6940,
    34995 => -6943,
    34996 => -6946,
    34997 => -6949,
    34998 => -6952,
    34999 => -6955,
    35000 => -6958,
    35001 => -6961,
    35002 => -6965,
    35003 => -6968,
    35004 => -6971,
    35005 => -6974,
    35006 => -6977,
    35007 => -6980,
    35008 => -6983,
    35009 => -6986,
    35010 => -6989,
    35011 => -6992,
    35012 => -6995,
    35013 => -6998,
    35014 => -7001,
    35015 => -7004,
    35016 => -7008,
    35017 => -7011,
    35018 => -7014,
    35019 => -7017,
    35020 => -7020,
    35021 => -7023,
    35022 => -7026,
    35023 => -7029,
    35024 => -7032,
    35025 => -7035,
    35026 => -7038,
    35027 => -7041,
    35028 => -7044,
    35029 => -7047,
    35030 => -7050,
    35031 => -7054,
    35032 => -7057,
    35033 => -7060,
    35034 => -7063,
    35035 => -7066,
    35036 => -7069,
    35037 => -7072,
    35038 => -7075,
    35039 => -7078,
    35040 => -7081,
    35041 => -7084,
    35042 => -7087,
    35043 => -7090,
    35044 => -7093,
    35045 => -7097,
    35046 => -7100,
    35047 => -7103,
    35048 => -7106,
    35049 => -7109,
    35050 => -7112,
    35051 => -7115,
    35052 => -7118,
    35053 => -7121,
    35054 => -7124,
    35055 => -7127,
    35056 => -7130,
    35057 => -7133,
    35058 => -7136,
    35059 => -7139,
    35060 => -7143,
    35061 => -7146,
    35062 => -7149,
    35063 => -7152,
    35064 => -7155,
    35065 => -7158,
    35066 => -7161,
    35067 => -7164,
    35068 => -7167,
    35069 => -7170,
    35070 => -7173,
    35071 => -7176,
    35072 => -7179,
    35073 => -7182,
    35074 => -7185,
    35075 => -7188,
    35076 => -7192,
    35077 => -7195,
    35078 => -7198,
    35079 => -7201,
    35080 => -7204,
    35081 => -7207,
    35082 => -7210,
    35083 => -7213,
    35084 => -7216,
    35085 => -7219,
    35086 => -7222,
    35087 => -7225,
    35088 => -7228,
    35089 => -7231,
    35090 => -7234,
    35091 => -7238,
    35092 => -7241,
    35093 => -7244,
    35094 => -7247,
    35095 => -7250,
    35096 => -7253,
    35097 => -7256,
    35098 => -7259,
    35099 => -7262,
    35100 => -7265,
    35101 => -7268,
    35102 => -7271,
    35103 => -7274,
    35104 => -7277,
    35105 => -7280,
    35106 => -7283,
    35107 => -7287,
    35108 => -7290,
    35109 => -7293,
    35110 => -7296,
    35111 => -7299,
    35112 => -7302,
    35113 => -7305,
    35114 => -7308,
    35115 => -7311,
    35116 => -7314,
    35117 => -7317,
    35118 => -7320,
    35119 => -7323,
    35120 => -7326,
    35121 => -7329,
    35122 => -7332,
    35123 => -7336,
    35124 => -7339,
    35125 => -7342,
    35126 => -7345,
    35127 => -7348,
    35128 => -7351,
    35129 => -7354,
    35130 => -7357,
    35131 => -7360,
    35132 => -7363,
    35133 => -7366,
    35134 => -7369,
    35135 => -7372,
    35136 => -7375,
    35137 => -7378,
    35138 => -7381,
    35139 => -7385,
    35140 => -7388,
    35141 => -7391,
    35142 => -7394,
    35143 => -7397,
    35144 => -7400,
    35145 => -7403,
    35146 => -7406,
    35147 => -7409,
    35148 => -7412,
    35149 => -7415,
    35150 => -7418,
    35151 => -7421,
    35152 => -7424,
    35153 => -7427,
    35154 => -7430,
    35155 => -7433,
    35156 => -7437,
    35157 => -7440,
    35158 => -7443,
    35159 => -7446,
    35160 => -7449,
    35161 => -7452,
    35162 => -7455,
    35163 => -7458,
    35164 => -7461,
    35165 => -7464,
    35166 => -7467,
    35167 => -7470,
    35168 => -7473,
    35169 => -7476,
    35170 => -7479,
    35171 => -7482,
    35172 => -7485,
    35173 => -7489,
    35174 => -7492,
    35175 => -7495,
    35176 => -7498,
    35177 => -7501,
    35178 => -7504,
    35179 => -7507,
    35180 => -7510,
    35181 => -7513,
    35182 => -7516,
    35183 => -7519,
    35184 => -7522,
    35185 => -7525,
    35186 => -7528,
    35187 => -7531,
    35188 => -7534,
    35189 => -7537,
    35190 => -7541,
    35191 => -7544,
    35192 => -7547,
    35193 => -7550,
    35194 => -7553,
    35195 => -7556,
    35196 => -7559,
    35197 => -7562,
    35198 => -7565,
    35199 => -7568,
    35200 => -7571,
    35201 => -7574,
    35202 => -7577,
    35203 => -7580,
    35204 => -7583,
    35205 => -7586,
    35206 => -7589,
    35207 => -7592,
    35208 => -7596,
    35209 => -7599,
    35210 => -7602,
    35211 => -7605,
    35212 => -7608,
    35213 => -7611,
    35214 => -7614,
    35215 => -7617,
    35216 => -7620,
    35217 => -7623,
    35218 => -7626,
    35219 => -7629,
    35220 => -7632,
    35221 => -7635,
    35222 => -7638,
    35223 => -7641,
    35224 => -7644,
    35225 => -7647,
    35226 => -7651,
    35227 => -7654,
    35228 => -7657,
    35229 => -7660,
    35230 => -7663,
    35231 => -7666,
    35232 => -7669,
    35233 => -7672,
    35234 => -7675,
    35235 => -7678,
    35236 => -7681,
    35237 => -7684,
    35238 => -7687,
    35239 => -7690,
    35240 => -7693,
    35241 => -7696,
    35242 => -7699,
    35243 => -7702,
    35244 => -7705,
    35245 => -7709,
    35246 => -7712,
    35247 => -7715,
    35248 => -7718,
    35249 => -7721,
    35250 => -7724,
    35251 => -7727,
    35252 => -7730,
    35253 => -7733,
    35254 => -7736,
    35255 => -7739,
    35256 => -7742,
    35257 => -7745,
    35258 => -7748,
    35259 => -7751,
    35260 => -7754,
    35261 => -7757,
    35262 => -7760,
    35263 => -7764,
    35264 => -7767,
    35265 => -7770,
    35266 => -7773,
    35267 => -7776,
    35268 => -7779,
    35269 => -7782,
    35270 => -7785,
    35271 => -7788,
    35272 => -7791,
    35273 => -7794,
    35274 => -7797,
    35275 => -7800,
    35276 => -7803,
    35277 => -7806,
    35278 => -7809,
    35279 => -7812,
    35280 => -7815,
    35281 => -7818,
    35282 => -7821,
    35283 => -7825,
    35284 => -7828,
    35285 => -7831,
    35286 => -7834,
    35287 => -7837,
    35288 => -7840,
    35289 => -7843,
    35290 => -7846,
    35291 => -7849,
    35292 => -7852,
    35293 => -7855,
    35294 => -7858,
    35295 => -7861,
    35296 => -7864,
    35297 => -7867,
    35298 => -7870,
    35299 => -7873,
    35300 => -7876,
    35301 => -7879,
    35302 => -7882,
    35303 => -7886,
    35304 => -7889,
    35305 => -7892,
    35306 => -7895,
    35307 => -7898,
    35308 => -7901,
    35309 => -7904,
    35310 => -7907,
    35311 => -7910,
    35312 => -7913,
    35313 => -7916,
    35314 => -7919,
    35315 => -7922,
    35316 => -7925,
    35317 => -7928,
    35318 => -7931,
    35319 => -7934,
    35320 => -7937,
    35321 => -7940,
    35322 => -7943,
    35323 => -7946,
    35324 => -7950,
    35325 => -7953,
    35326 => -7956,
    35327 => -7959,
    35328 => -7962,
    35329 => -7965,
    35330 => -7968,
    35331 => -7971,
    35332 => -7974,
    35333 => -7977,
    35334 => -7980,
    35335 => -7983,
    35336 => -7986,
    35337 => -7989,
    35338 => -7992,
    35339 => -7995,
    35340 => -7998,
    35341 => -8001,
    35342 => -8004,
    35343 => -8007,
    35344 => -8010,
    35345 => -8014,
    35346 => -8017,
    35347 => -8020,
    35348 => -8023,
    35349 => -8026,
    35350 => -8029,
    35351 => -8032,
    35352 => -8035,
    35353 => -8038,
    35354 => -8041,
    35355 => -8044,
    35356 => -8047,
    35357 => -8050,
    35358 => -8053,
    35359 => -8056,
    35360 => -8059,
    35361 => -8062,
    35362 => -8065,
    35363 => -8068,
    35364 => -8071,
    35365 => -8074,
    35366 => -8077,
    35367 => -8081,
    35368 => -8084,
    35369 => -8087,
    35370 => -8090,
    35371 => -8093,
    35372 => -8096,
    35373 => -8099,
    35374 => -8102,
    35375 => -8105,
    35376 => -8108,
    35377 => -8111,
    35378 => -8114,
    35379 => -8117,
    35380 => -8120,
    35381 => -8123,
    35382 => -8126,
    35383 => -8129,
    35384 => -8132,
    35385 => -8135,
    35386 => -8138,
    35387 => -8141,
    35388 => -8144,
    35389 => -8147,
    35390 => -8151,
    35391 => -8154,
    35392 => -8157,
    35393 => -8160,
    35394 => -8163,
    35395 => -8166,
    35396 => -8169,
    35397 => -8172,
    35398 => -8175,
    35399 => -8178,
    35400 => -8181,
    35401 => -8184,
    35402 => -8187,
    35403 => -8190,
    35404 => -8193,
    35405 => -8196,
    35406 => -8199,
    35407 => -8202,
    35408 => -8205,
    35409 => -8208,
    35410 => -8211,
    35411 => -8214,
    35412 => -8217,
    35413 => -8220,
    35414 => -8224,
    35415 => -8227,
    35416 => -8230,
    35417 => -8233,
    35418 => -8236,
    35419 => -8239,
    35420 => -8242,
    35421 => -8245,
    35422 => -8248,
    35423 => -8251,
    35424 => -8254,
    35425 => -8257,
    35426 => -8260,
    35427 => -8263,
    35428 => -8266,
    35429 => -8269,
    35430 => -8272,
    35431 => -8275,
    35432 => -8278,
    35433 => -8281,
    35434 => -8284,
    35435 => -8287,
    35436 => -8290,
    35437 => -8293,
    35438 => -8296,
    35439 => -8300,
    35440 => -8303,
    35441 => -8306,
    35442 => -8309,
    35443 => -8312,
    35444 => -8315,
    35445 => -8318,
    35446 => -8321,
    35447 => -8324,
    35448 => -8327,
    35449 => -8330,
    35450 => -8333,
    35451 => -8336,
    35452 => -8339,
    35453 => -8342,
    35454 => -8345,
    35455 => -8348,
    35456 => -8351,
    35457 => -8354,
    35458 => -8357,
    35459 => -8360,
    35460 => -8363,
    35461 => -8366,
    35462 => -8369,
    35463 => -8372,
    35464 => -8375,
    35465 => -8379,
    35466 => -8382,
    35467 => -8385,
    35468 => -8388,
    35469 => -8391,
    35470 => -8394,
    35471 => -8397,
    35472 => -8400,
    35473 => -8403,
    35474 => -8406,
    35475 => -8409,
    35476 => -8412,
    35477 => -8415,
    35478 => -8418,
    35479 => -8421,
    35480 => -8424,
    35481 => -8427,
    35482 => -8430,
    35483 => -8433,
    35484 => -8436,
    35485 => -8439,
    35486 => -8442,
    35487 => -8445,
    35488 => -8448,
    35489 => -8451,
    35490 => -8454,
    35491 => -8457,
    35492 => -8460,
    35493 => -8464,
    35494 => -8467,
    35495 => -8470,
    35496 => -8473,
    35497 => -8476,
    35498 => -8479,
    35499 => -8482,
    35500 => -8485,
    35501 => -8488,
    35502 => -8491,
    35503 => -8494,
    35504 => -8497,
    35505 => -8500,
    35506 => -8503,
    35507 => -8506,
    35508 => -8509,
    35509 => -8512,
    35510 => -8515,
    35511 => -8518,
    35512 => -8521,
    35513 => -8524,
    35514 => -8527,
    35515 => -8530,
    35516 => -8533,
    35517 => -8536,
    35518 => -8539,
    35519 => -8542,
    35520 => -8545,
    35521 => -8548,
    35522 => -8552,
    35523 => -8555,
    35524 => -8558,
    35525 => -8561,
    35526 => -8564,
    35527 => -8567,
    35528 => -8570,
    35529 => -8573,
    35530 => -8576,
    35531 => -8579,
    35532 => -8582,
    35533 => -8585,
    35534 => -8588,
    35535 => -8591,
    35536 => -8594,
    35537 => -8597,
    35538 => -8600,
    35539 => -8603,
    35540 => -8606,
    35541 => -8609,
    35542 => -8612,
    35543 => -8615,
    35544 => -8618,
    35545 => -8621,
    35546 => -8624,
    35547 => -8627,
    35548 => -8630,
    35549 => -8633,
    35550 => -8636,
    35551 => -8639,
    35552 => -8642,
    35553 => -8645,
    35554 => -8649,
    35555 => -8652,
    35556 => -8655,
    35557 => -8658,
    35558 => -8661,
    35559 => -8664,
    35560 => -8667,
    35561 => -8670,
    35562 => -8673,
    35563 => -8676,
    35564 => -8679,
    35565 => -8682,
    35566 => -8685,
    35567 => -8688,
    35568 => -8691,
    35569 => -8694,
    35570 => -8697,
    35571 => -8700,
    35572 => -8703,
    35573 => -8706,
    35574 => -8709,
    35575 => -8712,
    35576 => -8715,
    35577 => -8718,
    35578 => -8721,
    35579 => -8724,
    35580 => -8727,
    35581 => -8730,
    35582 => -8733,
    35583 => -8736,
    35584 => -8739,
    35585 => -8742,
    35586 => -8745,
    35587 => -8748,
    35588 => -8751,
    35589 => -8755,
    35590 => -8758,
    35591 => -8761,
    35592 => -8764,
    35593 => -8767,
    35594 => -8770,
    35595 => -8773,
    35596 => -8776,
    35597 => -8779,
    35598 => -8782,
    35599 => -8785,
    35600 => -8788,
    35601 => -8791,
    35602 => -8794,
    35603 => -8797,
    35604 => -8800,
    35605 => -8803,
    35606 => -8806,
    35607 => -8809,
    35608 => -8812,
    35609 => -8815,
    35610 => -8818,
    35611 => -8821,
    35612 => -8824,
    35613 => -8827,
    35614 => -8830,
    35615 => -8833,
    35616 => -8836,
    35617 => -8839,
    35618 => -8842,
    35619 => -8845,
    35620 => -8848,
    35621 => -8851,
    35622 => -8854,
    35623 => -8857,
    35624 => -8860,
    35625 => -8863,
    35626 => -8866,
    35627 => -8869,
    35628 => -8873,
    35629 => -8876,
    35630 => -8879,
    35631 => -8882,
    35632 => -8885,
    35633 => -8888,
    35634 => -8891,
    35635 => -8894,
    35636 => -8897,
    35637 => -8900,
    35638 => -8903,
    35639 => -8906,
    35640 => -8909,
    35641 => -8912,
    35642 => -8915,
    35643 => -8918,
    35644 => -8921,
    35645 => -8924,
    35646 => -8927,
    35647 => -8930,
    35648 => -8933,
    35649 => -8936,
    35650 => -8939,
    35651 => -8942,
    35652 => -8945,
    35653 => -8948,
    35654 => -8951,
    35655 => -8954,
    35656 => -8957,
    35657 => -8960,
    35658 => -8963,
    35659 => -8966,
    35660 => -8969,
    35661 => -8972,
    35662 => -8975,
    35663 => -8978,
    35664 => -8981,
    35665 => -8984,
    35666 => -8987,
    35667 => -8990,
    35668 => -8993,
    35669 => -8996,
    35670 => -8999,
    35671 => -9002,
    35672 => -9006,
    35673 => -9009,
    35674 => -9012,
    35675 => -9015,
    35676 => -9018,
    35677 => -9021,
    35678 => -9024,
    35679 => -9027,
    35680 => -9030,
    35681 => -9033,
    35682 => -9036,
    35683 => -9039,
    35684 => -9042,
    35685 => -9045,
    35686 => -9048,
    35687 => -9051,
    35688 => -9054,
    35689 => -9057,
    35690 => -9060,
    35691 => -9063,
    35692 => -9066,
    35693 => -9069,
    35694 => -9072,
    35695 => -9075,
    35696 => -9078,
    35697 => -9081,
    35698 => -9084,
    35699 => -9087,
    35700 => -9090,
    35701 => -9093,
    35702 => -9096,
    35703 => -9099,
    35704 => -9102,
    35705 => -9105,
    35706 => -9108,
    35707 => -9111,
    35708 => -9114,
    35709 => -9117,
    35710 => -9120,
    35711 => -9123,
    35712 => -9126,
    35713 => -9129,
    35714 => -9132,
    35715 => -9135,
    35716 => -9138,
    35717 => -9141,
    35718 => -9144,
    35719 => -9147,
    35720 => -9150,
    35721 => -9153,
    35722 => -9156,
    35723 => -9159,
    35724 => -9162,
    35725 => -9165,
    35726 => -9168,
    35727 => -9172,
    35728 => -9175,
    35729 => -9178,
    35730 => -9181,
    35731 => -9184,
    35732 => -9187,
    35733 => -9190,
    35734 => -9193,
    35735 => -9196,
    35736 => -9199,
    35737 => -9202,
    35738 => -9205,
    35739 => -9208,
    35740 => -9211,
    35741 => -9214,
    35742 => -9217,
    35743 => -9220,
    35744 => -9223,
    35745 => -9226,
    35746 => -9229,
    35747 => -9232,
    35748 => -9235,
    35749 => -9238,
    35750 => -9241,
    35751 => -9244,
    35752 => -9247,
    35753 => -9250,
    35754 => -9253,
    35755 => -9256,
    35756 => -9259,
    35757 => -9262,
    35758 => -9265,
    35759 => -9268,
    35760 => -9271,
    35761 => -9274,
    35762 => -9277,
    35763 => -9280,
    35764 => -9283,
    35765 => -9286,
    35766 => -9289,
    35767 => -9292,
    35768 => -9295,
    35769 => -9298,
    35770 => -9301,
    35771 => -9304,
    35772 => -9307,
    35773 => -9310,
    35774 => -9313,
    35775 => -9316,
    35776 => -9319,
    35777 => -9322,
    35778 => -9325,
    35779 => -9328,
    35780 => -9331,
    35781 => -9334,
    35782 => -9337,
    35783 => -9340,
    35784 => -9343,
    35785 => -9346,
    35786 => -9349,
    35787 => -9352,
    35788 => -9355,
    35789 => -9358,
    35790 => -9361,
    35791 => -9364,
    35792 => -9367,
    35793 => -9370,
    35794 => -9373,
    35795 => -9376,
    35796 => -9379,
    35797 => -9382,
    35798 => -9385,
    35799 => -9388,
    35800 => -9391,
    35801 => -9394,
    35802 => -9397,
    35803 => -9400,
    35804 => -9403,
    35805 => -9406,
    35806 => -9409,
    35807 => -9413,
    35808 => -9416,
    35809 => -9419,
    35810 => -9422,
    35811 => -9425,
    35812 => -9428,
    35813 => -9431,
    35814 => -9434,
    35815 => -9437,
    35816 => -9440,
    35817 => -9443,
    35818 => -9446,
    35819 => -9449,
    35820 => -9452,
    35821 => -9455,
    35822 => -9458,
    35823 => -9461,
    35824 => -9464,
    35825 => -9467,
    35826 => -9470,
    35827 => -9473,
    35828 => -9476,
    35829 => -9479,
    35830 => -9482,
    35831 => -9485,
    35832 => -9488,
    35833 => -9491,
    35834 => -9494,
    35835 => -9497,
    35836 => -9500,
    35837 => -9503,
    35838 => -9506,
    35839 => -9509,
    35840 => -9512,
    35841 => -9515,
    35842 => -9518,
    35843 => -9521,
    35844 => -9524,
    35845 => -9527,
    35846 => -9530,
    35847 => -9533,
    35848 => -9536,
    35849 => -9539,
    35850 => -9542,
    35851 => -9545,
    35852 => -9548,
    35853 => -9551,
    35854 => -9554,
    35855 => -9557,
    35856 => -9560,
    35857 => -9563,
    35858 => -9566,
    35859 => -9569,
    35860 => -9572,
    35861 => -9575,
    35862 => -9578,
    35863 => -9581,
    35864 => -9584,
    35865 => -9587,
    35866 => -9590,
    35867 => -9593,
    35868 => -9596,
    35869 => -9599,
    35870 => -9602,
    35871 => -9605,
    35872 => -9608,
    35873 => -9611,
    35874 => -9614,
    35875 => -9617,
    35876 => -9620,
    35877 => -9623,
    35878 => -9626,
    35879 => -9629,
    35880 => -9632,
    35881 => -9635,
    35882 => -9638,
    35883 => -9641,
    35884 => -9644,
    35885 => -9647,
    35886 => -9650,
    35887 => -9653,
    35888 => -9656,
    35889 => -9659,
    35890 => -9662,
    35891 => -9665,
    35892 => -9668,
    35893 => -9671,
    35894 => -9674,
    35895 => -9677,
    35896 => -9680,
    35897 => -9683,
    35898 => -9686,
    35899 => -9689,
    35900 => -9692,
    35901 => -9695,
    35902 => -9698,
    35903 => -9701,
    35904 => -9704,
    35905 => -9707,
    35906 => -9710,
    35907 => -9713,
    35908 => -9716,
    35909 => -9719,
    35910 => -9722,
    35911 => -9725,
    35912 => -9728,
    35913 => -9731,
    35914 => -9734,
    35915 => -9737,
    35916 => -9740,
    35917 => -9743,
    35918 => -9746,
    35919 => -9749,
    35920 => -9752,
    35921 => -9755,
    35922 => -9758,
    35923 => -9761,
    35924 => -9764,
    35925 => -9767,
    35926 => -9770,
    35927 => -9773,
    35928 => -9776,
    35929 => -9779,
    35930 => -9782,
    35931 => -9785,
    35932 => -9788,
    35933 => -9791,
    35934 => -9794,
    35935 => -9797,
    35936 => -9800,
    35937 => -9803,
    35938 => -9806,
    35939 => -9809,
    35940 => -9812,
    35941 => -9815,
    35942 => -9818,
    35943 => -9821,
    35944 => -9824,
    35945 => -9827,
    35946 => -9830,
    35947 => -9833,
    35948 => -9836,
    35949 => -9839,
    35950 => -9842,
    35951 => -9845,
    35952 => -9848,
    35953 => -9851,
    35954 => -9854,
    35955 => -9857,
    35956 => -9860,
    35957 => -9863,
    35958 => -9866,
    35959 => -9869,
    35960 => -9872,
    35961 => -9875,
    35962 => -9878,
    35963 => -9881,
    35964 => -9884,
    35965 => -9887,
    35966 => -9890,
    35967 => -9893,
    35968 => -9896,
    35969 => -9899,
    35970 => -9902,
    35971 => -9905,
    35972 => -9908,
    35973 => -9911,
    35974 => -9914,
    35975 => -9917,
    35976 => -9920,
    35977 => -9923,
    35978 => -9926,
    35979 => -9929,
    35980 => -9932,
    35981 => -9935,
    35982 => -9938,
    35983 => -9941,
    35984 => -9944,
    35985 => -9947,
    35986 => -9950,
    35987 => -9953,
    35988 => -9956,
    35989 => -9959,
    35990 => -9962,
    35991 => -9965,
    35992 => -9968,
    35993 => -9971,
    35994 => -9974,
    35995 => -9977,
    35996 => -9980,
    35997 => -9983,
    35998 => -9986,
    35999 => -9989,
    36000 => -9992,
    36001 => -9995,
    36002 => -9998,
    36003 => -10001,
    36004 => -10004,
    36005 => -10007,
    36006 => -10010,
    36007 => -10013,
    36008 => -10016,
    36009 => -10019,
    36010 => -10022,
    36011 => -10025,
    36012 => -10028,
    36013 => -10031,
    36014 => -10033,
    36015 => -10036,
    36016 => -10039,
    36017 => -10042,
    36018 => -10045,
    36019 => -10048,
    36020 => -10051,
    36021 => -10054,
    36022 => -10057,
    36023 => -10060,
    36024 => -10063,
    36025 => -10066,
    36026 => -10069,
    36027 => -10072,
    36028 => -10075,
    36029 => -10078,
    36030 => -10081,
    36031 => -10084,
    36032 => -10087,
    36033 => -10090,
    36034 => -10093,
    36035 => -10096,
    36036 => -10099,
    36037 => -10102,
    36038 => -10105,
    36039 => -10108,
    36040 => -10111,
    36041 => -10114,
    36042 => -10117,
    36043 => -10120,
    36044 => -10123,
    36045 => -10126,
    36046 => -10129,
    36047 => -10132,
    36048 => -10135,
    36049 => -10138,
    36050 => -10141,
    36051 => -10144,
    36052 => -10147,
    36053 => -10150,
    36054 => -10153,
    36055 => -10156,
    36056 => -10159,
    36057 => -10162,
    36058 => -10165,
    36059 => -10168,
    36060 => -10171,
    36061 => -10174,
    36062 => -10177,
    36063 => -10180,
    36064 => -10183,
    36065 => -10186,
    36066 => -10189,
    36067 => -10192,
    36068 => -10195,
    36069 => -10198,
    36070 => -10201,
    36071 => -10204,
    36072 => -10207,
    36073 => -10210,
    36074 => -10213,
    36075 => -10216,
    36076 => -10219,
    36077 => -10222,
    36078 => -10225,
    36079 => -10228,
    36080 => -10231,
    36081 => -10234,
    36082 => -10237,
    36083 => -10240,
    36084 => -10243,
    36085 => -10246,
    36086 => -10249,
    36087 => -10252,
    36088 => -10255,
    36089 => -10258,
    36090 => -10261,
    36091 => -10263,
    36092 => -10266,
    36093 => -10269,
    36094 => -10272,
    36095 => -10275,
    36096 => -10278,
    36097 => -10281,
    36098 => -10284,
    36099 => -10287,
    36100 => -10290,
    36101 => -10293,
    36102 => -10296,
    36103 => -10299,
    36104 => -10302,
    36105 => -10305,
    36106 => -10308,
    36107 => -10311,
    36108 => -10314,
    36109 => -10317,
    36110 => -10320,
    36111 => -10323,
    36112 => -10326,
    36113 => -10329,
    36114 => -10332,
    36115 => -10335,
    36116 => -10338,
    36117 => -10341,
    36118 => -10344,
    36119 => -10347,
    36120 => -10350,
    36121 => -10353,
    36122 => -10356,
    36123 => -10359,
    36124 => -10362,
    36125 => -10365,
    36126 => -10368,
    36127 => -10371,
    36128 => -10374,
    36129 => -10377,
    36130 => -10380,
    36131 => -10383,
    36132 => -10386,
    36133 => -10389,
    36134 => -10392,
    36135 => -10395,
    36136 => -10398,
    36137 => -10401,
    36138 => -10404,
    36139 => -10407,
    36140 => -10410,
    36141 => -10413,
    36142 => -10416,
    36143 => -10419,
    36144 => -10421,
    36145 => -10424,
    36146 => -10427,
    36147 => -10430,
    36148 => -10433,
    36149 => -10436,
    36150 => -10439,
    36151 => -10442,
    36152 => -10445,
    36153 => -10448,
    36154 => -10451,
    36155 => -10454,
    36156 => -10457,
    36157 => -10460,
    36158 => -10463,
    36159 => -10466,
    36160 => -10469,
    36161 => -10472,
    36162 => -10475,
    36163 => -10478,
    36164 => -10481,
    36165 => -10484,
    36166 => -10487,
    36167 => -10490,
    36168 => -10493,
    36169 => -10496,
    36170 => -10499,
    36171 => -10502,
    36172 => -10505,
    36173 => -10508,
    36174 => -10511,
    36175 => -10514,
    36176 => -10517,
    36177 => -10520,
    36178 => -10523,
    36179 => -10526,
    36180 => -10529,
    36181 => -10532,
    36182 => -10535,
    36183 => -10538,
    36184 => -10541,
    36185 => -10544,
    36186 => -10546,
    36187 => -10549,
    36188 => -10552,
    36189 => -10555,
    36190 => -10558,
    36191 => -10561,
    36192 => -10564,
    36193 => -10567,
    36194 => -10570,
    36195 => -10573,
    36196 => -10576,
    36197 => -10579,
    36198 => -10582,
    36199 => -10585,
    36200 => -10588,
    36201 => -10591,
    36202 => -10594,
    36203 => -10597,
    36204 => -10600,
    36205 => -10603,
    36206 => -10606,
    36207 => -10609,
    36208 => -10612,
    36209 => -10615,
    36210 => -10618,
    36211 => -10621,
    36212 => -10624,
    36213 => -10627,
    36214 => -10630,
    36215 => -10633,
    36216 => -10636,
    36217 => -10639,
    36218 => -10642,
    36219 => -10645,
    36220 => -10648,
    36221 => -10651,
    36222 => -10654,
    36223 => -10656,
    36224 => -10659,
    36225 => -10662,
    36226 => -10665,
    36227 => -10668,
    36228 => -10671,
    36229 => -10674,
    36230 => -10677,
    36231 => -10680,
    36232 => -10683,
    36233 => -10686,
    36234 => -10689,
    36235 => -10692,
    36236 => -10695,
    36237 => -10698,
    36238 => -10701,
    36239 => -10704,
    36240 => -10707,
    36241 => -10710,
    36242 => -10713,
    36243 => -10716,
    36244 => -10719,
    36245 => -10722,
    36246 => -10725,
    36247 => -10728,
    36248 => -10731,
    36249 => -10734,
    36250 => -10737,
    36251 => -10740,
    36252 => -10743,
    36253 => -10746,
    36254 => -10749,
    36255 => -10751,
    36256 => -10754,
    36257 => -10757,
    36258 => -10760,
    36259 => -10763,
    36260 => -10766,
    36261 => -10769,
    36262 => -10772,
    36263 => -10775,
    36264 => -10778,
    36265 => -10781,
    36266 => -10784,
    36267 => -10787,
    36268 => -10790,
    36269 => -10793,
    36270 => -10796,
    36271 => -10799,
    36272 => -10802,
    36273 => -10805,
    36274 => -10808,
    36275 => -10811,
    36276 => -10814,
    36277 => -10817,
    36278 => -10820,
    36279 => -10823,
    36280 => -10826,
    36281 => -10829,
    36282 => -10832,
    36283 => -10835,
    36284 => -10838,
    36285 => -10840,
    36286 => -10843,
    36287 => -10846,
    36288 => -10849,
    36289 => -10852,
    36290 => -10855,
    36291 => -10858,
    36292 => -10861,
    36293 => -10864,
    36294 => -10867,
    36295 => -10870,
    36296 => -10873,
    36297 => -10876,
    36298 => -10879,
    36299 => -10882,
    36300 => -10885,
    36301 => -10888,
    36302 => -10891,
    36303 => -10894,
    36304 => -10897,
    36305 => -10900,
    36306 => -10903,
    36307 => -10906,
    36308 => -10909,
    36309 => -10912,
    36310 => -10915,
    36311 => -10918,
    36312 => -10920,
    36313 => -10923,
    36314 => -10926,
    36315 => -10929,
    36316 => -10932,
    36317 => -10935,
    36318 => -10938,
    36319 => -10941,
    36320 => -10944,
    36321 => -10947,
    36322 => -10950,
    36323 => -10953,
    36324 => -10956,
    36325 => -10959,
    36326 => -10962,
    36327 => -10965,
    36328 => -10968,
    36329 => -10971,
    36330 => -10974,
    36331 => -10977,
    36332 => -10980,
    36333 => -10983,
    36334 => -10986,
    36335 => -10989,
    36336 => -10992,
    36337 => -10994,
    36338 => -10997,
    36339 => -11000,
    36340 => -11003,
    36341 => -11006,
    36342 => -11009,
    36343 => -11012,
    36344 => -11015,
    36345 => -11018,
    36346 => -11021,
    36347 => -11024,
    36348 => -11027,
    36349 => -11030,
    36350 => -11033,
    36351 => -11036,
    36352 => -11039,
    36353 => -11042,
    36354 => -11045,
    36355 => -11048,
    36356 => -11051,
    36357 => -11054,
    36358 => -11057,
    36359 => -11060,
    36360 => -11063,
    36361 => -11065,
    36362 => -11068,
    36363 => -11071,
    36364 => -11074,
    36365 => -11077,
    36366 => -11080,
    36367 => -11083,
    36368 => -11086,
    36369 => -11089,
    36370 => -11092,
    36371 => -11095,
    36372 => -11098,
    36373 => -11101,
    36374 => -11104,
    36375 => -11107,
    36376 => -11110,
    36377 => -11113,
    36378 => -11116,
    36379 => -11119,
    36380 => -11122,
    36381 => -11125,
    36382 => -11128,
    36383 => -11131,
    36384 => -11133,
    36385 => -11136,
    36386 => -11139,
    36387 => -11142,
    36388 => -11145,
    36389 => -11148,
    36390 => -11151,
    36391 => -11154,
    36392 => -11157,
    36393 => -11160,
    36394 => -11163,
    36395 => -11166,
    36396 => -11169,
    36397 => -11172,
    36398 => -11175,
    36399 => -11178,
    36400 => -11181,
    36401 => -11184,
    36402 => -11187,
    36403 => -11190,
    36404 => -11193,
    36405 => -11195,
    36406 => -11198,
    36407 => -11201,
    36408 => -11204,
    36409 => -11207,
    36410 => -11210,
    36411 => -11213,
    36412 => -11216,
    36413 => -11219,
    36414 => -11222,
    36415 => -11225,
    36416 => -11228,
    36417 => -11231,
    36418 => -11234,
    36419 => -11237,
    36420 => -11240,
    36421 => -11243,
    36422 => -11246,
    36423 => -11249,
    36424 => -11252,
    36425 => -11255,
    36426 => -11257,
    36427 => -11260,
    36428 => -11263,
    36429 => -11266,
    36430 => -11269,
    36431 => -11272,
    36432 => -11275,
    36433 => -11278,
    36434 => -11281,
    36435 => -11284,
    36436 => -11287,
    36437 => -11290,
    36438 => -11293,
    36439 => -11296,
    36440 => -11299,
    36441 => -11302,
    36442 => -11305,
    36443 => -11308,
    36444 => -11311,
    36445 => -11314,
    36446 => -11316,
    36447 => -11319,
    36448 => -11322,
    36449 => -11325,
    36450 => -11328,
    36451 => -11331,
    36452 => -11334,
    36453 => -11337,
    36454 => -11340,
    36455 => -11343,
    36456 => -11346,
    36457 => -11349,
    36458 => -11352,
    36459 => -11355,
    36460 => -11358,
    36461 => -11361,
    36462 => -11364,
    36463 => -11367,
    36464 => -11370,
    36465 => -11372,
    36466 => -11375,
    36467 => -11378,
    36468 => -11381,
    36469 => -11384,
    36470 => -11387,
    36471 => -11390,
    36472 => -11393,
    36473 => -11396,
    36474 => -11399,
    36475 => -11402,
    36476 => -11405,
    36477 => -11408,
    36478 => -11411,
    36479 => -11414,
    36480 => -11417,
    36481 => -11420,
    36482 => -11423,
    36483 => -11425,
    36484 => -11428,
    36485 => -11431,
    36486 => -11434,
    36487 => -11437,
    36488 => -11440,
    36489 => -11443,
    36490 => -11446,
    36491 => -11449,
    36492 => -11452,
    36493 => -11455,
    36494 => -11458,
    36495 => -11461,
    36496 => -11464,
    36497 => -11467,
    36498 => -11470,
    36499 => -11473,
    36500 => -11476,
    36501 => -11478,
    36502 => -11481,
    36503 => -11484,
    36504 => -11487,
    36505 => -11490,
    36506 => -11493,
    36507 => -11496,
    36508 => -11499,
    36509 => -11502,
    36510 => -11505,
    36511 => -11508,
    36512 => -11511,
    36513 => -11514,
    36514 => -11517,
    36515 => -11520,
    36516 => -11523,
    36517 => -11526,
    36518 => -11528,
    36519 => -11531,
    36520 => -11534,
    36521 => -11537,
    36522 => -11540,
    36523 => -11543,
    36524 => -11546,
    36525 => -11549,
    36526 => -11552,
    36527 => -11555,
    36528 => -11558,
    36529 => -11561,
    36530 => -11564,
    36531 => -11567,
    36532 => -11570,
    36533 => -11573,
    36534 => -11575,
    36535 => -11578,
    36536 => -11581,
    36537 => -11584,
    36538 => -11587,
    36539 => -11590,
    36540 => -11593,
    36541 => -11596,
    36542 => -11599,
    36543 => -11602,
    36544 => -11605,
    36545 => -11608,
    36546 => -11611,
    36547 => -11614,
    36548 => -11617,
    36549 => -11620,
    36550 => -11623,
    36551 => -11625,
    36552 => -11628,
    36553 => -11631,
    36554 => -11634,
    36555 => -11637,
    36556 => -11640,
    36557 => -11643,
    36558 => -11646,
    36559 => -11649,
    36560 => -11652,
    36561 => -11655,
    36562 => -11658,
    36563 => -11661,
    36564 => -11664,
    36565 => -11667,
    36566 => -11669,
    36567 => -11672,
    36568 => -11675,
    36569 => -11678,
    36570 => -11681,
    36571 => -11684,
    36572 => -11687,
    36573 => -11690,
    36574 => -11693,
    36575 => -11696,
    36576 => -11699,
    36577 => -11702,
    36578 => -11705,
    36579 => -11708,
    36580 => -11711,
    36581 => -11714,
    36582 => -11716,
    36583 => -11719,
    36584 => -11722,
    36585 => -11725,
    36586 => -11728,
    36587 => -11731,
    36588 => -11734,
    36589 => -11737,
    36590 => -11740,
    36591 => -11743,
    36592 => -11746,
    36593 => -11749,
    36594 => -11752,
    36595 => -11755,
    36596 => -11758,
    36597 => -11760,
    36598 => -11763,
    36599 => -11766,
    36600 => -11769,
    36601 => -11772,
    36602 => -11775,
    36603 => -11778,
    36604 => -11781,
    36605 => -11784,
    36606 => -11787,
    36607 => -11790,
    36608 => -11793,
    36609 => -11796,
    36610 => -11799,
    36611 => -11801,
    36612 => -11804,
    36613 => -11807,
    36614 => -11810,
    36615 => -11813,
    36616 => -11816,
    36617 => -11819,
    36618 => -11822,
    36619 => -11825,
    36620 => -11828,
    36621 => -11831,
    36622 => -11834,
    36623 => -11837,
    36624 => -11840,
    36625 => -11842,
    36626 => -11845,
    36627 => -11848,
    36628 => -11851,
    36629 => -11854,
    36630 => -11857,
    36631 => -11860,
    36632 => -11863,
    36633 => -11866,
    36634 => -11869,
    36635 => -11872,
    36636 => -11875,
    36637 => -11878,
    36638 => -11881,
    36639 => -11883,
    36640 => -11886,
    36641 => -11889,
    36642 => -11892,
    36643 => -11895,
    36644 => -11898,
    36645 => -11901,
    36646 => -11904,
    36647 => -11907,
    36648 => -11910,
    36649 => -11913,
    36650 => -11916,
    36651 => -11919,
    36652 => -11922,
    36653 => -11924,
    36654 => -11927,
    36655 => -11930,
    36656 => -11933,
    36657 => -11936,
    36658 => -11939,
    36659 => -11942,
    36660 => -11945,
    36661 => -11948,
    36662 => -11951,
    36663 => -11954,
    36664 => -11957,
    36665 => -11960,
    36666 => -11962,
    36667 => -11965,
    36668 => -11968,
    36669 => -11971,
    36670 => -11974,
    36671 => -11977,
    36672 => -11980,
    36673 => -11983,
    36674 => -11986,
    36675 => -11989,
    36676 => -11992,
    36677 => -11995,
    36678 => -11998,
    36679 => -12001,
    36680 => -12003,
    36681 => -12006,
    36682 => -12009,
    36683 => -12012,
    36684 => -12015,
    36685 => -12018,
    36686 => -12021,
    36687 => -12024,
    36688 => -12027,
    36689 => -12030,
    36690 => -12033,
    36691 => -12036,
    36692 => -12038,
    36693 => -12041,
    36694 => -12044,
    36695 => -12047,
    36696 => -12050,
    36697 => -12053,
    36698 => -12056,
    36699 => -12059,
    36700 => -12062,
    36701 => -12065,
    36702 => -12068,
    36703 => -12071,
    36704 => -12074,
    36705 => -12076,
    36706 => -12079,
    36707 => -12082,
    36708 => -12085,
    36709 => -12088,
    36710 => -12091,
    36711 => -12094,
    36712 => -12097,
    36713 => -12100,
    36714 => -12103,
    36715 => -12106,
    36716 => -12109,
    36717 => -12112,
    36718 => -12114,
    36719 => -12117,
    36720 => -12120,
    36721 => -12123,
    36722 => -12126,
    36723 => -12129,
    36724 => -12132,
    36725 => -12135,
    36726 => -12138,
    36727 => -12141,
    36728 => -12144,
    36729 => -12147,
    36730 => -12149,
    36731 => -12152,
    36732 => -12155,
    36733 => -12158,
    36734 => -12161,
    36735 => -12164,
    36736 => -12167,
    36737 => -12170,
    36738 => -12173,
    36739 => -12176,
    36740 => -12179,
    36741 => -12182,
    36742 => -12184,
    36743 => -12187,
    36744 => -12190,
    36745 => -12193,
    36746 => -12196,
    36747 => -12199,
    36748 => -12202,
    36749 => -12205,
    36750 => -12208,
    36751 => -12211,
    36752 => -12214,
    36753 => -12217,
    36754 => -12219,
    36755 => -12222,
    36756 => -12225,
    36757 => -12228,
    36758 => -12231,
    36759 => -12234,
    36760 => -12237,
    36761 => -12240,
    36762 => -12243,
    36763 => -12246,
    36764 => -12249,
    36765 => -12251,
    36766 => -12254,
    36767 => -12257,
    36768 => -12260,
    36769 => -12263,
    36770 => -12266,
    36771 => -12269,
    36772 => -12272,
    36773 => -12275,
    36774 => -12278,
    36775 => -12281,
    36776 => -12284,
    36777 => -12286,
    36778 => -12289,
    36779 => -12292,
    36780 => -12295,
    36781 => -12298,
    36782 => -12301,
    36783 => -12304,
    36784 => -12307,
    36785 => -12310,
    36786 => -12313,
    36787 => -12316,
    36788 => -12318,
    36789 => -12321,
    36790 => -12324,
    36791 => -12327,
    36792 => -12330,
    36793 => -12333,
    36794 => -12336,
    36795 => -12339,
    36796 => -12342,
    36797 => -12345,
    36798 => -12348,
    36799 => -12350,
    36800 => -12353,
    36801 => -12356,
    36802 => -12359,
    36803 => -12362,
    36804 => -12365,
    36805 => -12368,
    36806 => -12371,
    36807 => -12374,
    36808 => -12377,
    36809 => -12380,
    36810 => -12382,
    36811 => -12385,
    36812 => -12388,
    36813 => -12391,
    36814 => -12394,
    36815 => -12397,
    36816 => -12400,
    36817 => -12403,
    36818 => -12406,
    36819 => -12409,
    36820 => -12412,
    36821 => -12414,
    36822 => -12417,
    36823 => -12420,
    36824 => -12423,
    36825 => -12426,
    36826 => -12429,
    36827 => -12432,
    36828 => -12435,
    36829 => -12438,
    36830 => -12441,
    36831 => -12444,
    36832 => -12446,
    36833 => -12449,
    36834 => -12452,
    36835 => -12455,
    36836 => -12458,
    36837 => -12461,
    36838 => -12464,
    36839 => -12467,
    36840 => -12470,
    36841 => -12473,
    36842 => -12476,
    36843 => -12478,
    36844 => -12481,
    36845 => -12484,
    36846 => -12487,
    36847 => -12490,
    36848 => -12493,
    36849 => -12496,
    36850 => -12499,
    36851 => -12502,
    36852 => -12505,
    36853 => -12507,
    36854 => -12510,
    36855 => -12513,
    36856 => -12516,
    36857 => -12519,
    36858 => -12522,
    36859 => -12525,
    36860 => -12528,
    36861 => -12531,
    36862 => -12534,
    36863 => -12536,
    36864 => -12539,
    36865 => -12542,
    36866 => -12545,
    36867 => -12548,
    36868 => -12551,
    36869 => -12554,
    36870 => -12557,
    36871 => -12560,
    36872 => -12563,
    36873 => -12566,
    36874 => -12568,
    36875 => -12571,
    36876 => -12574,
    36877 => -12577,
    36878 => -12580,
    36879 => -12583,
    36880 => -12586,
    36881 => -12589,
    36882 => -12592,
    36883 => -12595,
    36884 => -12597,
    36885 => -12600,
    36886 => -12603,
    36887 => -12606,
    36888 => -12609,
    36889 => -12612,
    36890 => -12615,
    36891 => -12618,
    36892 => -12621,
    36893 => -12624,
    36894 => -12626,
    36895 => -12629,
    36896 => -12632,
    36897 => -12635,
    36898 => -12638,
    36899 => -12641,
    36900 => -12644,
    36901 => -12647,
    36902 => -12650,
    36903 => -12652,
    36904 => -12655,
    36905 => -12658,
    36906 => -12661,
    36907 => -12664,
    36908 => -12667,
    36909 => -12670,
    36910 => -12673,
    36911 => -12676,
    36912 => -12679,
    36913 => -12681,
    36914 => -12684,
    36915 => -12687,
    36916 => -12690,
    36917 => -12693,
    36918 => -12696,
    36919 => -12699,
    36920 => -12702,
    36921 => -12705,
    36922 => -12708,
    36923 => -12710,
    36924 => -12713,
    36925 => -12716,
    36926 => -12719,
    36927 => -12722,
    36928 => -12725,
    36929 => -12728,
    36930 => -12731,
    36931 => -12734,
    36932 => -12736,
    36933 => -12739,
    36934 => -12742,
    36935 => -12745,
    36936 => -12748,
    36937 => -12751,
    36938 => -12754,
    36939 => -12757,
    36940 => -12760,
    36941 => -12763,
    36942 => -12765,
    36943 => -12768,
    36944 => -12771,
    36945 => -12774,
    36946 => -12777,
    36947 => -12780,
    36948 => -12783,
    36949 => -12786,
    36950 => -12789,
    36951 => -12791,
    36952 => -12794,
    36953 => -12797,
    36954 => -12800,
    36955 => -12803,
    36956 => -12806,
    36957 => -12809,
    36958 => -12812,
    36959 => -12815,
    36960 => -12817,
    36961 => -12820,
    36962 => -12823,
    36963 => -12826,
    36964 => -12829,
    36965 => -12832,
    36966 => -12835,
    36967 => -12838,
    36968 => -12841,
    36969 => -12843,
    36970 => -12846,
    36971 => -12849,
    36972 => -12852,
    36973 => -12855,
    36974 => -12858,
    36975 => -12861,
    36976 => -12864,
    36977 => -12867,
    36978 => -12870,
    36979 => -12872,
    36980 => -12875,
    36981 => -12878,
    36982 => -12881,
    36983 => -12884,
    36984 => -12887,
    36985 => -12890,
    36986 => -12893,
    36987 => -12895,
    36988 => -12898,
    36989 => -12901,
    36990 => -12904,
    36991 => -12907,
    36992 => -12910,
    36993 => -12913,
    36994 => -12916,
    36995 => -12919,
    36996 => -12921,
    36997 => -12924,
    36998 => -12927,
    36999 => -12930,
    37000 => -12933,
    37001 => -12936,
    37002 => -12939,
    37003 => -12942,
    37004 => -12945,
    37005 => -12947,
    37006 => -12950,
    37007 => -12953,
    37008 => -12956,
    37009 => -12959,
    37010 => -12962,
    37011 => -12965,
    37012 => -12968,
    37013 => -12971,
    37014 => -12973,
    37015 => -12976,
    37016 => -12979,
    37017 => -12982,
    37018 => -12985,
    37019 => -12988,
    37020 => -12991,
    37021 => -12994,
    37022 => -12997,
    37023 => -12999,
    37024 => -13002,
    37025 => -13005,
    37026 => -13008,
    37027 => -13011,
    37028 => -13014,
    37029 => -13017,
    37030 => -13020,
    37031 => -13022,
    37032 => -13025,
    37033 => -13028,
    37034 => -13031,
    37035 => -13034,
    37036 => -13037,
    37037 => -13040,
    37038 => -13043,
    37039 => -13046,
    37040 => -13048,
    37041 => -13051,
    37042 => -13054,
    37043 => -13057,
    37044 => -13060,
    37045 => -13063,
    37046 => -13066,
    37047 => -13069,
    37048 => -13071,
    37049 => -13074,
    37050 => -13077,
    37051 => -13080,
    37052 => -13083,
    37053 => -13086,
    37054 => -13089,
    37055 => -13092,
    37056 => -13094,
    37057 => -13097,
    37058 => -13100,
    37059 => -13103,
    37060 => -13106,
    37061 => -13109,
    37062 => -13112,
    37063 => -13115,
    37064 => -13118,
    37065 => -13120,
    37066 => -13123,
    37067 => -13126,
    37068 => -13129,
    37069 => -13132,
    37070 => -13135,
    37071 => -13138,
    37072 => -13141,
    37073 => -13143,
    37074 => -13146,
    37075 => -13149,
    37076 => -13152,
    37077 => -13155,
    37078 => -13158,
    37079 => -13161,
    37080 => -13164,
    37081 => -13166,
    37082 => -13169,
    37083 => -13172,
    37084 => -13175,
    37085 => -13178,
    37086 => -13181,
    37087 => -13184,
    37088 => -13187,
    37089 => -13189,
    37090 => -13192,
    37091 => -13195,
    37092 => -13198,
    37093 => -13201,
    37094 => -13204,
    37095 => -13207,
    37096 => -13210,
    37097 => -13212,
    37098 => -13215,
    37099 => -13218,
    37100 => -13221,
    37101 => -13224,
    37102 => -13227,
    37103 => -13230,
    37104 => -13233,
    37105 => -13235,
    37106 => -13238,
    37107 => -13241,
    37108 => -13244,
    37109 => -13247,
    37110 => -13250,
    37111 => -13253,
    37112 => -13256,
    37113 => -13258,
    37114 => -13261,
    37115 => -13264,
    37116 => -13267,
    37117 => -13270,
    37118 => -13273,
    37119 => -13276,
    37120 => -13279,
    37121 => -13281,
    37122 => -13284,
    37123 => -13287,
    37124 => -13290,
    37125 => -13293,
    37126 => -13296,
    37127 => -13299,
    37128 => -13302,
    37129 => -13304,
    37130 => -13307,
    37131 => -13310,
    37132 => -13313,
    37133 => -13316,
    37134 => -13319,
    37135 => -13322,
    37136 => -13324,
    37137 => -13327,
    37138 => -13330,
    37139 => -13333,
    37140 => -13336,
    37141 => -13339,
    37142 => -13342,
    37143 => -13345,
    37144 => -13347,
    37145 => -13350,
    37146 => -13353,
    37147 => -13356,
    37148 => -13359,
    37149 => -13362,
    37150 => -13365,
    37151 => -13368,
    37152 => -13370,
    37153 => -13373,
    37154 => -13376,
    37155 => -13379,
    37156 => -13382,
    37157 => -13385,
    37158 => -13388,
    37159 => -13390,
    37160 => -13393,
    37161 => -13396,
    37162 => -13399,
    37163 => -13402,
    37164 => -13405,
    37165 => -13408,
    37166 => -13411,
    37167 => -13413,
    37168 => -13416,
    37169 => -13419,
    37170 => -13422,
    37171 => -13425,
    37172 => -13428,
    37173 => -13431,
    37174 => -13433,
    37175 => -13436,
    37176 => -13439,
    37177 => -13442,
    37178 => -13445,
    37179 => -13448,
    37180 => -13451,
    37181 => -13454,
    37182 => -13456,
    37183 => -13459,
    37184 => -13462,
    37185 => -13465,
    37186 => -13468,
    37187 => -13471,
    37188 => -13474,
    37189 => -13476,
    37190 => -13479,
    37191 => -13482,
    37192 => -13485,
    37193 => -13488,
    37194 => -13491,
    37195 => -13494,
    37196 => -13496,
    37197 => -13499,
    37198 => -13502,
    37199 => -13505,
    37200 => -13508,
    37201 => -13511,
    37202 => -13514,
    37203 => -13516,
    37204 => -13519,
    37205 => -13522,
    37206 => -13525,
    37207 => -13528,
    37208 => -13531,
    37209 => -13534,
    37210 => -13537,
    37211 => -13539,
    37212 => -13542,
    37213 => -13545,
    37214 => -13548,
    37215 => -13551,
    37216 => -13554,
    37217 => -13557,
    37218 => -13559,
    37219 => -13562,
    37220 => -13565,
    37221 => -13568,
    37222 => -13571,
    37223 => -13574,
    37224 => -13577,
    37225 => -13579,
    37226 => -13582,
    37227 => -13585,
    37228 => -13588,
    37229 => -13591,
    37230 => -13594,
    37231 => -13597,
    37232 => -13599,
    37233 => -13602,
    37234 => -13605,
    37235 => -13608,
    37236 => -13611,
    37237 => -13614,
    37238 => -13617,
    37239 => -13619,
    37240 => -13622,
    37241 => -13625,
    37242 => -13628,
    37243 => -13631,
    37244 => -13634,
    37245 => -13637,
    37246 => -13639,
    37247 => -13642,
    37248 => -13645,
    37249 => -13648,
    37250 => -13651,
    37251 => -13654,
    37252 => -13657,
    37253 => -13659,
    37254 => -13662,
    37255 => -13665,
    37256 => -13668,
    37257 => -13671,
    37258 => -13674,
    37259 => -13677,
    37260 => -13679,
    37261 => -13682,
    37262 => -13685,
    37263 => -13688,
    37264 => -13691,
    37265 => -13694,
    37266 => -13697,
    37267 => -13699,
    37268 => -13702,
    37269 => -13705,
    37270 => -13708,
    37271 => -13711,
    37272 => -13714,
    37273 => -13717,
    37274 => -13719,
    37275 => -13722,
    37276 => -13725,
    37277 => -13728,
    37278 => -13731,
    37279 => -13734,
    37280 => -13736,
    37281 => -13739,
    37282 => -13742,
    37283 => -13745,
    37284 => -13748,
    37285 => -13751,
    37286 => -13754,
    37287 => -13756,
    37288 => -13759,
    37289 => -13762,
    37290 => -13765,
    37291 => -13768,
    37292 => -13771,
    37293 => -13774,
    37294 => -13776,
    37295 => -13779,
    37296 => -13782,
    37297 => -13785,
    37298 => -13788,
    37299 => -13791,
    37300 => -13793,
    37301 => -13796,
    37302 => -13799,
    37303 => -13802,
    37304 => -13805,
    37305 => -13808,
    37306 => -13811,
    37307 => -13813,
    37308 => -13816,
    37309 => -13819,
    37310 => -13822,
    37311 => -13825,
    37312 => -13828,
    37313 => -13831,
    37314 => -13833,
    37315 => -13836,
    37316 => -13839,
    37317 => -13842,
    37318 => -13845,
    37319 => -13848,
    37320 => -13850,
    37321 => -13853,
    37322 => -13856,
    37323 => -13859,
    37324 => -13862,
    37325 => -13865,
    37326 => -13868,
    37327 => -13870,
    37328 => -13873,
    37329 => -13876,
    37330 => -13879,
    37331 => -13882,
    37332 => -13885,
    37333 => -13887,
    37334 => -13890,
    37335 => -13893,
    37336 => -13896,
    37337 => -13899,
    37338 => -13902,
    37339 => -13905,
    37340 => -13907,
    37341 => -13910,
    37342 => -13913,
    37343 => -13916,
    37344 => -13919,
    37345 => -13922,
    37346 => -13924,
    37347 => -13927,
    37348 => -13930,
    37349 => -13933,
    37350 => -13936,
    37351 => -13939,
    37352 => -13942,
    37353 => -13944,
    37354 => -13947,
    37355 => -13950,
    37356 => -13953,
    37357 => -13956,
    37358 => -13959,
    37359 => -13961,
    37360 => -13964,
    37361 => -13967,
    37362 => -13970,
    37363 => -13973,
    37364 => -13976,
    37365 => -13978,
    37366 => -13981,
    37367 => -13984,
    37368 => -13987,
    37369 => -13990,
    37370 => -13993,
    37371 => -13995,
    37372 => -13998,
    37373 => -14001,
    37374 => -14004,
    37375 => -14007,
    37376 => -14010,
    37377 => -14013,
    37378 => -14015,
    37379 => -14018,
    37380 => -14021,
    37381 => -14024,
    37382 => -14027,
    37383 => -14030,
    37384 => -14032,
    37385 => -14035,
    37386 => -14038,
    37387 => -14041,
    37388 => -14044,
    37389 => -14047,
    37390 => -14049,
    37391 => -14052,
    37392 => -14055,
    37393 => -14058,
    37394 => -14061,
    37395 => -14064,
    37396 => -14066,
    37397 => -14069,
    37398 => -14072,
    37399 => -14075,
    37400 => -14078,
    37401 => -14081,
    37402 => -14083,
    37403 => -14086,
    37404 => -14089,
    37405 => -14092,
    37406 => -14095,
    37407 => -14098,
    37408 => -14101,
    37409 => -14103,
    37410 => -14106,
    37411 => -14109,
    37412 => -14112,
    37413 => -14115,
    37414 => -14118,
    37415 => -14120,
    37416 => -14123,
    37417 => -14126,
    37418 => -14129,
    37419 => -14132,
    37420 => -14135,
    37421 => -14137,
    37422 => -14140,
    37423 => -14143,
    37424 => -14146,
    37425 => -14149,
    37426 => -14152,
    37427 => -14154,
    37428 => -14157,
    37429 => -14160,
    37430 => -14163,
    37431 => -14166,
    37432 => -14169,
    37433 => -14171,
    37434 => -14174,
    37435 => -14177,
    37436 => -14180,
    37437 => -14183,
    37438 => -14186,
    37439 => -14188,
    37440 => -14191,
    37441 => -14194,
    37442 => -14197,
    37443 => -14200,
    37444 => -14203,
    37445 => -14205,
    37446 => -14208,
    37447 => -14211,
    37448 => -14214,
    37449 => -14217,
    37450 => -14219,
    37451 => -14222,
    37452 => -14225,
    37453 => -14228,
    37454 => -14231,
    37455 => -14234,
    37456 => -14236,
    37457 => -14239,
    37458 => -14242,
    37459 => -14245,
    37460 => -14248,
    37461 => -14251,
    37462 => -14253,
    37463 => -14256,
    37464 => -14259,
    37465 => -14262,
    37466 => -14265,
    37467 => -14268,
    37468 => -14270,
    37469 => -14273,
    37470 => -14276,
    37471 => -14279,
    37472 => -14282,
    37473 => -14285,
    37474 => -14287,
    37475 => -14290,
    37476 => -14293,
    37477 => -14296,
    37478 => -14299,
    37479 => -14302,
    37480 => -14304,
    37481 => -14307,
    37482 => -14310,
    37483 => -14313,
    37484 => -14316,
    37485 => -14318,
    37486 => -14321,
    37487 => -14324,
    37488 => -14327,
    37489 => -14330,
    37490 => -14333,
    37491 => -14335,
    37492 => -14338,
    37493 => -14341,
    37494 => -14344,
    37495 => -14347,
    37496 => -14350,
    37497 => -14352,
    37498 => -14355,
    37499 => -14358,
    37500 => -14361,
    37501 => -14364,
    37502 => -14366,
    37503 => -14369,
    37504 => -14372,
    37505 => -14375,
    37506 => -14378,
    37507 => -14381,
    37508 => -14383,
    37509 => -14386,
    37510 => -14389,
    37511 => -14392,
    37512 => -14395,
    37513 => -14398,
    37514 => -14400,
    37515 => -14403,
    37516 => -14406,
    37517 => -14409,
    37518 => -14412,
    37519 => -14414,
    37520 => -14417,
    37521 => -14420,
    37522 => -14423,
    37523 => -14426,
    37524 => -14429,
    37525 => -14431,
    37526 => -14434,
    37527 => -14437,
    37528 => -14440,
    37529 => -14443,
    37530 => -14445,
    37531 => -14448,
    37532 => -14451,
    37533 => -14454,
    37534 => -14457,
    37535 => -14460,
    37536 => -14462,
    37537 => -14465,
    37538 => -14468,
    37539 => -14471,
    37540 => -14474,
    37541 => -14477,
    37542 => -14479,
    37543 => -14482,
    37544 => -14485,
    37545 => -14488,
    37546 => -14491,
    37547 => -14493,
    37548 => -14496,
    37549 => -14499,
    37550 => -14502,
    37551 => -14505,
    37552 => -14507,
    37553 => -14510,
    37554 => -14513,
    37555 => -14516,
    37556 => -14519,
    37557 => -14522,
    37558 => -14524,
    37559 => -14527,
    37560 => -14530,
    37561 => -14533,
    37562 => -14536,
    37563 => -14538,
    37564 => -14541,
    37565 => -14544,
    37566 => -14547,
    37567 => -14550,
    37568 => -14553,
    37569 => -14555,
    37570 => -14558,
    37571 => -14561,
    37572 => -14564,
    37573 => -14567,
    37574 => -14569,
    37575 => -14572,
    37576 => -14575,
    37577 => -14578,
    37578 => -14581,
    37579 => -14584,
    37580 => -14586,
    37581 => -14589,
    37582 => -14592,
    37583 => -14595,
    37584 => -14598,
    37585 => -14600,
    37586 => -14603,
    37587 => -14606,
    37588 => -14609,
    37589 => -14612,
    37590 => -14614,
    37591 => -14617,
    37592 => -14620,
    37593 => -14623,
    37594 => -14626,
    37595 => -14628,
    37596 => -14631,
    37597 => -14634,
    37598 => -14637,
    37599 => -14640,
    37600 => -14643,
    37601 => -14645,
    37602 => -14648,
    37603 => -14651,
    37604 => -14654,
    37605 => -14657,
    37606 => -14659,
    37607 => -14662,
    37608 => -14665,
    37609 => -14668,
    37610 => -14671,
    37611 => -14673,
    37612 => -14676,
    37613 => -14679,
    37614 => -14682,
    37615 => -14685,
    37616 => -14688,
    37617 => -14690,
    37618 => -14693,
    37619 => -14696,
    37620 => -14699,
    37621 => -14702,
    37622 => -14704,
    37623 => -14707,
    37624 => -14710,
    37625 => -14713,
    37626 => -14716,
    37627 => -14718,
    37628 => -14721,
    37629 => -14724,
    37630 => -14727,
    37631 => -14730,
    37632 => -14732,
    37633 => -14735,
    37634 => -14738,
    37635 => -14741,
    37636 => -14744,
    37637 => -14746,
    37638 => -14749,
    37639 => -14752,
    37640 => -14755,
    37641 => -14758,
    37642 => -14760,
    37643 => -14763,
    37644 => -14766,
    37645 => -14769,
    37646 => -14772,
    37647 => -14774,
    37648 => -14777,
    37649 => -14780,
    37650 => -14783,
    37651 => -14786,
    37652 => -14789,
    37653 => -14791,
    37654 => -14794,
    37655 => -14797,
    37656 => -14800,
    37657 => -14803,
    37658 => -14805,
    37659 => -14808,
    37660 => -14811,
    37661 => -14814,
    37662 => -14817,
    37663 => -14819,
    37664 => -14822,
    37665 => -14825,
    37666 => -14828,
    37667 => -14831,
    37668 => -14833,
    37669 => -14836,
    37670 => -14839,
    37671 => -14842,
    37672 => -14845,
    37673 => -14847,
    37674 => -14850,
    37675 => -14853,
    37676 => -14856,
    37677 => -14859,
    37678 => -14861,
    37679 => -14864,
    37680 => -14867,
    37681 => -14870,
    37682 => -14873,
    37683 => -14875,
    37684 => -14878,
    37685 => -14881,
    37686 => -14884,
    37687 => -14887,
    37688 => -14889,
    37689 => -14892,
    37690 => -14895,
    37691 => -14898,
    37692 => -14901,
    37693 => -14903,
    37694 => -14906,
    37695 => -14909,
    37696 => -14912,
    37697 => -14915,
    37698 => -14917,
    37699 => -14920,
    37700 => -14923,
    37701 => -14926,
    37702 => -14929,
    37703 => -14931,
    37704 => -14934,
    37705 => -14937,
    37706 => -14940,
    37707 => -14942,
    37708 => -14945,
    37709 => -14948,
    37710 => -14951,
    37711 => -14954,
    37712 => -14956,
    37713 => -14959,
    37714 => -14962,
    37715 => -14965,
    37716 => -14968,
    37717 => -14970,
    37718 => -14973,
    37719 => -14976,
    37720 => -14979,
    37721 => -14982,
    37722 => -14984,
    37723 => -14987,
    37724 => -14990,
    37725 => -14993,
    37726 => -14996,
    37727 => -14998,
    37728 => -15001,
    37729 => -15004,
    37730 => -15007,
    37731 => -15010,
    37732 => -15012,
    37733 => -15015,
    37734 => -15018,
    37735 => -15021,
    37736 => -15024,
    37737 => -15026,
    37738 => -15029,
    37739 => -15032,
    37740 => -15035,
    37741 => -15037,
    37742 => -15040,
    37743 => -15043,
    37744 => -15046,
    37745 => -15049,
    37746 => -15051,
    37747 => -15054,
    37748 => -15057,
    37749 => -15060,
    37750 => -15063,
    37751 => -15065,
    37752 => -15068,
    37753 => -15071,
    37754 => -15074,
    37755 => -15077,
    37756 => -15079,
    37757 => -15082,
    37758 => -15085,
    37759 => -15088,
    37760 => -15090,
    37761 => -15093,
    37762 => -15096,
    37763 => -15099,
    37764 => -15102,
    37765 => -15104,
    37766 => -15107,
    37767 => -15110,
    37768 => -15113,
    37769 => -15116,
    37770 => -15118,
    37771 => -15121,
    37772 => -15124,
    37773 => -15127,
    37774 => -15129,
    37775 => -15132,
    37776 => -15135,
    37777 => -15138,
    37778 => -15141,
    37779 => -15143,
    37780 => -15146,
    37781 => -15149,
    37782 => -15152,
    37783 => -15155,
    37784 => -15157,
    37785 => -15160,
    37786 => -15163,
    37787 => -15166,
    37788 => -15168,
    37789 => -15171,
    37790 => -15174,
    37791 => -15177,
    37792 => -15180,
    37793 => -15182,
    37794 => -15185,
    37795 => -15188,
    37796 => -15191,
    37797 => -15194,
    37798 => -15196,
    37799 => -15199,
    37800 => -15202,
    37801 => -15205,
    37802 => -15207,
    37803 => -15210,
    37804 => -15213,
    37805 => -15216,
    37806 => -15219,
    37807 => -15221,
    37808 => -15224,
    37809 => -15227,
    37810 => -15230,
    37811 => -15233,
    37812 => -15235,
    37813 => -15238,
    37814 => -15241,
    37815 => -15244,
    37816 => -15246,
    37817 => -15249,
    37818 => -15252,
    37819 => -15255,
    37820 => -15258,
    37821 => -15260,
    37822 => -15263,
    37823 => -15266,
    37824 => -15269,
    37825 => -15271,
    37826 => -15274,
    37827 => -15277,
    37828 => -15280,
    37829 => -15283,
    37830 => -15285,
    37831 => -15288,
    37832 => -15291,
    37833 => -15294,
    37834 => -15296,
    37835 => -15299,
    37836 => -15302,
    37837 => -15305,
    37838 => -15308,
    37839 => -15310,
    37840 => -15313,
    37841 => -15316,
    37842 => -15319,
    37843 => -15321,
    37844 => -15324,
    37845 => -15327,
    37846 => -15330,
    37847 => -15333,
    37848 => -15335,
    37849 => -15338,
    37850 => -15341,
    37851 => -15344,
    37852 => -15346,
    37853 => -15349,
    37854 => -15352,
    37855 => -15355,
    37856 => -15358,
    37857 => -15360,
    37858 => -15363,
    37859 => -15366,
    37860 => -15369,
    37861 => -15371,
    37862 => -15374,
    37863 => -15377,
    37864 => -15380,
    37865 => -15382,
    37866 => -15385,
    37867 => -15388,
    37868 => -15391,
    37869 => -15394,
    37870 => -15396,
    37871 => -15399,
    37872 => -15402,
    37873 => -15405,
    37874 => -15407,
    37875 => -15410,
    37876 => -15413,
    37877 => -15416,
    37878 => -15419,
    37879 => -15421,
    37880 => -15424,
    37881 => -15427,
    37882 => -15430,
    37883 => -15432,
    37884 => -15435,
    37885 => -15438,
    37886 => -15441,
    37887 => -15443,
    37888 => -15446,
    37889 => -15449,
    37890 => -15452,
    37891 => -15455,
    37892 => -15457,
    37893 => -15460,
    37894 => -15463,
    37895 => -15466,
    37896 => -15468,
    37897 => -15471,
    37898 => -15474,
    37899 => -15477,
    37900 => -15479,
    37901 => -15482,
    37902 => -15485,
    37903 => -15488,
    37904 => -15491,
    37905 => -15493,
    37906 => -15496,
    37907 => -15499,
    37908 => -15502,
    37909 => -15504,
    37910 => -15507,
    37911 => -15510,
    37912 => -15513,
    37913 => -15515,
    37914 => -15518,
    37915 => -15521,
    37916 => -15524,
    37917 => -15527,
    37918 => -15529,
    37919 => -15532,
    37920 => -15535,
    37921 => -15538,
    37922 => -15540,
    37923 => -15543,
    37924 => -15546,
    37925 => -15549,
    37926 => -15551,
    37927 => -15554,
    37928 => -15557,
    37929 => -15560,
    37930 => -15562,
    37931 => -15565,
    37932 => -15568,
    37933 => -15571,
    37934 => -15574,
    37935 => -15576,
    37936 => -15579,
    37937 => -15582,
    37938 => -15585,
    37939 => -15587,
    37940 => -15590,
    37941 => -15593,
    37942 => -15596,
    37943 => -15598,
    37944 => -15601,
    37945 => -15604,
    37946 => -15607,
    37947 => -15609,
    37948 => -15612,
    37949 => -15615,
    37950 => -15618,
    37951 => -15621,
    37952 => -15623,
    37953 => -15626,
    37954 => -15629,
    37955 => -15632,
    37956 => -15634,
    37957 => -15637,
    37958 => -15640,
    37959 => -15643,
    37960 => -15645,
    37961 => -15648,
    37962 => -15651,
    37963 => -15654,
    37964 => -15656,
    37965 => -15659,
    37966 => -15662,
    37967 => -15665,
    37968 => -15667,
    37969 => -15670,
    37970 => -15673,
    37971 => -15676,
    37972 => -15678,
    37973 => -15681,
    37974 => -15684,
    37975 => -15687,
    37976 => -15690,
    37977 => -15692,
    37978 => -15695,
    37979 => -15698,
    37980 => -15701,
    37981 => -15703,
    37982 => -15706,
    37983 => -15709,
    37984 => -15712,
    37985 => -15714,
    37986 => -15717,
    37987 => -15720,
    37988 => -15723,
    37989 => -15725,
    37990 => -15728,
    37991 => -15731,
    37992 => -15734,
    37993 => -15736,
    37994 => -15739,
    37995 => -15742,
    37996 => -15745,
    37997 => -15747,
    37998 => -15750,
    37999 => -15753,
    38000 => -15756,
    38001 => -15758,
    38002 => -15761,
    38003 => -15764,
    38004 => -15767,
    38005 => -15769,
    38006 => -15772,
    38007 => -15775,
    38008 => -15778,
    38009 => -15780,
    38010 => -15783,
    38011 => -15786,
    38012 => -15789,
    38013 => -15791,
    38014 => -15794,
    38015 => -15797,
    38016 => -15800,
    38017 => -15802,
    38018 => -15805,
    38019 => -15808,
    38020 => -15811,
    38021 => -15813,
    38022 => -15816,
    38023 => -15819,
    38024 => -15822,
    38025 => -15824,
    38026 => -15827,
    38027 => -15830,
    38028 => -15833,
    38029 => -15835,
    38030 => -15838,
    38031 => -15841,
    38032 => -15844,
    38033 => -15846,
    38034 => -15849,
    38035 => -15852,
    38036 => -15855,
    38037 => -15857,
    38038 => -15860,
    38039 => -15863,
    38040 => -15866,
    38041 => -15868,
    38042 => -15871,
    38043 => -15874,
    38044 => -15877,
    38045 => -15879,
    38046 => -15882,
    38047 => -15885,
    38048 => -15888,
    38049 => -15890,
    38050 => -15893,
    38051 => -15896,
    38052 => -15899,
    38053 => -15901,
    38054 => -15904,
    38055 => -15907,
    38056 => -15910,
    38057 => -15912,
    38058 => -15915,
    38059 => -15918,
    38060 => -15921,
    38061 => -15923,
    38062 => -15926,
    38063 => -15929,
    38064 => -15932,
    38065 => -15934,
    38066 => -15937,
    38067 => -15940,
    38068 => -15943,
    38069 => -15945,
    38070 => -15948,
    38071 => -15951,
    38072 => -15954,
    38073 => -15956,
    38074 => -15959,
    38075 => -15962,
    38076 => -15965,
    38077 => -15967,
    38078 => -15970,
    38079 => -15973,
    38080 => -15976,
    38081 => -15978,
    38082 => -15981,
    38083 => -15984,
    38084 => -15987,
    38085 => -15989,
    38086 => -15992,
    38087 => -15995,
    38088 => -15997,
    38089 => -16000,
    38090 => -16003,
    38091 => -16006,
    38092 => -16008,
    38093 => -16011,
    38094 => -16014,
    38095 => -16017,
    38096 => -16019,
    38097 => -16022,
    38098 => -16025,
    38099 => -16028,
    38100 => -16030,
    38101 => -16033,
    38102 => -16036,
    38103 => -16039,
    38104 => -16041,
    38105 => -16044,
    38106 => -16047,
    38107 => -16050,
    38108 => -16052,
    38109 => -16055,
    38110 => -16058,
    38111 => -16061,
    38112 => -16063,
    38113 => -16066,
    38114 => -16069,
    38115 => -16071,
    38116 => -16074,
    38117 => -16077,
    38118 => -16080,
    38119 => -16082,
    38120 => -16085,
    38121 => -16088,
    38122 => -16091,
    38123 => -16093,
    38124 => -16096,
    38125 => -16099,
    38126 => -16102,
    38127 => -16104,
    38128 => -16107,
    38129 => -16110,
    38130 => -16113,
    38131 => -16115,
    38132 => -16118,
    38133 => -16121,
    38134 => -16123,
    38135 => -16126,
    38136 => -16129,
    38137 => -16132,
    38138 => -16134,
    38139 => -16137,
    38140 => -16140,
    38141 => -16143,
    38142 => -16145,
    38143 => -16148,
    38144 => -16151,
    38145 => -16154,
    38146 => -16156,
    38147 => -16159,
    38148 => -16162,
    38149 => -16164,
    38150 => -16167,
    38151 => -16170,
    38152 => -16173,
    38153 => -16175,
    38154 => -16178,
    38155 => -16181,
    38156 => -16184,
    38157 => -16186,
    38158 => -16189,
    38159 => -16192,
    38160 => -16195,
    38161 => -16197,
    38162 => -16200,
    38163 => -16203,
    38164 => -16205,
    38165 => -16208,
    38166 => -16211,
    38167 => -16214,
    38168 => -16216,
    38169 => -16219,
    38170 => -16222,
    38171 => -16225,
    38172 => -16227,
    38173 => -16230,
    38174 => -16233,
    38175 => -16235,
    38176 => -16238,
    38177 => -16241,
    38178 => -16244,
    38179 => -16246,
    38180 => -16249,
    38181 => -16252,
    38182 => -16255,
    38183 => -16257,
    38184 => -16260,
    38185 => -16263,
    38186 => -16265,
    38187 => -16268,
    38188 => -16271,
    38189 => -16274,
    38190 => -16276,
    38191 => -16279,
    38192 => -16282,
    38193 => -16285,
    38194 => -16287,
    38195 => -16290,
    38196 => -16293,
    38197 => -16295,
    38198 => -16298,
    38199 => -16301,
    38200 => -16304,
    38201 => -16306,
    38202 => -16309,
    38203 => -16312,
    38204 => -16315,
    38205 => -16317,
    38206 => -16320,
    38207 => -16323,
    38208 => -16325,
    38209 => -16328,
    38210 => -16331,
    38211 => -16334,
    38212 => -16336,
    38213 => -16339,
    38214 => -16342,
    38215 => -16344,
    38216 => -16347,
    38217 => -16350,
    38218 => -16353,
    38219 => -16355,
    38220 => -16358,
    38221 => -16361,
    38222 => -16364,
    38223 => -16366,
    38224 => -16369,
    38225 => -16372,
    38226 => -16374,
    38227 => -16377,
    38228 => -16380,
    38229 => -16383,
    38230 => -16385,
    38231 => -16388,
    38232 => -16391,
    38233 => -16393,
    38234 => -16396,
    38235 => -16399,
    38236 => -16402,
    38237 => -16404,
    38238 => -16407,
    38239 => -16410,
    38240 => -16413,
    38241 => -16415,
    38242 => -16418,
    38243 => -16421,
    38244 => -16423,
    38245 => -16426,
    38246 => -16429,
    38247 => -16432,
    38248 => -16434,
    38249 => -16437,
    38250 => -16440,
    38251 => -16442,
    38252 => -16445,
    38253 => -16448,
    38254 => -16451,
    38255 => -16453,
    38256 => -16456,
    38257 => -16459,
    38258 => -16461,
    38259 => -16464,
    38260 => -16467,
    38261 => -16470,
    38262 => -16472,
    38263 => -16475,
    38264 => -16478,
    38265 => -16480,
    38266 => -16483,
    38267 => -16486,
    38268 => -16489,
    38269 => -16491,
    38270 => -16494,
    38271 => -16497,
    38272 => -16499,
    38273 => -16502,
    38274 => -16505,
    38275 => -16508,
    38276 => -16510,
    38277 => -16513,
    38278 => -16516,
    38279 => -16518,
    38280 => -16521,
    38281 => -16524,
    38282 => -16527,
    38283 => -16529,
    38284 => -16532,
    38285 => -16535,
    38286 => -16537,
    38287 => -16540,
    38288 => -16543,
    38289 => -16546,
    38290 => -16548,
    38291 => -16551,
    38292 => -16554,
    38293 => -16556,
    38294 => -16559,
    38295 => -16562,
    38296 => -16565,
    38297 => -16567,
    38298 => -16570,
    38299 => -16573,
    38300 => -16575,
    38301 => -16578,
    38302 => -16581,
    38303 => -16584,
    38304 => -16586,
    38305 => -16589,
    38306 => -16592,
    38307 => -16594,
    38308 => -16597,
    38309 => -16600,
    38310 => -16602,
    38311 => -16605,
    38312 => -16608,
    38313 => -16611,
    38314 => -16613,
    38315 => -16616,
    38316 => -16619,
    38317 => -16621,
    38318 => -16624,
    38319 => -16627,
    38320 => -16630,
    38321 => -16632,
    38322 => -16635,
    38323 => -16638,
    38324 => -16640,
    38325 => -16643,
    38326 => -16646,
    38327 => -16648,
    38328 => -16651,
    38329 => -16654,
    38330 => -16657,
    38331 => -16659,
    38332 => -16662,
    38333 => -16665,
    38334 => -16667,
    38335 => -16670,
    38336 => -16673,
    38337 => -16676,
    38338 => -16678,
    38339 => -16681,
    38340 => -16684,
    38341 => -16686,
    38342 => -16689,
    38343 => -16692,
    38344 => -16694,
    38345 => -16697,
    38346 => -16700,
    38347 => -16703,
    38348 => -16705,
    38349 => -16708,
    38350 => -16711,
    38351 => -16713,
    38352 => -16716,
    38353 => -16719,
    38354 => -16721,
    38355 => -16724,
    38356 => -16727,
    38357 => -16730,
    38358 => -16732,
    38359 => -16735,
    38360 => -16738,
    38361 => -16740,
    38362 => -16743,
    38363 => -16746,
    38364 => -16749,
    38365 => -16751,
    38366 => -16754,
    38367 => -16757,
    38368 => -16759,
    38369 => -16762,
    38370 => -16765,
    38371 => -16767,
    38372 => -16770,
    38373 => -16773,
    38374 => -16775,
    38375 => -16778,
    38376 => -16781,
    38377 => -16784,
    38378 => -16786,
    38379 => -16789,
    38380 => -16792,
    38381 => -16794,
    38382 => -16797,
    38383 => -16800,
    38384 => -16802,
    38385 => -16805,
    38386 => -16808,
    38387 => -16811,
    38388 => -16813,
    38389 => -16816,
    38390 => -16819,
    38391 => -16821,
    38392 => -16824,
    38393 => -16827,
    38394 => -16829,
    38395 => -16832,
    38396 => -16835,
    38397 => -16838,
    38398 => -16840,
    38399 => -16843,
    38400 => -16846,
    38401 => -16848,
    38402 => -16851,
    38403 => -16854,
    38404 => -16856,
    38405 => -16859,
    38406 => -16862,
    38407 => -16864,
    38408 => -16867,
    38409 => -16870,
    38410 => -16873,
    38411 => -16875,
    38412 => -16878,
    38413 => -16881,
    38414 => -16883,
    38415 => -16886,
    38416 => -16889,
    38417 => -16891,
    38418 => -16894,
    38419 => -16897,
    38420 => -16899,
    38421 => -16902,
    38422 => -16905,
    38423 => -16908,
    38424 => -16910,
    38425 => -16913,
    38426 => -16916,
    38427 => -16918,
    38428 => -16921,
    38429 => -16924,
    38430 => -16926,
    38431 => -16929,
    38432 => -16932,
    38433 => -16934,
    38434 => -16937,
    38435 => -16940,
    38436 => -16943,
    38437 => -16945,
    38438 => -16948,
    38439 => -16951,
    38440 => -16953,
    38441 => -16956,
    38442 => -16959,
    38443 => -16961,
    38444 => -16964,
    38445 => -16967,
    38446 => -16969,
    38447 => -16972,
    38448 => -16975,
    38449 => -16977,
    38450 => -16980,
    38451 => -16983,
    38452 => -16986,
    38453 => -16988,
    38454 => -16991,
    38455 => -16994,
    38456 => -16996,
    38457 => -16999,
    38458 => -17002,
    38459 => -17004,
    38460 => -17007,
    38461 => -17010,
    38462 => -17012,
    38463 => -17015,
    38464 => -17018,
    38465 => -17020,
    38466 => -17023,
    38467 => -17026,
    38468 => -17028,
    38469 => -17031,
    38470 => -17034,
    38471 => -17037,
    38472 => -17039,
    38473 => -17042,
    38474 => -17045,
    38475 => -17047,
    38476 => -17050,
    38477 => -17053,
    38478 => -17055,
    38479 => -17058,
    38480 => -17061,
    38481 => -17063,
    38482 => -17066,
    38483 => -17069,
    38484 => -17071,
    38485 => -17074,
    38486 => -17077,
    38487 => -17079,
    38488 => -17082,
    38489 => -17085,
    38490 => -17087,
    38491 => -17090,
    38492 => -17093,
    38493 => -17096,
    38494 => -17098,
    38495 => -17101,
    38496 => -17104,
    38497 => -17106,
    38498 => -17109,
    38499 => -17112,
    38500 => -17114,
    38501 => -17117,
    38502 => -17120,
    38503 => -17122,
    38504 => -17125,
    38505 => -17128,
    38506 => -17130,
    38507 => -17133,
    38508 => -17136,
    38509 => -17138,
    38510 => -17141,
    38511 => -17144,
    38512 => -17146,
    38513 => -17149,
    38514 => -17152,
    38515 => -17154,
    38516 => -17157,
    38517 => -17160,
    38518 => -17162,
    38519 => -17165,
    38520 => -17168,
    38521 => -17171,
    38522 => -17173,
    38523 => -17176,
    38524 => -17179,
    38525 => -17181,
    38526 => -17184,
    38527 => -17187,
    38528 => -17189,
    38529 => -17192,
    38530 => -17195,
    38531 => -17197,
    38532 => -17200,
    38533 => -17203,
    38534 => -17205,
    38535 => -17208,
    38536 => -17211,
    38537 => -17213,
    38538 => -17216,
    38539 => -17219,
    38540 => -17221,
    38541 => -17224,
    38542 => -17227,
    38543 => -17229,
    38544 => -17232,
    38545 => -17235,
    38546 => -17237,
    38547 => -17240,
    38548 => -17243,
    38549 => -17245,
    38550 => -17248,
    38551 => -17251,
    38552 => -17253,
    38553 => -17256,
    38554 => -17259,
    38555 => -17261,
    38556 => -17264,
    38557 => -17267,
    38558 => -17269,
    38559 => -17272,
    38560 => -17275,
    38561 => -17277,
    38562 => -17280,
    38563 => -17283,
    38564 => -17285,
    38565 => -17288,
    38566 => -17291,
    38567 => -17293,
    38568 => -17296,
    38569 => -17299,
    38570 => -17301,
    38571 => -17304,
    38572 => -17307,
    38573 => -17309,
    38574 => -17312,
    38575 => -17315,
    38576 => -17317,
    38577 => -17320,
    38578 => -17323,
    38579 => -17325,
    38580 => -17328,
    38581 => -17331,
    38582 => -17333,
    38583 => -17336,
    38584 => -17339,
    38585 => -17341,
    38586 => -17344,
    38587 => -17347,
    38588 => -17349,
    38589 => -17352,
    38590 => -17355,
    38591 => -17357,
    38592 => -17360,
    38593 => -17363,
    38594 => -17365,
    38595 => -17368,
    38596 => -17371,
    38597 => -17373,
    38598 => -17376,
    38599 => -17379,
    38600 => -17381,
    38601 => -17384,
    38602 => -17387,
    38603 => -17389,
    38604 => -17392,
    38605 => -17395,
    38606 => -17397,
    38607 => -17400,
    38608 => -17403,
    38609 => -17405,
    38610 => -17408,
    38611 => -17411,
    38612 => -17413,
    38613 => -17416,
    38614 => -17419,
    38615 => -17421,
    38616 => -17424,
    38617 => -17427,
    38618 => -17429,
    38619 => -17432,
    38620 => -17435,
    38621 => -17437,
    38622 => -17440,
    38623 => -17443,
    38624 => -17445,
    38625 => -17448,
    38626 => -17451,
    38627 => -17453,
    38628 => -17456,
    38629 => -17459,
    38630 => -17461,
    38631 => -17464,
    38632 => -17467,
    38633 => -17469,
    38634 => -17472,
    38635 => -17474,
    38636 => -17477,
    38637 => -17480,
    38638 => -17482,
    38639 => -17485,
    38640 => -17488,
    38641 => -17490,
    38642 => -17493,
    38643 => -17496,
    38644 => -17498,
    38645 => -17501,
    38646 => -17504,
    38647 => -17506,
    38648 => -17509,
    38649 => -17512,
    38650 => -17514,
    38651 => -17517,
    38652 => -17520,
    38653 => -17522,
    38654 => -17525,
    38655 => -17528,
    38656 => -17530,
    38657 => -17533,
    38658 => -17536,
    38659 => -17538,
    38660 => -17541,
    38661 => -17544,
    38662 => -17546,
    38663 => -17549,
    38664 => -17551,
    38665 => -17554,
    38666 => -17557,
    38667 => -17559,
    38668 => -17562,
    38669 => -17565,
    38670 => -17567,
    38671 => -17570,
    38672 => -17573,
    38673 => -17575,
    38674 => -17578,
    38675 => -17581,
    38676 => -17583,
    38677 => -17586,
    38678 => -17589,
    38679 => -17591,
    38680 => -17594,
    38681 => -17597,
    38682 => -17599,
    38683 => -17602,
    38684 => -17605,
    38685 => -17607,
    38686 => -17610,
    38687 => -17612,
    38688 => -17615,
    38689 => -17618,
    38690 => -17620,
    38691 => -17623,
    38692 => -17626,
    38693 => -17628,
    38694 => -17631,
    38695 => -17634,
    38696 => -17636,
    38697 => -17639,
    38698 => -17642,
    38699 => -17644,
    38700 => -17647,
    38701 => -17650,
    38702 => -17652,
    38703 => -17655,
    38704 => -17657,
    38705 => -17660,
    38706 => -17663,
    38707 => -17665,
    38708 => -17668,
    38709 => -17671,
    38710 => -17673,
    38711 => -17676,
    38712 => -17679,
    38713 => -17681,
    38714 => -17684,
    38715 => -17687,
    38716 => -17689,
    38717 => -17692,
    38718 => -17695,
    38719 => -17697,
    38720 => -17700,
    38721 => -17702,
    38722 => -17705,
    38723 => -17708,
    38724 => -17710,
    38725 => -17713,
    38726 => -17716,
    38727 => -17718,
    38728 => -17721,
    38729 => -17724,
    38730 => -17726,
    38731 => -17729,
    38732 => -17732,
    38733 => -17734,
    38734 => -17737,
    38735 => -17739,
    38736 => -17742,
    38737 => -17745,
    38738 => -17747,
    38739 => -17750,
    38740 => -17753,
    38741 => -17755,
    38742 => -17758,
    38743 => -17761,
    38744 => -17763,
    38745 => -17766,
    38746 => -17768,
    38747 => -17771,
    38748 => -17774,
    38749 => -17776,
    38750 => -17779,
    38751 => -17782,
    38752 => -17784,
    38753 => -17787,
    38754 => -17790,
    38755 => -17792,
    38756 => -17795,
    38757 => -17798,
    38758 => -17800,
    38759 => -17803,
    38760 => -17805,
    38761 => -17808,
    38762 => -17811,
    38763 => -17813,
    38764 => -17816,
    38765 => -17819,
    38766 => -17821,
    38767 => -17824,
    38768 => -17827,
    38769 => -17829,
    38770 => -17832,
    38771 => -17834,
    38772 => -17837,
    38773 => -17840,
    38774 => -17842,
    38775 => -17845,
    38776 => -17848,
    38777 => -17850,
    38778 => -17853,
    38779 => -17855,
    38780 => -17858,
    38781 => -17861,
    38782 => -17863,
    38783 => -17866,
    38784 => -17869,
    38785 => -17871,
    38786 => -17874,
    38787 => -17877,
    38788 => -17879,
    38789 => -17882,
    38790 => -17884,
    38791 => -17887,
    38792 => -17890,
    38793 => -17892,
    38794 => -17895,
    38795 => -17898,
    38796 => -17900,
    38797 => -17903,
    38798 => -17906,
    38799 => -17908,
    38800 => -17911,
    38801 => -17913,
    38802 => -17916,
    38803 => -17919,
    38804 => -17921,
    38805 => -17924,
    38806 => -17927,
    38807 => -17929,
    38808 => -17932,
    38809 => -17934,
    38810 => -17937,
    38811 => -17940,
    38812 => -17942,
    38813 => -17945,
    38814 => -17948,
    38815 => -17950,
    38816 => -17953,
    38817 => -17955,
    38818 => -17958,
    38819 => -17961,
    38820 => -17963,
    38821 => -17966,
    38822 => -17969,
    38823 => -17971,
    38824 => -17974,
    38825 => -17976,
    38826 => -17979,
    38827 => -17982,
    38828 => -17984,
    38829 => -17987,
    38830 => -17990,
    38831 => -17992,
    38832 => -17995,
    38833 => -17997,
    38834 => -18000,
    38835 => -18003,
    38836 => -18005,
    38837 => -18008,
    38838 => -18011,
    38839 => -18013,
    38840 => -18016,
    38841 => -18018,
    38842 => -18021,
    38843 => -18024,
    38844 => -18026,
    38845 => -18029,
    38846 => -18032,
    38847 => -18034,
    38848 => -18037,
    38849 => -18039,
    38850 => -18042,
    38851 => -18045,
    38852 => -18047,
    38853 => -18050,
    38854 => -18053,
    38855 => -18055,
    38856 => -18058,
    38857 => -18060,
    38858 => -18063,
    38859 => -18066,
    38860 => -18068,
    38861 => -18071,
    38862 => -18074,
    38863 => -18076,
    38864 => -18079,
    38865 => -18081,
    38866 => -18084,
    38867 => -18087,
    38868 => -18089,
    38869 => -18092,
    38870 => -18095,
    38871 => -18097,
    38872 => -18100,
    38873 => -18102,
    38874 => -18105,
    38875 => -18108,
    38876 => -18110,
    38877 => -18113,
    38878 => -18115,
    38879 => -18118,
    38880 => -18121,
    38881 => -18123,
    38882 => -18126,
    38883 => -18129,
    38884 => -18131,
    38885 => -18134,
    38886 => -18136,
    38887 => -18139,
    38888 => -18142,
    38889 => -18144,
    38890 => -18147,
    38891 => -18149,
    38892 => -18152,
    38893 => -18155,
    38894 => -18157,
    38895 => -18160,
    38896 => -18163,
    38897 => -18165,
    38898 => -18168,
    38899 => -18170,
    38900 => -18173,
    38901 => -18176,
    38902 => -18178,
    38903 => -18181,
    38904 => -18183,
    38905 => -18186,
    38906 => -18189,
    38907 => -18191,
    38908 => -18194,
    38909 => -18197,
    38910 => -18199,
    38911 => -18202,
    38912 => -18204,
    38913 => -18207,
    38914 => -18210,
    38915 => -18212,
    38916 => -18215,
    38917 => -18217,
    38918 => -18220,
    38919 => -18223,
    38920 => -18225,
    38921 => -18228,
    38922 => -18230,
    38923 => -18233,
    38924 => -18236,
    38925 => -18238,
    38926 => -18241,
    38927 => -18244,
    38928 => -18246,
    38929 => -18249,
    38930 => -18251,
    38931 => -18254,
    38932 => -18257,
    38933 => -18259,
    38934 => -18262,
    38935 => -18264,
    38936 => -18267,
    38937 => -18270,
    38938 => -18272,
    38939 => -18275,
    38940 => -18277,
    38941 => -18280,
    38942 => -18283,
    38943 => -18285,
    38944 => -18288,
    38945 => -18290,
    38946 => -18293,
    38947 => -18296,
    38948 => -18298,
    38949 => -18301,
    38950 => -18304,
    38951 => -18306,
    38952 => -18309,
    38953 => -18311,
    38954 => -18314,
    38955 => -18317,
    38956 => -18319,
    38957 => -18322,
    38958 => -18324,
    38959 => -18327,
    38960 => -18330,
    38961 => -18332,
    38962 => -18335,
    38963 => -18337,
    38964 => -18340,
    38965 => -18343,
    38966 => -18345,
    38967 => -18348,
    38968 => -18350,
    38969 => -18353,
    38970 => -18356,
    38971 => -18358,
    38972 => -18361,
    38973 => -18363,
    38974 => -18366,
    38975 => -18369,
    38976 => -18371,
    38977 => -18374,
    38978 => -18376,
    38979 => -18379,
    38980 => -18382,
    38981 => -18384,
    38982 => -18387,
    38983 => -18389,
    38984 => -18392,
    38985 => -18395,
    38986 => -18397,
    38987 => -18400,
    38988 => -18402,
    38989 => -18405,
    38990 => -18408,
    38991 => -18410,
    38992 => -18413,
    38993 => -18415,
    38994 => -18418,
    38995 => -18421,
    38996 => -18423,
    38997 => -18426,
    38998 => -18428,
    38999 => -18431,
    39000 => -18434,
    39001 => -18436,
    39002 => -18439,
    39003 => -18441,
    39004 => -18444,
    39005 => -18447,
    39006 => -18449,
    39007 => -18452,
    39008 => -18454,
    39009 => -18457,
    39010 => -18460,
    39011 => -18462,
    39012 => -18465,
    39013 => -18467,
    39014 => -18470,
    39015 => -18473,
    39016 => -18475,
    39017 => -18478,
    39018 => -18480,
    39019 => -18483,
    39020 => -18485,
    39021 => -18488,
    39022 => -18491,
    39023 => -18493,
    39024 => -18496,
    39025 => -18498,
    39026 => -18501,
    39027 => -18504,
    39028 => -18506,
    39029 => -18509,
    39030 => -18511,
    39031 => -18514,
    39032 => -18517,
    39033 => -18519,
    39034 => -18522,
    39035 => -18524,
    39036 => -18527,
    39037 => -18530,
    39038 => -18532,
    39039 => -18535,
    39040 => -18537,
    39041 => -18540,
    39042 => -18543,
    39043 => -18545,
    39044 => -18548,
    39045 => -18550,
    39046 => -18553,
    39047 => -18555,
    39048 => -18558,
    39049 => -18561,
    39050 => -18563,
    39051 => -18566,
    39052 => -18568,
    39053 => -18571,
    39054 => -18574,
    39055 => -18576,
    39056 => -18579,
    39057 => -18581,
    39058 => -18584,
    39059 => -18587,
    39060 => -18589,
    39061 => -18592,
    39062 => -18594,
    39063 => -18597,
    39064 => -18599,
    39065 => -18602,
    39066 => -18605,
    39067 => -18607,
    39068 => -18610,
    39069 => -18612,
    39070 => -18615,
    39071 => -18618,
    39072 => -18620,
    39073 => -18623,
    39074 => -18625,
    39075 => -18628,
    39076 => -18630,
    39077 => -18633,
    39078 => -18636,
    39079 => -18638,
    39080 => -18641,
    39081 => -18643,
    39082 => -18646,
    39083 => -18649,
    39084 => -18651,
    39085 => -18654,
    39086 => -18656,
    39087 => -18659,
    39088 => -18661,
    39089 => -18664,
    39090 => -18667,
    39091 => -18669,
    39092 => -18672,
    39093 => -18674,
    39094 => -18677,
    39095 => -18680,
    39096 => -18682,
    39097 => -18685,
    39098 => -18687,
    39099 => -18690,
    39100 => -18692,
    39101 => -18695,
    39102 => -18698,
    39103 => -18700,
    39104 => -18703,
    39105 => -18705,
    39106 => -18708,
    39107 => -18711,
    39108 => -18713,
    39109 => -18716,
    39110 => -18718,
    39111 => -18721,
    39112 => -18723,
    39113 => -18726,
    39114 => -18729,
    39115 => -18731,
    39116 => -18734,
    39117 => -18736,
    39118 => -18739,
    39119 => -18741,
    39120 => -18744,
    39121 => -18747,
    39122 => -18749,
    39123 => -18752,
    39124 => -18754,
    39125 => -18757,
    39126 => -18759,
    39127 => -18762,
    39128 => -18765,
    39129 => -18767,
    39130 => -18770,
    39131 => -18772,
    39132 => -18775,
    39133 => -18778,
    39134 => -18780,
    39135 => -18783,
    39136 => -18785,
    39137 => -18788,
    39138 => -18790,
    39139 => -18793,
    39140 => -18796,
    39141 => -18798,
    39142 => -18801,
    39143 => -18803,
    39144 => -18806,
    39145 => -18808,
    39146 => -18811,
    39147 => -18814,
    39148 => -18816,
    39149 => -18819,
    39150 => -18821,
    39151 => -18824,
    39152 => -18826,
    39153 => -18829,
    39154 => -18832,
    39155 => -18834,
    39156 => -18837,
    39157 => -18839,
    39158 => -18842,
    39159 => -18844,
    39160 => -18847,
    39161 => -18850,
    39162 => -18852,
    39163 => -18855,
    39164 => -18857,
    39165 => -18860,
    39166 => -18862,
    39167 => -18865,
    39168 => -18868,
    39169 => -18870,
    39170 => -18873,
    39171 => -18875,
    39172 => -18878,
    39173 => -18880,
    39174 => -18883,
    39175 => -18885,
    39176 => -18888,
    39177 => -18891,
    39178 => -18893,
    39179 => -18896,
    39180 => -18898,
    39181 => -18901,
    39182 => -18903,
    39183 => -18906,
    39184 => -18909,
    39185 => -18911,
    39186 => -18914,
    39187 => -18916,
    39188 => -18919,
    39189 => -18921,
    39190 => -18924,
    39191 => -18927,
    39192 => -18929,
    39193 => -18932,
    39194 => -18934,
    39195 => -18937,
    39196 => -18939,
    39197 => -18942,
    39198 => -18944,
    39199 => -18947,
    39200 => -18950,
    39201 => -18952,
    39202 => -18955,
    39203 => -18957,
    39204 => -18960,
    39205 => -18962,
    39206 => -18965,
    39207 => -18968,
    39208 => -18970,
    39209 => -18973,
    39210 => -18975,
    39211 => -18978,
    39212 => -18980,
    39213 => -18983,
    39214 => -18985,
    39215 => -18988,
    39216 => -18991,
    39217 => -18993,
    39218 => -18996,
    39219 => -18998,
    39220 => -19001,
    39221 => -19003,
    39222 => -19006,
    39223 => -19009,
    39224 => -19011,
    39225 => -19014,
    39226 => -19016,
    39227 => -19019,
    39228 => -19021,
    39229 => -19024,
    39230 => -19026,
    39231 => -19029,
    39232 => -19032,
    39233 => -19034,
    39234 => -19037,
    39235 => -19039,
    39236 => -19042,
    39237 => -19044,
    39238 => -19047,
    39239 => -19049,
    39240 => -19052,
    39241 => -19055,
    39242 => -19057,
    39243 => -19060,
    39244 => -19062,
    39245 => -19065,
    39246 => -19067,
    39247 => -19070,
    39248 => -19072,
    39249 => -19075,
    39250 => -19078,
    39251 => -19080,
    39252 => -19083,
    39253 => -19085,
    39254 => -19088,
    39255 => -19090,
    39256 => -19093,
    39257 => -19095,
    39258 => -19098,
    39259 => -19101,
    39260 => -19103,
    39261 => -19106,
    39262 => -19108,
    39263 => -19111,
    39264 => -19113,
    39265 => -19116,
    39266 => -19118,
    39267 => -19121,
    39268 => -19123,
    39269 => -19126,
    39270 => -19129,
    39271 => -19131,
    39272 => -19134,
    39273 => -19136,
    39274 => -19139,
    39275 => -19141,
    39276 => -19144,
    39277 => -19146,
    39278 => -19149,
    39279 => -19152,
    39280 => -19154,
    39281 => -19157,
    39282 => -19159,
    39283 => -19162,
    39284 => -19164,
    39285 => -19167,
    39286 => -19169,
    39287 => -19172,
    39288 => -19174,
    39289 => -19177,
    39290 => -19180,
    39291 => -19182,
    39292 => -19185,
    39293 => -19187,
    39294 => -19190,
    39295 => -19192,
    39296 => -19195,
    39297 => -19197,
    39298 => -19200,
    39299 => -19202,
    39300 => -19205,
    39301 => -19208,
    39302 => -19210,
    39303 => -19213,
    39304 => -19215,
    39305 => -19218,
    39306 => -19220,
    39307 => -19223,
    39308 => -19225,
    39309 => -19228,
    39310 => -19230,
    39311 => -19233,
    39312 => -19236,
    39313 => -19238,
    39314 => -19241,
    39315 => -19243,
    39316 => -19246,
    39317 => -19248,
    39318 => -19251,
    39319 => -19253,
    39320 => -19256,
    39321 => -19258,
    39322 => -19261,
    39323 => -19264,
    39324 => -19266,
    39325 => -19269,
    39326 => -19271,
    39327 => -19274,
    39328 => -19276,
    39329 => -19279,
    39330 => -19281,
    39331 => -19284,
    39332 => -19286,
    39333 => -19289,
    39334 => -19291,
    39335 => -19294,
    39336 => -19297,
    39337 => -19299,
    39338 => -19302,
    39339 => -19304,
    39340 => -19307,
    39341 => -19309,
    39342 => -19312,
    39343 => -19314,
    39344 => -19317,
    39345 => -19319,
    39346 => -19322,
    39347 => -19324,
    39348 => -19327,
    39349 => -19330,
    39350 => -19332,
    39351 => -19335,
    39352 => -19337,
    39353 => -19340,
    39354 => -19342,
    39355 => -19345,
    39356 => -19347,
    39357 => -19350,
    39358 => -19352,
    39359 => -19355,
    39360 => -19357,
    39361 => -19360,
    39362 => -19362,
    39363 => -19365,
    39364 => -19368,
    39365 => -19370,
    39366 => -19373,
    39367 => -19375,
    39368 => -19378,
    39369 => -19380,
    39370 => -19383,
    39371 => -19385,
    39372 => -19388,
    39373 => -19390,
    39374 => -19393,
    39375 => -19395,
    39376 => -19398,
    39377 => -19400,
    39378 => -19403,
    39379 => -19406,
    39380 => -19408,
    39381 => -19411,
    39382 => -19413,
    39383 => -19416,
    39384 => -19418,
    39385 => -19421,
    39386 => -19423,
    39387 => -19426,
    39388 => -19428,
    39389 => -19431,
    39390 => -19433,
    39391 => -19436,
    39392 => -19438,
    39393 => -19441,
    39394 => -19444,
    39395 => -19446,
    39396 => -19449,
    39397 => -19451,
    39398 => -19454,
    39399 => -19456,
    39400 => -19459,
    39401 => -19461,
    39402 => -19464,
    39403 => -19466,
    39404 => -19469,
    39405 => -19471,
    39406 => -19474,
    39407 => -19476,
    39408 => -19479,
    39409 => -19481,
    39410 => -19484,
    39411 => -19486,
    39412 => -19489,
    39413 => -19492,
    39414 => -19494,
    39415 => -19497,
    39416 => -19499,
    39417 => -19502,
    39418 => -19504,
    39419 => -19507,
    39420 => -19509,
    39421 => -19512,
    39422 => -19514,
    39423 => -19517,
    39424 => -19519,
    39425 => -19522,
    39426 => -19524,
    39427 => -19527,
    39428 => -19529,
    39429 => -19532,
    39430 => -19534,
    39431 => -19537,
    39432 => -19539,
    39433 => -19542,
    39434 => -19545,
    39435 => -19547,
    39436 => -19550,
    39437 => -19552,
    39438 => -19555,
    39439 => -19557,
    39440 => -19560,
    39441 => -19562,
    39442 => -19565,
    39443 => -19567,
    39444 => -19570,
    39445 => -19572,
    39446 => -19575,
    39447 => -19577,
    39448 => -19580,
    39449 => -19582,
    39450 => -19585,
    39451 => -19587,
    39452 => -19590,
    39453 => -19592,
    39454 => -19595,
    39455 => -19597,
    39456 => -19600,
    39457 => -19602,
    39458 => -19605,
    39459 => -19607,
    39460 => -19610,
    39461 => -19613,
    39462 => -19615,
    39463 => -19618,
    39464 => -19620,
    39465 => -19623,
    39466 => -19625,
    39467 => -19628,
    39468 => -19630,
    39469 => -19633,
    39470 => -19635,
    39471 => -19638,
    39472 => -19640,
    39473 => -19643,
    39474 => -19645,
    39475 => -19648,
    39476 => -19650,
    39477 => -19653,
    39478 => -19655,
    39479 => -19658,
    39480 => -19660,
    39481 => -19663,
    39482 => -19665,
    39483 => -19668,
    39484 => -19670,
    39485 => -19673,
    39486 => -19675,
    39487 => -19678,
    39488 => -19680,
    39489 => -19683,
    39490 => -19685,
    39491 => -19688,
    39492 => -19690,
    39493 => -19693,
    39494 => -19695,
    39495 => -19698,
    39496 => -19700,
    39497 => -19703,
    39498 => -19706,
    39499 => -19708,
    39500 => -19711,
    39501 => -19713,
    39502 => -19716,
    39503 => -19718,
    39504 => -19721,
    39505 => -19723,
    39506 => -19726,
    39507 => -19728,
    39508 => -19731,
    39509 => -19733,
    39510 => -19736,
    39511 => -19738,
    39512 => -19741,
    39513 => -19743,
    39514 => -19746,
    39515 => -19748,
    39516 => -19751,
    39517 => -19753,
    39518 => -19756,
    39519 => -19758,
    39520 => -19761,
    39521 => -19763,
    39522 => -19766,
    39523 => -19768,
    39524 => -19771,
    39525 => -19773,
    39526 => -19776,
    39527 => -19778,
    39528 => -19781,
    39529 => -19783,
    39530 => -19786,
    39531 => -19788,
    39532 => -19791,
    39533 => -19793,
    39534 => -19796,
    39535 => -19798,
    39536 => -19801,
    39537 => -19803,
    39538 => -19806,
    39539 => -19808,
    39540 => -19811,
    39541 => -19813,
    39542 => -19816,
    39543 => -19818,
    39544 => -19821,
    39545 => -19823,
    39546 => -19826,
    39547 => -19828,
    39548 => -19831,
    39549 => -19833,
    39550 => -19836,
    39551 => -19838,
    39552 => -19841,
    39553 => -19843,
    39554 => -19846,
    39555 => -19848,
    39556 => -19851,
    39557 => -19853,
    39558 => -19856,
    39559 => -19858,
    39560 => -19861,
    39561 => -19863,
    39562 => -19866,
    39563 => -19868,
    39564 => -19871,
    39565 => -19873,
    39566 => -19876,
    39567 => -19878,
    39568 => -19881,
    39569 => -19883,
    39570 => -19886,
    39571 => -19888,
    39572 => -19891,
    39573 => -19893,
    39574 => -19896,
    39575 => -19898,
    39576 => -19901,
    39577 => -19903,
    39578 => -19906,
    39579 => -19908,
    39580 => -19911,
    39581 => -19913,
    39582 => -19916,
    39583 => -19918,
    39584 => -19921,
    39585 => -19923,
    39586 => -19926,
    39587 => -19928,
    39588 => -19931,
    39589 => -19933,
    39590 => -19936,
    39591 => -19938,
    39592 => -19941,
    39593 => -19943,
    39594 => -19946,
    39595 => -19948,
    39596 => -19951,
    39597 => -19953,
    39598 => -19956,
    39599 => -19958,
    39600 => -19961,
    39601 => -19963,
    39602 => -19966,
    39603 => -19968,
    39604 => -19971,
    39605 => -19973,
    39606 => -19976,
    39607 => -19978,
    39608 => -19981,
    39609 => -19983,
    39610 => -19985,
    39611 => -19988,
    39612 => -19990,
    39613 => -19993,
    39614 => -19995,
    39615 => -19998,
    39616 => -20000,
    39617 => -20003,
    39618 => -20005,
    39619 => -20008,
    39620 => -20010,
    39621 => -20013,
    39622 => -20015,
    39623 => -20018,
    39624 => -20020,
    39625 => -20023,
    39626 => -20025,
    39627 => -20028,
    39628 => -20030,
    39629 => -20033,
    39630 => -20035,
    39631 => -20038,
    39632 => -20040,
    39633 => -20043,
    39634 => -20045,
    39635 => -20048,
    39636 => -20050,
    39637 => -20053,
    39638 => -20055,
    39639 => -20058,
    39640 => -20060,
    39641 => -20063,
    39642 => -20065,
    39643 => -20068,
    39644 => -20070,
    39645 => -20072,
    39646 => -20075,
    39647 => -20077,
    39648 => -20080,
    39649 => -20082,
    39650 => -20085,
    39651 => -20087,
    39652 => -20090,
    39653 => -20092,
    39654 => -20095,
    39655 => -20097,
    39656 => -20100,
    39657 => -20102,
    39658 => -20105,
    39659 => -20107,
    39660 => -20110,
    39661 => -20112,
    39662 => -20115,
    39663 => -20117,
    39664 => -20120,
    39665 => -20122,
    39666 => -20125,
    39667 => -20127,
    39668 => -20130,
    39669 => -20132,
    39670 => -20135,
    39671 => -20137,
    39672 => -20139,
    39673 => -20142,
    39674 => -20144,
    39675 => -20147,
    39676 => -20149,
    39677 => -20152,
    39678 => -20154,
    39679 => -20157,
    39680 => -20159,
    39681 => -20162,
    39682 => -20164,
    39683 => -20167,
    39684 => -20169,
    39685 => -20172,
    39686 => -20174,
    39687 => -20177,
    39688 => -20179,
    39689 => -20182,
    39690 => -20184,
    39691 => -20187,
    39692 => -20189,
    39693 => -20191,
    39694 => -20194,
    39695 => -20196,
    39696 => -20199,
    39697 => -20201,
    39698 => -20204,
    39699 => -20206,
    39700 => -20209,
    39701 => -20211,
    39702 => -20214,
    39703 => -20216,
    39704 => -20219,
    39705 => -20221,
    39706 => -20224,
    39707 => -20226,
    39708 => -20229,
    39709 => -20231,
    39710 => -20234,
    39711 => -20236,
    39712 => -20238,
    39713 => -20241,
    39714 => -20243,
    39715 => -20246,
    39716 => -20248,
    39717 => -20251,
    39718 => -20253,
    39719 => -20256,
    39720 => -20258,
    39721 => -20261,
    39722 => -20263,
    39723 => -20266,
    39724 => -20268,
    39725 => -20271,
    39726 => -20273,
    39727 => -20275,
    39728 => -20278,
    39729 => -20280,
    39730 => -20283,
    39731 => -20285,
    39732 => -20288,
    39733 => -20290,
    39734 => -20293,
    39735 => -20295,
    39736 => -20298,
    39737 => -20300,
    39738 => -20303,
    39739 => -20305,
    39740 => -20308,
    39741 => -20310,
    39742 => -20312,
    39743 => -20315,
    39744 => -20317,
    39745 => -20320,
    39746 => -20322,
    39747 => -20325,
    39748 => -20327,
    39749 => -20330,
    39750 => -20332,
    39751 => -20335,
    39752 => -20337,
    39753 => -20340,
    39754 => -20342,
    39755 => -20345,
    39756 => -20347,
    39757 => -20349,
    39758 => -20352,
    39759 => -20354,
    39760 => -20357,
    39761 => -20359,
    39762 => -20362,
    39763 => -20364,
    39764 => -20367,
    39765 => -20369,
    39766 => -20372,
    39767 => -20374,
    39768 => -20377,
    39769 => -20379,
    39770 => -20381,
    39771 => -20384,
    39772 => -20386,
    39773 => -20389,
    39774 => -20391,
    39775 => -20394,
    39776 => -20396,
    39777 => -20399,
    39778 => -20401,
    39779 => -20404,
    39780 => -20406,
    39781 => -20408,
    39782 => -20411,
    39783 => -20413,
    39784 => -20416,
    39785 => -20418,
    39786 => -20421,
    39787 => -20423,
    39788 => -20426,
    39789 => -20428,
    39790 => -20431,
    39791 => -20433,
    39792 => -20436,
    39793 => -20438,
    39794 => -20440,
    39795 => -20443,
    39796 => -20445,
    39797 => -20448,
    39798 => -20450,
    39799 => -20453,
    39800 => -20455,
    39801 => -20458,
    39802 => -20460,
    39803 => -20463,
    39804 => -20465,
    39805 => -20467,
    39806 => -20470,
    39807 => -20472,
    39808 => -20475,
    39809 => -20477,
    39810 => -20480,
    39811 => -20482,
    39812 => -20485,
    39813 => -20487,
    39814 => -20489,
    39815 => -20492,
    39816 => -20494,
    39817 => -20497,
    39818 => -20499,
    39819 => -20502,
    39820 => -20504,
    39821 => -20507,
    39822 => -20509,
    39823 => -20512,
    39824 => -20514,
    39825 => -20516,
    39826 => -20519,
    39827 => -20521,
    39828 => -20524,
    39829 => -20526,
    39830 => -20529,
    39831 => -20531,
    39832 => -20534,
    39833 => -20536,
    39834 => -20538,
    39835 => -20541,
    39836 => -20543,
    39837 => -20546,
    39838 => -20548,
    39839 => -20551,
    39840 => -20553,
    39841 => -20556,
    39842 => -20558,
    39843 => -20560,
    39844 => -20563,
    39845 => -20565,
    39846 => -20568,
    39847 => -20570,
    39848 => -20573,
    39849 => -20575,
    39850 => -20578,
    39851 => -20580,
    39852 => -20583,
    39853 => -20585,
    39854 => -20587,
    39855 => -20590,
    39856 => -20592,
    39857 => -20595,
    39858 => -20597,
    39859 => -20600,
    39860 => -20602,
    39861 => -20604,
    39862 => -20607,
    39863 => -20609,
    39864 => -20612,
    39865 => -20614,
    39866 => -20617,
    39867 => -20619,
    39868 => -20622,
    39869 => -20624,
    39870 => -20626,
    39871 => -20629,
    39872 => -20631,
    39873 => -20634,
    39874 => -20636,
    39875 => -20639,
    39876 => -20641,
    39877 => -20644,
    39878 => -20646,
    39879 => -20648,
    39880 => -20651,
    39881 => -20653,
    39882 => -20656,
    39883 => -20658,
    39884 => -20661,
    39885 => -20663,
    39886 => -20666,
    39887 => -20668,
    39888 => -20670,
    39889 => -20673,
    39890 => -20675,
    39891 => -20678,
    39892 => -20680,
    39893 => -20683,
    39894 => -20685,
    39895 => -20687,
    39896 => -20690,
    39897 => -20692,
    39898 => -20695,
    39899 => -20697,
    39900 => -20700,
    39901 => -20702,
    39902 => -20704,
    39903 => -20707,
    39904 => -20709,
    39905 => -20712,
    39906 => -20714,
    39907 => -20717,
    39908 => -20719,
    39909 => -20722,
    39910 => -20724,
    39911 => -20726,
    39912 => -20729,
    39913 => -20731,
    39914 => -20734,
    39915 => -20736,
    39916 => -20739,
    39917 => -20741,
    39918 => -20743,
    39919 => -20746,
    39920 => -20748,
    39921 => -20751,
    39922 => -20753,
    39923 => -20756,
    39924 => -20758,
    39925 => -20760,
    39926 => -20763,
    39927 => -20765,
    39928 => -20768,
    39929 => -20770,
    39930 => -20773,
    39931 => -20775,
    39932 => -20777,
    39933 => -20780,
    39934 => -20782,
    39935 => -20785,
    39936 => -20787,
    39937 => -20790,
    39938 => -20792,
    39939 => -20794,
    39940 => -20797,
    39941 => -20799,
    39942 => -20802,
    39943 => -20804,
    39944 => -20807,
    39945 => -20809,
    39946 => -20811,
    39947 => -20814,
    39948 => -20816,
    39949 => -20819,
    39950 => -20821,
    39951 => -20824,
    39952 => -20826,
    39953 => -20828,
    39954 => -20831,
    39955 => -20833,
    39956 => -20836,
    39957 => -20838,
    39958 => -20841,
    39959 => -20843,
    39960 => -20845,
    39961 => -20848,
    39962 => -20850,
    39963 => -20853,
    39964 => -20855,
    39965 => -20858,
    39966 => -20860,
    39967 => -20862,
    39968 => -20865,
    39969 => -20867,
    39970 => -20870,
    39971 => -20872,
    39972 => -20874,
    39973 => -20877,
    39974 => -20879,
    39975 => -20882,
    39976 => -20884,
    39977 => -20887,
    39978 => -20889,
    39979 => -20891,
    39980 => -20894,
    39981 => -20896,
    39982 => -20899,
    39983 => -20901,
    39984 => -20904,
    39985 => -20906,
    39986 => -20908,
    39987 => -20911,
    39988 => -20913,
    39989 => -20916,
    39990 => -20918,
    39991 => -20920,
    39992 => -20923,
    39993 => -20925,
    39994 => -20928,
    39995 => -20930,
    39996 => -20933,
    39997 => -20935,
    39998 => -20937,
    39999 => -20940,
    40000 => -20942,
    40001 => -20945,
    40002 => -20947,
    40003 => -20949,
    40004 => -20952,
    40005 => -20954,
    40006 => -20957,
    40007 => -20959,
    40008 => -20962,
    40009 => -20964,
    40010 => -20966,
    40011 => -20969,
    40012 => -20971,
    40013 => -20974,
    40014 => -20976,
    40015 => -20978,
    40016 => -20981,
    40017 => -20983,
    40018 => -20986,
    40019 => -20988,
    40020 => -20990,
    40021 => -20993,
    40022 => -20995,
    40023 => -20998,
    40024 => -21000,
    40025 => -21003,
    40026 => -21005,
    40027 => -21007,
    40028 => -21010,
    40029 => -21012,
    40030 => -21015,
    40031 => -21017,
    40032 => -21019,
    40033 => -21022,
    40034 => -21024,
    40035 => -21027,
    40036 => -21029,
    40037 => -21031,
    40038 => -21034,
    40039 => -21036,
    40040 => -21039,
    40041 => -21041,
    40042 => -21043,
    40043 => -21046,
    40044 => -21048,
    40045 => -21051,
    40046 => -21053,
    40047 => -21056,
    40048 => -21058,
    40049 => -21060,
    40050 => -21063,
    40051 => -21065,
    40052 => -21068,
    40053 => -21070,
    40054 => -21072,
    40055 => -21075,
    40056 => -21077,
    40057 => -21080,
    40058 => -21082,
    40059 => -21084,
    40060 => -21087,
    40061 => -21089,
    40062 => -21092,
    40063 => -21094,
    40064 => -21096,
    40065 => -21099,
    40066 => -21101,
    40067 => -21104,
    40068 => -21106,
    40069 => -21108,
    40070 => -21111,
    40071 => -21113,
    40072 => -21116,
    40073 => -21118,
    40074 => -21120,
    40075 => -21123,
    40076 => -21125,
    40077 => -21128,
    40078 => -21130,
    40079 => -21132,
    40080 => -21135,
    40081 => -21137,
    40082 => -21140,
    40083 => -21142,
    40084 => -21144,
    40085 => -21147,
    40086 => -21149,
    40087 => -21152,
    40088 => -21154,
    40089 => -21156,
    40090 => -21159,
    40091 => -21161,
    40092 => -21164,
    40093 => -21166,
    40094 => -21168,
    40095 => -21171,
    40096 => -21173,
    40097 => -21176,
    40098 => -21178,
    40099 => -21180,
    40100 => -21183,
    40101 => -21185,
    40102 => -21188,
    40103 => -21190,
    40104 => -21192,
    40105 => -21195,
    40106 => -21197,
    40107 => -21200,
    40108 => -21202,
    40109 => -21204,
    40110 => -21207,
    40111 => -21209,
    40112 => -21212,
    40113 => -21214,
    40114 => -21216,
    40115 => -21219,
    40116 => -21221,
    40117 => -21224,
    40118 => -21226,
    40119 => -21228,
    40120 => -21231,
    40121 => -21233,
    40122 => -21236,
    40123 => -21238,
    40124 => -21240,
    40125 => -21243,
    40126 => -21245,
    40127 => -21247,
    40128 => -21250,
    40129 => -21252,
    40130 => -21255,
    40131 => -21257,
    40132 => -21259,
    40133 => -21262,
    40134 => -21264,
    40135 => -21267,
    40136 => -21269,
    40137 => -21271,
    40138 => -21274,
    40139 => -21276,
    40140 => -21279,
    40141 => -21281,
    40142 => -21283,
    40143 => -21286,
    40144 => -21288,
    40145 => -21290,
    40146 => -21293,
    40147 => -21295,
    40148 => -21298,
    40149 => -21300,
    40150 => -21302,
    40151 => -21305,
    40152 => -21307,
    40153 => -21310,
    40154 => -21312,
    40155 => -21314,
    40156 => -21317,
    40157 => -21319,
    40158 => -21322,
    40159 => -21324,
    40160 => -21326,
    40161 => -21329,
    40162 => -21331,
    40163 => -21333,
    40164 => -21336,
    40165 => -21338,
    40166 => -21341,
    40167 => -21343,
    40168 => -21345,
    40169 => -21348,
    40170 => -21350,
    40171 => -21353,
    40172 => -21355,
    40173 => -21357,
    40174 => -21360,
    40175 => -21362,
    40176 => -21364,
    40177 => -21367,
    40178 => -21369,
    40179 => -21372,
    40180 => -21374,
    40181 => -21376,
    40182 => -21379,
    40183 => -21381,
    40184 => -21383,
    40185 => -21386,
    40186 => -21388,
    40187 => -21391,
    40188 => -21393,
    40189 => -21395,
    40190 => -21398,
    40191 => -21400,
    40192 => -21403,
    40193 => -21405,
    40194 => -21407,
    40195 => -21410,
    40196 => -21412,
    40197 => -21414,
    40198 => -21417,
    40199 => -21419,
    40200 => -21422,
    40201 => -21424,
    40202 => -21426,
    40203 => -21429,
    40204 => -21431,
    40205 => -21433,
    40206 => -21436,
    40207 => -21438,
    40208 => -21441,
    40209 => -21443,
    40210 => -21445,
    40211 => -21448,
    40212 => -21450,
    40213 => -21452,
    40214 => -21455,
    40215 => -21457,
    40216 => -21460,
    40217 => -21462,
    40218 => -21464,
    40219 => -21467,
    40220 => -21469,
    40221 => -21471,
    40222 => -21474,
    40223 => -21476,
    40224 => -21479,
    40225 => -21481,
    40226 => -21483,
    40227 => -21486,
    40228 => -21488,
    40229 => -21490,
    40230 => -21493,
    40231 => -21495,
    40232 => -21498,
    40233 => -21500,
    40234 => -21502,
    40235 => -21505,
    40236 => -21507,
    40237 => -21509,
    40238 => -21512,
    40239 => -21514,
    40240 => -21516,
    40241 => -21519,
    40242 => -21521,
    40243 => -21524,
    40244 => -21526,
    40245 => -21528,
    40246 => -21531,
    40247 => -21533,
    40248 => -21535,
    40249 => -21538,
    40250 => -21540,
    40251 => -21543,
    40252 => -21545,
    40253 => -21547,
    40254 => -21550,
    40255 => -21552,
    40256 => -21554,
    40257 => -21557,
    40258 => -21559,
    40259 => -21561,
    40260 => -21564,
    40261 => -21566,
    40262 => -21569,
    40263 => -21571,
    40264 => -21573,
    40265 => -21576,
    40266 => -21578,
    40267 => -21580,
    40268 => -21583,
    40269 => -21585,
    40270 => -21587,
    40271 => -21590,
    40272 => -21592,
    40273 => -21595,
    40274 => -21597,
    40275 => -21599,
    40276 => -21602,
    40277 => -21604,
    40278 => -21606,
    40279 => -21609,
    40280 => -21611,
    40281 => -21613,
    40282 => -21616,
    40283 => -21618,
    40284 => -21621,
    40285 => -21623,
    40286 => -21625,
    40287 => -21628,
    40288 => -21630,
    40289 => -21632,
    40290 => -21635,
    40291 => -21637,
    40292 => -21639,
    40293 => -21642,
    40294 => -21644,
    40295 => -21646,
    40296 => -21649,
    40297 => -21651,
    40298 => -21654,
    40299 => -21656,
    40300 => -21658,
    40301 => -21661,
    40302 => -21663,
    40303 => -21665,
    40304 => -21668,
    40305 => -21670,
    40306 => -21672,
    40307 => -21675,
    40308 => -21677,
    40309 => -21679,
    40310 => -21682,
    40311 => -21684,
    40312 => -21687,
    40313 => -21689,
    40314 => -21691,
    40315 => -21694,
    40316 => -21696,
    40317 => -21698,
    40318 => -21701,
    40319 => -21703,
    40320 => -21705,
    40321 => -21708,
    40322 => -21710,
    40323 => -21712,
    40324 => -21715,
    40325 => -21717,
    40326 => -21719,
    40327 => -21722,
    40328 => -21724,
    40329 => -21727,
    40330 => -21729,
    40331 => -21731,
    40332 => -21734,
    40333 => -21736,
    40334 => -21738,
    40335 => -21741,
    40336 => -21743,
    40337 => -21745,
    40338 => -21748,
    40339 => -21750,
    40340 => -21752,
    40341 => -21755,
    40342 => -21757,
    40343 => -21759,
    40344 => -21762,
    40345 => -21764,
    40346 => -21766,
    40347 => -21769,
    40348 => -21771,
    40349 => -21774,
    40350 => -21776,
    40351 => -21778,
    40352 => -21781,
    40353 => -21783,
    40354 => -21785,
    40355 => -21788,
    40356 => -21790,
    40357 => -21792,
    40358 => -21795,
    40359 => -21797,
    40360 => -21799,
    40361 => -21802,
    40362 => -21804,
    40363 => -21806,
    40364 => -21809,
    40365 => -21811,
    40366 => -21813,
    40367 => -21816,
    40368 => -21818,
    40369 => -21820,
    40370 => -21823,
    40371 => -21825,
    40372 => -21827,
    40373 => -21830,
    40374 => -21832,
    40375 => -21835,
    40376 => -21837,
    40377 => -21839,
    40378 => -21842,
    40379 => -21844,
    40380 => -21846,
    40381 => -21849,
    40382 => -21851,
    40383 => -21853,
    40384 => -21856,
    40385 => -21858,
    40386 => -21860,
    40387 => -21863,
    40388 => -21865,
    40389 => -21867,
    40390 => -21870,
    40391 => -21872,
    40392 => -21874,
    40393 => -21877,
    40394 => -21879,
    40395 => -21881,
    40396 => -21884,
    40397 => -21886,
    40398 => -21888,
    40399 => -21891,
    40400 => -21893,
    40401 => -21895,
    40402 => -21898,
    40403 => -21900,
    40404 => -21902,
    40405 => -21905,
    40406 => -21907,
    40407 => -21909,
    40408 => -21912,
    40409 => -21914,
    40410 => -21916,
    40411 => -21919,
    40412 => -21921,
    40413 => -21923,
    40414 => -21926,
    40415 => -21928,
    40416 => -21930,
    40417 => -21933,
    40418 => -21935,
    40419 => -21937,
    40420 => -21940,
    40421 => -21942,
    40422 => -21944,
    40423 => -21947,
    40424 => -21949,
    40425 => -21951,
    40426 => -21954,
    40427 => -21956,
    40428 => -21958,
    40429 => -21961,
    40430 => -21963,
    40431 => -21965,
    40432 => -21968,
    40433 => -21970,
    40434 => -21972,
    40435 => -21975,
    40436 => -21977,
    40437 => -21979,
    40438 => -21982,
    40439 => -21984,
    40440 => -21986,
    40441 => -21989,
    40442 => -21991,
    40443 => -21993,
    40444 => -21996,
    40445 => -21998,
    40446 => -22000,
    40447 => -22003,
    40448 => -22005,
    40449 => -22007,
    40450 => -22010,
    40451 => -22012,
    40452 => -22014,
    40453 => -22017,
    40454 => -22019,
    40455 => -22021,
    40456 => -22024,
    40457 => -22026,
    40458 => -22028,
    40459 => -22031,
    40460 => -22033,
    40461 => -22035,
    40462 => -22038,
    40463 => -22040,
    40464 => -22042,
    40465 => -22045,
    40466 => -22047,
    40467 => -22049,
    40468 => -22051,
    40469 => -22054,
    40470 => -22056,
    40471 => -22058,
    40472 => -22061,
    40473 => -22063,
    40474 => -22065,
    40475 => -22068,
    40476 => -22070,
    40477 => -22072,
    40478 => -22075,
    40479 => -22077,
    40480 => -22079,
    40481 => -22082,
    40482 => -22084,
    40483 => -22086,
    40484 => -22089,
    40485 => -22091,
    40486 => -22093,
    40487 => -22096,
    40488 => -22098,
    40489 => -22100,
    40490 => -22103,
    40491 => -22105,
    40492 => -22107,
    40493 => -22110,
    40494 => -22112,
    40495 => -22114,
    40496 => -22116,
    40497 => -22119,
    40498 => -22121,
    40499 => -22123,
    40500 => -22126,
    40501 => -22128,
    40502 => -22130,
    40503 => -22133,
    40504 => -22135,
    40505 => -22137,
    40506 => -22140,
    40507 => -22142,
    40508 => -22144,
    40509 => -22147,
    40510 => -22149,
    40511 => -22151,
    40512 => -22154,
    40513 => -22156,
    40514 => -22158,
    40515 => -22160,
    40516 => -22163,
    40517 => -22165,
    40518 => -22167,
    40519 => -22170,
    40520 => -22172,
    40521 => -22174,
    40522 => -22177,
    40523 => -22179,
    40524 => -22181,
    40525 => -22184,
    40526 => -22186,
    40527 => -22188,
    40528 => -22191,
    40529 => -22193,
    40530 => -22195,
    40531 => -22197,
    40532 => -22200,
    40533 => -22202,
    40534 => -22204,
    40535 => -22207,
    40536 => -22209,
    40537 => -22211,
    40538 => -22214,
    40539 => -22216,
    40540 => -22218,
    40541 => -22221,
    40542 => -22223,
    40543 => -22225,
    40544 => -22227,
    40545 => -22230,
    40546 => -22232,
    40547 => -22234,
    40548 => -22237,
    40549 => -22239,
    40550 => -22241,
    40551 => -22244,
    40552 => -22246,
    40553 => -22248,
    40554 => -22251,
    40555 => -22253,
    40556 => -22255,
    40557 => -22257,
    40558 => -22260,
    40559 => -22262,
    40560 => -22264,
    40561 => -22267,
    40562 => -22269,
    40563 => -22271,
    40564 => -22274,
    40565 => -22276,
    40566 => -22278,
    40567 => -22281,
    40568 => -22283,
    40569 => -22285,
    40570 => -22287,
    40571 => -22290,
    40572 => -22292,
    40573 => -22294,
    40574 => -22297,
    40575 => -22299,
    40576 => -22301,
    40577 => -22304,
    40578 => -22306,
    40579 => -22308,
    40580 => -22310,
    40581 => -22313,
    40582 => -22315,
    40583 => -22317,
    40584 => -22320,
    40585 => -22322,
    40586 => -22324,
    40587 => -22327,
    40588 => -22329,
    40589 => -22331,
    40590 => -22333,
    40591 => -22336,
    40592 => -22338,
    40593 => -22340,
    40594 => -22343,
    40595 => -22345,
    40596 => -22347,
    40597 => -22350,
    40598 => -22352,
    40599 => -22354,
    40600 => -22356,
    40601 => -22359,
    40602 => -22361,
    40603 => -22363,
    40604 => -22366,
    40605 => -22368,
    40606 => -22370,
    40607 => -22373,
    40608 => -22375,
    40609 => -22377,
    40610 => -22379,
    40611 => -22382,
    40612 => -22384,
    40613 => -22386,
    40614 => -22389,
    40615 => -22391,
    40616 => -22393,
    40617 => -22395,
    40618 => -22398,
    40619 => -22400,
    40620 => -22402,
    40621 => -22405,
    40622 => -22407,
    40623 => -22409,
    40624 => -22411,
    40625 => -22414,
    40626 => -22416,
    40627 => -22418,
    40628 => -22421,
    40629 => -22423,
    40630 => -22425,
    40631 => -22428,
    40632 => -22430,
    40633 => -22432,
    40634 => -22434,
    40635 => -22437,
    40636 => -22439,
    40637 => -22441,
    40638 => -22444,
    40639 => -22446,
    40640 => -22448,
    40641 => -22450,
    40642 => -22453,
    40643 => -22455,
    40644 => -22457,
    40645 => -22460,
    40646 => -22462,
    40647 => -22464,
    40648 => -22466,
    40649 => -22469,
    40650 => -22471,
    40651 => -22473,
    40652 => -22476,
    40653 => -22478,
    40654 => -22480,
    40655 => -22482,
    40656 => -22485,
    40657 => -22487,
    40658 => -22489,
    40659 => -22492,
    40660 => -22494,
    40661 => -22496,
    40662 => -22498,
    40663 => -22501,
    40664 => -22503,
    40665 => -22505,
    40666 => -22508,
    40667 => -22510,
    40668 => -22512,
    40669 => -22514,
    40670 => -22517,
    40671 => -22519,
    40672 => -22521,
    40673 => -22524,
    40674 => -22526,
    40675 => -22528,
    40676 => -22530,
    40677 => -22533,
    40678 => -22535,
    40679 => -22537,
    40680 => -22540,
    40681 => -22542,
    40682 => -22544,
    40683 => -22546,
    40684 => -22549,
    40685 => -22551,
    40686 => -22553,
    40687 => -22555,
    40688 => -22558,
    40689 => -22560,
    40690 => -22562,
    40691 => -22565,
    40692 => -22567,
    40693 => -22569,
    40694 => -22571,
    40695 => -22574,
    40696 => -22576,
    40697 => -22578,
    40698 => -22581,
    40699 => -22583,
    40700 => -22585,
    40701 => -22587,
    40702 => -22590,
    40703 => -22592,
    40704 => -22594,
    40705 => -22596,
    40706 => -22599,
    40707 => -22601,
    40708 => -22603,
    40709 => -22606,
    40710 => -22608,
    40711 => -22610,
    40712 => -22612,
    40713 => -22615,
    40714 => -22617,
    40715 => -22619,
    40716 => -22621,
    40717 => -22624,
    40718 => -22626,
    40719 => -22628,
    40720 => -22631,
    40721 => -22633,
    40722 => -22635,
    40723 => -22637,
    40724 => -22640,
    40725 => -22642,
    40726 => -22644,
    40727 => -22646,
    40728 => -22649,
    40729 => -22651,
    40730 => -22653,
    40731 => -22656,
    40732 => -22658,
    40733 => -22660,
    40734 => -22662,
    40735 => -22665,
    40736 => -22667,
    40737 => -22669,
    40738 => -22671,
    40739 => -22674,
    40740 => -22676,
    40741 => -22678,
    40742 => -22680,
    40743 => -22683,
    40744 => -22685,
    40745 => -22687,
    40746 => -22690,
    40747 => -22692,
    40748 => -22694,
    40749 => -22696,
    40750 => -22699,
    40751 => -22701,
    40752 => -22703,
    40753 => -22705,
    40754 => -22708,
    40755 => -22710,
    40756 => -22712,
    40757 => -22714,
    40758 => -22717,
    40759 => -22719,
    40760 => -22721,
    40761 => -22724,
    40762 => -22726,
    40763 => -22728,
    40764 => -22730,
    40765 => -22733,
    40766 => -22735,
    40767 => -22737,
    40768 => -22739,
    40769 => -22742,
    40770 => -22744,
    40771 => -22746,
    40772 => -22748,
    40773 => -22751,
    40774 => -22753,
    40775 => -22755,
    40776 => -22757,
    40777 => -22760,
    40778 => -22762,
    40779 => -22764,
    40780 => -22766,
    40781 => -22769,
    40782 => -22771,
    40783 => -22773,
    40784 => -22776,
    40785 => -22778,
    40786 => -22780,
    40787 => -22782,
    40788 => -22785,
    40789 => -22787,
    40790 => -22789,
    40791 => -22791,
    40792 => -22794,
    40793 => -22796,
    40794 => -22798,
    40795 => -22800,
    40796 => -22803,
    40797 => -22805,
    40798 => -22807,
    40799 => -22809,
    40800 => -22812,
    40801 => -22814,
    40802 => -22816,
    40803 => -22818,
    40804 => -22821,
    40805 => -22823,
    40806 => -22825,
    40807 => -22827,
    40808 => -22830,
    40809 => -22832,
    40810 => -22834,
    40811 => -22836,
    40812 => -22839,
    40813 => -22841,
    40814 => -22843,
    40815 => -22845,
    40816 => -22848,
    40817 => -22850,
    40818 => -22852,
    40819 => -22854,
    40820 => -22857,
    40821 => -22859,
    40822 => -22861,
    40823 => -22863,
    40824 => -22866,
    40825 => -22868,
    40826 => -22870,
    40827 => -22872,
    40828 => -22875,
    40829 => -22877,
    40830 => -22879,
    40831 => -22881,
    40832 => -22884,
    40833 => -22886,
    40834 => -22888,
    40835 => -22890,
    40836 => -22893,
    40837 => -22895,
    40838 => -22897,
    40839 => -22899,
    40840 => -22902,
    40841 => -22904,
    40842 => -22906,
    40843 => -22908,
    40844 => -22911,
    40845 => -22913,
    40846 => -22915,
    40847 => -22917,
    40848 => -22920,
    40849 => -22922,
    40850 => -22924,
    40851 => -22926,
    40852 => -22929,
    40853 => -22931,
    40854 => -22933,
    40855 => -22935,
    40856 => -22938,
    40857 => -22940,
    40858 => -22942,
    40859 => -22944,
    40860 => -22947,
    40861 => -22949,
    40862 => -22951,
    40863 => -22953,
    40864 => -22956,
    40865 => -22958,
    40866 => -22960,
    40867 => -22962,
    40868 => -22965,
    40869 => -22967,
    40870 => -22969,
    40871 => -22971,
    40872 => -22973,
    40873 => -22976,
    40874 => -22978,
    40875 => -22980,
    40876 => -22982,
    40877 => -22985,
    40878 => -22987,
    40879 => -22989,
    40880 => -22991,
    40881 => -22994,
    40882 => -22996,
    40883 => -22998,
    40884 => -23000,
    40885 => -23003,
    40886 => -23005,
    40887 => -23007,
    40888 => -23009,
    40889 => -23012,
    40890 => -23014,
    40891 => -23016,
    40892 => -23018,
    40893 => -23020,
    40894 => -23023,
    40895 => -23025,
    40896 => -23027,
    40897 => -23029,
    40898 => -23032,
    40899 => -23034,
    40900 => -23036,
    40901 => -23038,
    40902 => -23041,
    40903 => -23043,
    40904 => -23045,
    40905 => -23047,
    40906 => -23050,
    40907 => -23052,
    40908 => -23054,
    40909 => -23056,
    40910 => -23058,
    40911 => -23061,
    40912 => -23063,
    40913 => -23065,
    40914 => -23067,
    40915 => -23070,
    40916 => -23072,
    40917 => -23074,
    40918 => -23076,
    40919 => -23079,
    40920 => -23081,
    40921 => -23083,
    40922 => -23085,
    40923 => -23087,
    40924 => -23090,
    40925 => -23092,
    40926 => -23094,
    40927 => -23096,
    40928 => -23099,
    40929 => -23101,
    40930 => -23103,
    40931 => -23105,
    40932 => -23107,
    40933 => -23110,
    40934 => -23112,
    40935 => -23114,
    40936 => -23116,
    40937 => -23119,
    40938 => -23121,
    40939 => -23123,
    40940 => -23125,
    40941 => -23128,
    40942 => -23130,
    40943 => -23132,
    40944 => -23134,
    40945 => -23136,
    40946 => -23139,
    40947 => -23141,
    40948 => -23143,
    40949 => -23145,
    40950 => -23148,
    40951 => -23150,
    40952 => -23152,
    40953 => -23154,
    40954 => -23156,
    40955 => -23159,
    40956 => -23161,
    40957 => -23163,
    40958 => -23165,
    40959 => -23168,
    40960 => -23170,
    40961 => -23172,
    40962 => -23174,
    40963 => -23176,
    40964 => -23179,
    40965 => -23181,
    40966 => -23183,
    40967 => -23185,
    40968 => -23188,
    40969 => -23190,
    40970 => -23192,
    40971 => -23194,
    40972 => -23196,
    40973 => -23199,
    40974 => -23201,
    40975 => -23203,
    40976 => -23205,
    40977 => -23208,
    40978 => -23210,
    40979 => -23212,
    40980 => -23214,
    40981 => -23216,
    40982 => -23219,
    40983 => -23221,
    40984 => -23223,
    40985 => -23225,
    40986 => -23227,
    40987 => -23230,
    40988 => -23232,
    40989 => -23234,
    40990 => -23236,
    40991 => -23239,
    40992 => -23241,
    40993 => -23243,
    40994 => -23245,
    40995 => -23247,
    40996 => -23250,
    40997 => -23252,
    40998 => -23254,
    40999 => -23256,
    41000 => -23258,
    41001 => -23261,
    41002 => -23263,
    41003 => -23265,
    41004 => -23267,
    41005 => -23270,
    41006 => -23272,
    41007 => -23274,
    41008 => -23276,
    41009 => -23278,
    41010 => -23281,
    41011 => -23283,
    41012 => -23285,
    41013 => -23287,
    41014 => -23289,
    41015 => -23292,
    41016 => -23294,
    41017 => -23296,
    41018 => -23298,
    41019 => -23300,
    41020 => -23303,
    41021 => -23305,
    41022 => -23307,
    41023 => -23309,
    41024 => -23311,
    41025 => -23314,
    41026 => -23316,
    41027 => -23318,
    41028 => -23320,
    41029 => -23323,
    41030 => -23325,
    41031 => -23327,
    41032 => -23329,
    41033 => -23331,
    41034 => -23334,
    41035 => -23336,
    41036 => -23338,
    41037 => -23340,
    41038 => -23342,
    41039 => -23345,
    41040 => -23347,
    41041 => -23349,
    41042 => -23351,
    41043 => -23353,
    41044 => -23356,
    41045 => -23358,
    41046 => -23360,
    41047 => -23362,
    41048 => -23364,
    41049 => -23367,
    41050 => -23369,
    41051 => -23371,
    41052 => -23373,
    41053 => -23375,
    41054 => -23378,
    41055 => -23380,
    41056 => -23382,
    41057 => -23384,
    41058 => -23386,
    41059 => -23389,
    41060 => -23391,
    41061 => -23393,
    41062 => -23395,
    41063 => -23397,
    41064 => -23400,
    41065 => -23402,
    41066 => -23404,
    41067 => -23406,
    41068 => -23408,
    41069 => -23411,
    41070 => -23413,
    41071 => -23415,
    41072 => -23417,
    41073 => -23419,
    41074 => -23422,
    41075 => -23424,
    41076 => -23426,
    41077 => -23428,
    41078 => -23430,
    41079 => -23433,
    41080 => -23435,
    41081 => -23437,
    41082 => -23439,
    41083 => -23441,
    41084 => -23444,
    41085 => -23446,
    41086 => -23448,
    41087 => -23450,
    41088 => -23452,
    41089 => -23455,
    41090 => -23457,
    41091 => -23459,
    41092 => -23461,
    41093 => -23463,
    41094 => -23466,
    41095 => -23468,
    41096 => -23470,
    41097 => -23472,
    41098 => -23474,
    41099 => -23476,
    41100 => -23479,
    41101 => -23481,
    41102 => -23483,
    41103 => -23485,
    41104 => -23487,
    41105 => -23490,
    41106 => -23492,
    41107 => -23494,
    41108 => -23496,
    41109 => -23498,
    41110 => -23501,
    41111 => -23503,
    41112 => -23505,
    41113 => -23507,
    41114 => -23509,
    41115 => -23512,
    41116 => -23514,
    41117 => -23516,
    41118 => -23518,
    41119 => -23520,
    41120 => -23522,
    41121 => -23525,
    41122 => -23527,
    41123 => -23529,
    41124 => -23531,
    41125 => -23533,
    41126 => -23536,
    41127 => -23538,
    41128 => -23540,
    41129 => -23542,
    41130 => -23544,
    41131 => -23546,
    41132 => -23549,
    41133 => -23551,
    41134 => -23553,
    41135 => -23555,
    41136 => -23557,
    41137 => -23560,
    41138 => -23562,
    41139 => -23564,
    41140 => -23566,
    41141 => -23568,
    41142 => -23571,
    41143 => -23573,
    41144 => -23575,
    41145 => -23577,
    41146 => -23579,
    41147 => -23581,
    41148 => -23584,
    41149 => -23586,
    41150 => -23588,
    41151 => -23590,
    41152 => -23592,
    41153 => -23595,
    41154 => -23597,
    41155 => -23599,
    41156 => -23601,
    41157 => -23603,
    41158 => -23605,
    41159 => -23608,
    41160 => -23610,
    41161 => -23612,
    41162 => -23614,
    41163 => -23616,
    41164 => -23618,
    41165 => -23621,
    41166 => -23623,
    41167 => -23625,
    41168 => -23627,
    41169 => -23629,
    41170 => -23632,
    41171 => -23634,
    41172 => -23636,
    41173 => -23638,
    41174 => -23640,
    41175 => -23642,
    41176 => -23645,
    41177 => -23647,
    41178 => -23649,
    41179 => -23651,
    41180 => -23653,
    41181 => -23655,
    41182 => -23658,
    41183 => -23660,
    41184 => -23662,
    41185 => -23664,
    41186 => -23666,
    41187 => -23668,
    41188 => -23671,
    41189 => -23673,
    41190 => -23675,
    41191 => -23677,
    41192 => -23679,
    41193 => -23682,
    41194 => -23684,
    41195 => -23686,
    41196 => -23688,
    41197 => -23690,
    41198 => -23692,
    41199 => -23695,
    41200 => -23697,
    41201 => -23699,
    41202 => -23701,
    41203 => -23703,
    41204 => -23705,
    41205 => -23708,
    41206 => -23710,
    41207 => -23712,
    41208 => -23714,
    41209 => -23716,
    41210 => -23718,
    41211 => -23721,
    41212 => -23723,
    41213 => -23725,
    41214 => -23727,
    41215 => -23729,
    41216 => -23731,
    41217 => -23734,
    41218 => -23736,
    41219 => -23738,
    41220 => -23740,
    41221 => -23742,
    41222 => -23744,
    41223 => -23747,
    41224 => -23749,
    41225 => -23751,
    41226 => -23753,
    41227 => -23755,
    41228 => -23757,
    41229 => -23760,
    41230 => -23762,
    41231 => -23764,
    41232 => -23766,
    41233 => -23768,
    41234 => -23770,
    41235 => -23773,
    41236 => -23775,
    41237 => -23777,
    41238 => -23779,
    41239 => -23781,
    41240 => -23783,
    41241 => -23785,
    41242 => -23788,
    41243 => -23790,
    41244 => -23792,
    41245 => -23794,
    41246 => -23796,
    41247 => -23798,
    41248 => -23801,
    41249 => -23803,
    41250 => -23805,
    41251 => -23807,
    41252 => -23809,
    41253 => -23811,
    41254 => -23814,
    41255 => -23816,
    41256 => -23818,
    41257 => -23820,
    41258 => -23822,
    41259 => -23824,
    41260 => -23827,
    41261 => -23829,
    41262 => -23831,
    41263 => -23833,
    41264 => -23835,
    41265 => -23837,
    41266 => -23839,
    41267 => -23842,
    41268 => -23844,
    41269 => -23846,
    41270 => -23848,
    41271 => -23850,
    41272 => -23852,
    41273 => -23855,
    41274 => -23857,
    41275 => -23859,
    41276 => -23861,
    41277 => -23863,
    41278 => -23865,
    41279 => -23867,
    41280 => -23870,
    41281 => -23872,
    41282 => -23874,
    41283 => -23876,
    41284 => -23878,
    41285 => -23880,
    41286 => -23883,
    41287 => -23885,
    41288 => -23887,
    41289 => -23889,
    41290 => -23891,
    41291 => -23893,
    41292 => -23895,
    41293 => -23898,
    41294 => -23900,
    41295 => -23902,
    41296 => -23904,
    41297 => -23906,
    41298 => -23908,
    41299 => -23910,
    41300 => -23913,
    41301 => -23915,
    41302 => -23917,
    41303 => -23919,
    41304 => -23921,
    41305 => -23923,
    41306 => -23925,
    41307 => -23928,
    41308 => -23930,
    41309 => -23932,
    41310 => -23934,
    41311 => -23936,
    41312 => -23938,
    41313 => -23940,
    41314 => -23943,
    41315 => -23945,
    41316 => -23947,
    41317 => -23949,
    41318 => -23951,
    41319 => -23953,
    41320 => -23956,
    41321 => -23958,
    41322 => -23960,
    41323 => -23962,
    41324 => -23964,
    41325 => -23966,
    41326 => -23968,
    41327 => -23971,
    41328 => -23973,
    41329 => -23975,
    41330 => -23977,
    41331 => -23979,
    41332 => -23981,
    41333 => -23983,
    41334 => -23985,
    41335 => -23988,
    41336 => -23990,
    41337 => -23992,
    41338 => -23994,
    41339 => -23996,
    41340 => -23998,
    41341 => -24000,
    41342 => -24003,
    41343 => -24005,
    41344 => -24007,
    41345 => -24009,
    41346 => -24011,
    41347 => -24013,
    41348 => -24015,
    41349 => -24018,
    41350 => -24020,
    41351 => -24022,
    41352 => -24024,
    41353 => -24026,
    41354 => -24028,
    41355 => -24030,
    41356 => -24033,
    41357 => -24035,
    41358 => -24037,
    41359 => -24039,
    41360 => -24041,
    41361 => -24043,
    41362 => -24045,
    41363 => -24047,
    41364 => -24050,
    41365 => -24052,
    41366 => -24054,
    41367 => -24056,
    41368 => -24058,
    41369 => -24060,
    41370 => -24062,
    41371 => -24065,
    41372 => -24067,
    41373 => -24069,
    41374 => -24071,
    41375 => -24073,
    41376 => -24075,
    41377 => -24077,
    41378 => -24079,
    41379 => -24082,
    41380 => -24084,
    41381 => -24086,
    41382 => -24088,
    41383 => -24090,
    41384 => -24092,
    41385 => -24094,
    41386 => -24096,
    41387 => -24099,
    41388 => -24101,
    41389 => -24103,
    41390 => -24105,
    41391 => -24107,
    41392 => -24109,
    41393 => -24111,
    41394 => -24114,
    41395 => -24116,
    41396 => -24118,
    41397 => -24120,
    41398 => -24122,
    41399 => -24124,
    41400 => -24126,
    41401 => -24128,
    41402 => -24131,
    41403 => -24133,
    41404 => -24135,
    41405 => -24137,
    41406 => -24139,
    41407 => -24141,
    41408 => -24143,
    41409 => -24145,
    41410 => -24148,
    41411 => -24150,
    41412 => -24152,
    41413 => -24154,
    41414 => -24156,
    41415 => -24158,
    41416 => -24160,
    41417 => -24162,
    41418 => -24164,
    41419 => -24167,
    41420 => -24169,
    41421 => -24171,
    41422 => -24173,
    41423 => -24175,
    41424 => -24177,
    41425 => -24179,
    41426 => -24181,
    41427 => -24184,
    41428 => -24186,
    41429 => -24188,
    41430 => -24190,
    41431 => -24192,
    41432 => -24194,
    41433 => -24196,
    41434 => -24198,
    41435 => -24201,
    41436 => -24203,
    41437 => -24205,
    41438 => -24207,
    41439 => -24209,
    41440 => -24211,
    41441 => -24213,
    41442 => -24215,
    41443 => -24217,
    41444 => -24220,
    41445 => -24222,
    41446 => -24224,
    41447 => -24226,
    41448 => -24228,
    41449 => -24230,
    41450 => -24232,
    41451 => -24234,
    41452 => -24237,
    41453 => -24239,
    41454 => -24241,
    41455 => -24243,
    41456 => -24245,
    41457 => -24247,
    41458 => -24249,
    41459 => -24251,
    41460 => -24253,
    41461 => -24256,
    41462 => -24258,
    41463 => -24260,
    41464 => -24262,
    41465 => -24264,
    41466 => -24266,
    41467 => -24268,
    41468 => -24270,
    41469 => -24272,
    41470 => -24275,
    41471 => -24277,
    41472 => -24279,
    41473 => -24281,
    41474 => -24283,
    41475 => -24285,
    41476 => -24287,
    41477 => -24289,
    41478 => -24291,
    41479 => -24294,
    41480 => -24296,
    41481 => -24298,
    41482 => -24300,
    41483 => -24302,
    41484 => -24304,
    41485 => -24306,
    41486 => -24308,
    41487 => -24310,
    41488 => -24312,
    41489 => -24315,
    41490 => -24317,
    41491 => -24319,
    41492 => -24321,
    41493 => -24323,
    41494 => -24325,
    41495 => -24327,
    41496 => -24329,
    41497 => -24331,
    41498 => -24334,
    41499 => -24336,
    41500 => -24338,
    41501 => -24340,
    41502 => -24342,
    41503 => -24344,
    41504 => -24346,
    41505 => -24348,
    41506 => -24350,
    41507 => -24352,
    41508 => -24355,
    41509 => -24357,
    41510 => -24359,
    41511 => -24361,
    41512 => -24363,
    41513 => -24365,
    41514 => -24367,
    41515 => -24369,
    41516 => -24371,
    41517 => -24373,
    41518 => -24376,
    41519 => -24378,
    41520 => -24380,
    41521 => -24382,
    41522 => -24384,
    41523 => -24386,
    41524 => -24388,
    41525 => -24390,
    41526 => -24392,
    41527 => -24394,
    41528 => -24397,
    41529 => -24399,
    41530 => -24401,
    41531 => -24403,
    41532 => -24405,
    41533 => -24407,
    41534 => -24409,
    41535 => -24411,
    41536 => -24413,
    41537 => -24415,
    41538 => -24417,
    41539 => -24420,
    41540 => -24422,
    41541 => -24424,
    41542 => -24426,
    41543 => -24428,
    41544 => -24430,
    41545 => -24432,
    41546 => -24434,
    41547 => -24436,
    41548 => -24438,
    41549 => -24441,
    41550 => -24443,
    41551 => -24445,
    41552 => -24447,
    41553 => -24449,
    41554 => -24451,
    41555 => -24453,
    41556 => -24455,
    41557 => -24457,
    41558 => -24459,
    41559 => -24461,
    41560 => -24464,
    41561 => -24466,
    41562 => -24468,
    41563 => -24470,
    41564 => -24472,
    41565 => -24474,
    41566 => -24476,
    41567 => -24478,
    41568 => -24480,
    41569 => -24482,
    41570 => -24484,
    41571 => -24487,
    41572 => -24489,
    41573 => -24491,
    41574 => -24493,
    41575 => -24495,
    41576 => -24497,
    41577 => -24499,
    41578 => -24501,
    41579 => -24503,
    41580 => -24505,
    41581 => -24507,
    41582 => -24509,
    41583 => -24512,
    41584 => -24514,
    41585 => -24516,
    41586 => -24518,
    41587 => -24520,
    41588 => -24522,
    41589 => -24524,
    41590 => -24526,
    41591 => -24528,
    41592 => -24530,
    41593 => -24532,
    41594 => -24534,
    41595 => -24537,
    41596 => -24539,
    41597 => -24541,
    41598 => -24543,
    41599 => -24545,
    41600 => -24547,
    41601 => -24549,
    41602 => -24551,
    41603 => -24553,
    41604 => -24555,
    41605 => -24557,
    41606 => -24559,
    41607 => -24562,
    41608 => -24564,
    41609 => -24566,
    41610 => -24568,
    41611 => -24570,
    41612 => -24572,
    41613 => -24574,
    41614 => -24576,
    41615 => -24578,
    41616 => -24580,
    41617 => -24582,
    41618 => -24584,
    41619 => -24586,
    41620 => -24589,
    41621 => -24591,
    41622 => -24593,
    41623 => -24595,
    41624 => -24597,
    41625 => -24599,
    41626 => -24601,
    41627 => -24603,
    41628 => -24605,
    41629 => -24607,
    41630 => -24609,
    41631 => -24611,
    41632 => -24613,
    41633 => -24616,
    41634 => -24618,
    41635 => -24620,
    41636 => -24622,
    41637 => -24624,
    41638 => -24626,
    41639 => -24628,
    41640 => -24630,
    41641 => -24632,
    41642 => -24634,
    41643 => -24636,
    41644 => -24638,
    41645 => -24640,
    41646 => -24642,
    41647 => -24645,
    41648 => -24647,
    41649 => -24649,
    41650 => -24651,
    41651 => -24653,
    41652 => -24655,
    41653 => -24657,
    41654 => -24659,
    41655 => -24661,
    41656 => -24663,
    41657 => -24665,
    41658 => -24667,
    41659 => -24669,
    41660 => -24671,
    41661 => -24673,
    41662 => -24676,
    41663 => -24678,
    41664 => -24680,
    41665 => -24682,
    41666 => -24684,
    41667 => -24686,
    41668 => -24688,
    41669 => -24690,
    41670 => -24692,
    41671 => -24694,
    41672 => -24696,
    41673 => -24698,
    41674 => -24700,
    41675 => -24702,
    41676 => -24704,
    41677 => -24707,
    41678 => -24709,
    41679 => -24711,
    41680 => -24713,
    41681 => -24715,
    41682 => -24717,
    41683 => -24719,
    41684 => -24721,
    41685 => -24723,
    41686 => -24725,
    41687 => -24727,
    41688 => -24729,
    41689 => -24731,
    41690 => -24733,
    41691 => -24735,
    41692 => -24737,
    41693 => -24740,
    41694 => -24742,
    41695 => -24744,
    41696 => -24746,
    41697 => -24748,
    41698 => -24750,
    41699 => -24752,
    41700 => -24754,
    41701 => -24756,
    41702 => -24758,
    41703 => -24760,
    41704 => -24762,
    41705 => -24764,
    41706 => -24766,
    41707 => -24768,
    41708 => -24770,
    41709 => -24772,
    41710 => -24774,
    41711 => -24777,
    41712 => -24779,
    41713 => -24781,
    41714 => -24783,
    41715 => -24785,
    41716 => -24787,
    41717 => -24789,
    41718 => -24791,
    41719 => -24793,
    41720 => -24795,
    41721 => -24797,
    41722 => -24799,
    41723 => -24801,
    41724 => -24803,
    41725 => -24805,
    41726 => -24807,
    41727 => -24809,
    41728 => -24811,
    41729 => -24814,
    41730 => -24816,
    41731 => -24818,
    41732 => -24820,
    41733 => -24822,
    41734 => -24824,
    41735 => -24826,
    41736 => -24828,
    41737 => -24830,
    41738 => -24832,
    41739 => -24834,
    41740 => -24836,
    41741 => -24838,
    41742 => -24840,
    41743 => -24842,
    41744 => -24844,
    41745 => -24846,
    41746 => -24848,
    41747 => -24850,
    41748 => -24852,
    41749 => -24855,
    41750 => -24857,
    41751 => -24859,
    41752 => -24861,
    41753 => -24863,
    41754 => -24865,
    41755 => -24867,
    41756 => -24869,
    41757 => -24871,
    41758 => -24873,
    41759 => -24875,
    41760 => -24877,
    41761 => -24879,
    41762 => -24881,
    41763 => -24883,
    41764 => -24885,
    41765 => -24887,
    41766 => -24889,
    41767 => -24891,
    41768 => -24893,
    41769 => -24895,
    41770 => -24897,
    41771 => -24899,
    41772 => -24902,
    41773 => -24904,
    41774 => -24906,
    41775 => -24908,
    41776 => -24910,
    41777 => -24912,
    41778 => -24914,
    41779 => -24916,
    41780 => -24918,
    41781 => -24920,
    41782 => -24922,
    41783 => -24924,
    41784 => -24926,
    41785 => -24928,
    41786 => -24930,
    41787 => -24932,
    41788 => -24934,
    41789 => -24936,
    41790 => -24938,
    41791 => -24940,
    41792 => -24942,
    41793 => -24944,
    41794 => -24946,
    41795 => -24948,
    41796 => -24950,
    41797 => -24953,
    41798 => -24955,
    41799 => -24957,
    41800 => -24959,
    41801 => -24961,
    41802 => -24963,
    41803 => -24965,
    41804 => -24967,
    41805 => -24969,
    41806 => -24971,
    41807 => -24973,
    41808 => -24975,
    41809 => -24977,
    41810 => -24979,
    41811 => -24981,
    41812 => -24983,
    41813 => -24985,
    41814 => -24987,
    41815 => -24989,
    41816 => -24991,
    41817 => -24993,
    41818 => -24995,
    41819 => -24997,
    41820 => -24999,
    41821 => -25001,
    41822 => -25003,
    41823 => -25005,
    41824 => -25007,
    41825 => -25009,
    41826 => -25011,
    41827 => -25013,
    41828 => -25016,
    41829 => -25018,
    41830 => -25020,
    41831 => -25022,
    41832 => -25024,
    41833 => -25026,
    41834 => -25028,
    41835 => -25030,
    41836 => -25032,
    41837 => -25034,
    41838 => -25036,
    41839 => -25038,
    41840 => -25040,
    41841 => -25042,
    41842 => -25044,
    41843 => -25046,
    41844 => -25048,
    41845 => -25050,
    41846 => -25052,
    41847 => -25054,
    41848 => -25056,
    41849 => -25058,
    41850 => -25060,
    41851 => -25062,
    41852 => -25064,
    41853 => -25066,
    41854 => -25068,
    41855 => -25070,
    41856 => -25072,
    41857 => -25074,
    41858 => -25076,
    41859 => -25078,
    41860 => -25080,
    41861 => -25082,
    41862 => -25084,
    41863 => -25086,
    41864 => -25088,
    41865 => -25090,
    41866 => -25092,
    41867 => -25094,
    41868 => -25096,
    41869 => -25099,
    41870 => -25101,
    41871 => -25103,
    41872 => -25105,
    41873 => -25107,
    41874 => -25109,
    41875 => -25111,
    41876 => -25113,
    41877 => -25115,
    41878 => -25117,
    41879 => -25119,
    41880 => -25121,
    41881 => -25123,
    41882 => -25125,
    41883 => -25127,
    41884 => -25129,
    41885 => -25131,
    41886 => -25133,
    41887 => -25135,
    41888 => -25137,
    41889 => -25139,
    41890 => -25141,
    41891 => -25143,
    41892 => -25145,
    41893 => -25147,
    41894 => -25149,
    41895 => -25151,
    41896 => -25153,
    41897 => -25155,
    41898 => -25157,
    41899 => -25159,
    41900 => -25161,
    41901 => -25163,
    41902 => -25165,
    41903 => -25167,
    41904 => -25169,
    41905 => -25171,
    41906 => -25173,
    41907 => -25175,
    41908 => -25177,
    41909 => -25179,
    41910 => -25181,
    41911 => -25183,
    41912 => -25185,
    41913 => -25187,
    41914 => -25189,
    41915 => -25191,
    41916 => -25193,
    41917 => -25195,
    41918 => -25197,
    41919 => -25199,
    41920 => -25201,
    41921 => -25203,
    41922 => -25205,
    41923 => -25207,
    41924 => -25209,
    41925 => -25211,
    41926 => -25213,
    41927 => -25215,
    41928 => -25217,
    41929 => -25219,
    41930 => -25221,
    41931 => -25223,
    41932 => -25225,
    41933 => -25227,
    41934 => -25229,
    41935 => -25231,
    41936 => -25233,
    41937 => -25235,
    41938 => -25237,
    41939 => -25239,
    41940 => -25241,
    41941 => -25243,
    41942 => -25245,
    41943 => -25247,
    41944 => -25249,
    41945 => -25251,
    41946 => -25253,
    41947 => -25255,
    41948 => -25257,
    41949 => -25259,
    41950 => -25261,
    41951 => -25263,
    41952 => -25265,
    41953 => -25267,
    41954 => -25269,
    41955 => -25271,
    41956 => -25273,
    41957 => -25275,
    41958 => -25277,
    41959 => -25279,
    41960 => -25281,
    41961 => -25283,
    41962 => -25285,
    41963 => -25287,
    41964 => -25289,
    41965 => -25291,
    41966 => -25293,
    41967 => -25295,
    41968 => -25297,
    41969 => -25299,
    41970 => -25301,
    41971 => -25303,
    41972 => -25305,
    41973 => -25307,
    41974 => -25309,
    41975 => -25311,
    41976 => -25313,
    41977 => -25315,
    41978 => -25317,
    41979 => -25319,
    41980 => -25321,
    41981 => -25323,
    41982 => -25325,
    41983 => -25327,
    41984 => -25329,
    41985 => -25331,
    41986 => -25333,
    41987 => -25335,
    41988 => -25337,
    41989 => -25339,
    41990 => -25341,
    41991 => -25343,
    41992 => -25345,
    41993 => -25347,
    41994 => -25349,
    41995 => -25351,
    41996 => -25353,
    41997 => -25355,
    41998 => -25357,
    41999 => -25359,
    42000 => -25361,
    42001 => -25363,
    42002 => -25365,
    42003 => -25367,
    42004 => -25369,
    42005 => -25371,
    42006 => -25373,
    42007 => -25375,
    42008 => -25377,
    42009 => -25379,
    42010 => -25381,
    42011 => -25383,
    42012 => -25385,
    42013 => -25387,
    42014 => -25389,
    42015 => -25391,
    42016 => -25393,
    42017 => -25395,
    42018 => -25397,
    42019 => -25399,
    42020 => -25401,
    42021 => -25403,
    42022 => -25405,
    42023 => -25407,
    42024 => -25409,
    42025 => -25411,
    42026 => -25413,
    42027 => -25415,
    42028 => -25417,
    42029 => -25419,
    42030 => -25421,
    42031 => -25423,
    42032 => -25425,
    42033 => -25427,
    42034 => -25429,
    42035 => -25431,
    42036 => -25433,
    42037 => -25435,
    42038 => -25437,
    42039 => -25438,
    42040 => -25440,
    42041 => -25442,
    42042 => -25444,
    42043 => -25446,
    42044 => -25448,
    42045 => -25450,
    42046 => -25452,
    42047 => -25454,
    42048 => -25456,
    42049 => -25458,
    42050 => -25460,
    42051 => -25462,
    42052 => -25464,
    42053 => -25466,
    42054 => -25468,
    42055 => -25470,
    42056 => -25472,
    42057 => -25474,
    42058 => -25476,
    42059 => -25478,
    42060 => -25480,
    42061 => -25482,
    42062 => -25484,
    42063 => -25486,
    42064 => -25488,
    42065 => -25490,
    42066 => -25492,
    42067 => -25494,
    42068 => -25496,
    42069 => -25498,
    42070 => -25500,
    42071 => -25502,
    42072 => -25504,
    42073 => -25506,
    42074 => -25508,
    42075 => -25510,
    42076 => -25512,
    42077 => -25514,
    42078 => -25516,
    42079 => -25518,
    42080 => -25519,
    42081 => -25521,
    42082 => -25523,
    42083 => -25525,
    42084 => -25527,
    42085 => -25529,
    42086 => -25531,
    42087 => -25533,
    42088 => -25535,
    42089 => -25537,
    42090 => -25539,
    42091 => -25541,
    42092 => -25543,
    42093 => -25545,
    42094 => -25547,
    42095 => -25549,
    42096 => -25551,
    42097 => -25553,
    42098 => -25555,
    42099 => -25557,
    42100 => -25559,
    42101 => -25561,
    42102 => -25563,
    42103 => -25565,
    42104 => -25567,
    42105 => -25569,
    42106 => -25571,
    42107 => -25573,
    42108 => -25575,
    42109 => -25577,
    42110 => -25578,
    42111 => -25580,
    42112 => -25582,
    42113 => -25584,
    42114 => -25586,
    42115 => -25588,
    42116 => -25590,
    42117 => -25592,
    42118 => -25594,
    42119 => -25596,
    42120 => -25598,
    42121 => -25600,
    42122 => -25602,
    42123 => -25604,
    42124 => -25606,
    42125 => -25608,
    42126 => -25610,
    42127 => -25612,
    42128 => -25614,
    42129 => -25616,
    42130 => -25618,
    42131 => -25620,
    42132 => -25622,
    42133 => -25624,
    42134 => -25626,
    42135 => -25628,
    42136 => -25629,
    42137 => -25631,
    42138 => -25633,
    42139 => -25635,
    42140 => -25637,
    42141 => -25639,
    42142 => -25641,
    42143 => -25643,
    42144 => -25645,
    42145 => -25647,
    42146 => -25649,
    42147 => -25651,
    42148 => -25653,
    42149 => -25655,
    42150 => -25657,
    42151 => -25659,
    42152 => -25661,
    42153 => -25663,
    42154 => -25665,
    42155 => -25667,
    42156 => -25669,
    42157 => -25671,
    42158 => -25672,
    42159 => -25674,
    42160 => -25676,
    42161 => -25678,
    42162 => -25680,
    42163 => -25682,
    42164 => -25684,
    42165 => -25686,
    42166 => -25688,
    42167 => -25690,
    42168 => -25692,
    42169 => -25694,
    42170 => -25696,
    42171 => -25698,
    42172 => -25700,
    42173 => -25702,
    42174 => -25704,
    42175 => -25706,
    42176 => -25708,
    42177 => -25710,
    42178 => -25711,
    42179 => -25713,
    42180 => -25715,
    42181 => -25717,
    42182 => -25719,
    42183 => -25721,
    42184 => -25723,
    42185 => -25725,
    42186 => -25727,
    42187 => -25729,
    42188 => -25731,
    42189 => -25733,
    42190 => -25735,
    42191 => -25737,
    42192 => -25739,
    42193 => -25741,
    42194 => -25743,
    42195 => -25745,
    42196 => -25746,
    42197 => -25748,
    42198 => -25750,
    42199 => -25752,
    42200 => -25754,
    42201 => -25756,
    42202 => -25758,
    42203 => -25760,
    42204 => -25762,
    42205 => -25764,
    42206 => -25766,
    42207 => -25768,
    42208 => -25770,
    42209 => -25772,
    42210 => -25774,
    42211 => -25776,
    42212 => -25778,
    42213 => -25779,
    42214 => -25781,
    42215 => -25783,
    42216 => -25785,
    42217 => -25787,
    42218 => -25789,
    42219 => -25791,
    42220 => -25793,
    42221 => -25795,
    42222 => -25797,
    42223 => -25799,
    42224 => -25801,
    42225 => -25803,
    42226 => -25805,
    42227 => -25807,
    42228 => -25809,
    42229 => -25810,
    42230 => -25812,
    42231 => -25814,
    42232 => -25816,
    42233 => -25818,
    42234 => -25820,
    42235 => -25822,
    42236 => -25824,
    42237 => -25826,
    42238 => -25828,
    42239 => -25830,
    42240 => -25832,
    42241 => -25834,
    42242 => -25836,
    42243 => -25838,
    42244 => -25839,
    42245 => -25841,
    42246 => -25843,
    42247 => -25845,
    42248 => -25847,
    42249 => -25849,
    42250 => -25851,
    42251 => -25853,
    42252 => -25855,
    42253 => -25857,
    42254 => -25859,
    42255 => -25861,
    42256 => -25863,
    42257 => -25865,
    42258 => -25866,
    42259 => -25868,
    42260 => -25870,
    42261 => -25872,
    42262 => -25874,
    42263 => -25876,
    42264 => -25878,
    42265 => -25880,
    42266 => -25882,
    42267 => -25884,
    42268 => -25886,
    42269 => -25888,
    42270 => -25890,
    42271 => -25892,
    42272 => -25893,
    42273 => -25895,
    42274 => -25897,
    42275 => -25899,
    42276 => -25901,
    42277 => -25903,
    42278 => -25905,
    42279 => -25907,
    42280 => -25909,
    42281 => -25911,
    42282 => -25913,
    42283 => -25915,
    42284 => -25917,
    42285 => -25918,
    42286 => -25920,
    42287 => -25922,
    42288 => -25924,
    42289 => -25926,
    42290 => -25928,
    42291 => -25930,
    42292 => -25932,
    42293 => -25934,
    42294 => -25936,
    42295 => -25938,
    42296 => -25940,
    42297 => -25942,
    42298 => -25943,
    42299 => -25945,
    42300 => -25947,
    42301 => -25949,
    42302 => -25951,
    42303 => -25953,
    42304 => -25955,
    42305 => -25957,
    42306 => -25959,
    42307 => -25961,
    42308 => -25963,
    42309 => -25965,
    42310 => -25966,
    42311 => -25968,
    42312 => -25970,
    42313 => -25972,
    42314 => -25974,
    42315 => -25976,
    42316 => -25978,
    42317 => -25980,
    42318 => -25982,
    42319 => -25984,
    42320 => -25986,
    42321 => -25988,
    42322 => -25989,
    42323 => -25991,
    42324 => -25993,
    42325 => -25995,
    42326 => -25997,
    42327 => -25999,
    42328 => -26001,
    42329 => -26003,
    42330 => -26005,
    42331 => -26007,
    42332 => -26009,
    42333 => -26010,
    42334 => -26012,
    42335 => -26014,
    42336 => -26016,
    42337 => -26018,
    42338 => -26020,
    42339 => -26022,
    42340 => -26024,
    42341 => -26026,
    42342 => -26028,
    42343 => -26030,
    42344 => -26031,
    42345 => -26033,
    42346 => -26035,
    42347 => -26037,
    42348 => -26039,
    42349 => -26041,
    42350 => -26043,
    42351 => -26045,
    42352 => -26047,
    42353 => -26049,
    42354 => -26051,
    42355 => -26052,
    42356 => -26054,
    42357 => -26056,
    42358 => -26058,
    42359 => -26060,
    42360 => -26062,
    42361 => -26064,
    42362 => -26066,
    42363 => -26068,
    42364 => -26070,
    42365 => -26071,
    42366 => -26073,
    42367 => -26075,
    42368 => -26077,
    42369 => -26079,
    42370 => -26081,
    42371 => -26083,
    42372 => -26085,
    42373 => -26087,
    42374 => -26089,
    42375 => -26090,
    42376 => -26092,
    42377 => -26094,
    42378 => -26096,
    42379 => -26098,
    42380 => -26100,
    42381 => -26102,
    42382 => -26104,
    42383 => -26106,
    42384 => -26108,
    42385 => -26109,
    42386 => -26111,
    42387 => -26113,
    42388 => -26115,
    42389 => -26117,
    42390 => -26119,
    42391 => -26121,
    42392 => -26123,
    42393 => -26125,
    42394 => -26127,
    42395 => -26128,
    42396 => -26130,
    42397 => -26132,
    42398 => -26134,
    42399 => -26136,
    42400 => -26138,
    42401 => -26140,
    42402 => -26142,
    42403 => -26144,
    42404 => -26146,
    42405 => -26147,
    42406 => -26149,
    42407 => -26151,
    42408 => -26153,
    42409 => -26155,
    42410 => -26157,
    42411 => -26159,
    42412 => -26161,
    42413 => -26163,
    42414 => -26164,
    42415 => -26166,
    42416 => -26168,
    42417 => -26170,
    42418 => -26172,
    42419 => -26174,
    42420 => -26176,
    42421 => -26178,
    42422 => -26180,
    42423 => -26181,
    42424 => -26183,
    42425 => -26185,
    42426 => -26187,
    42427 => -26189,
    42428 => -26191,
    42429 => -26193,
    42430 => -26195,
    42431 => -26197,
    42432 => -26198,
    42433 => -26200,
    42434 => -26202,
    42435 => -26204,
    42436 => -26206,
    42437 => -26208,
    42438 => -26210,
    42439 => -26212,
    42440 => -26214,
    42441 => -26215,
    42442 => -26217,
    42443 => -26219,
    42444 => -26221,
    42445 => -26223,
    42446 => -26225,
    42447 => -26227,
    42448 => -26229,
    42449 => -26230,
    42450 => -26232,
    42451 => -26234,
    42452 => -26236,
    42453 => -26238,
    42454 => -26240,
    42455 => -26242,
    42456 => -26244,
    42457 => -26246,
    42458 => -26247,
    42459 => -26249,
    42460 => -26251,
    42461 => -26253,
    42462 => -26255,
    42463 => -26257,
    42464 => -26259,
    42465 => -26261,
    42466 => -26262,
    42467 => -26264,
    42468 => -26266,
    42469 => -26268,
    42470 => -26270,
    42471 => -26272,
    42472 => -26274,
    42473 => -26276,
    42474 => -26277,
    42475 => -26279,
    42476 => -26281,
    42477 => -26283,
    42478 => -26285,
    42479 => -26287,
    42480 => -26289,
    42481 => -26291,
    42482 => -26292,
    42483 => -26294,
    42484 => -26296,
    42485 => -26298,
    42486 => -26300,
    42487 => -26302,
    42488 => -26304,
    42489 => -26306,
    42490 => -26307,
    42491 => -26309,
    42492 => -26311,
    42493 => -26313,
    42494 => -26315,
    42495 => -26317,
    42496 => -26319,
    42497 => -26321,
    42498 => -26322,
    42499 => -26324,
    42500 => -26326,
    42501 => -26328,
    42502 => -26330,
    42503 => -26332,
    42504 => -26334,
    42505 => -26336,
    42506 => -26337,
    42507 => -26339,
    42508 => -26341,
    42509 => -26343,
    42510 => -26345,
    42511 => -26347,
    42512 => -26349,
    42513 => -26350,
    42514 => -26352,
    42515 => -26354,
    42516 => -26356,
    42517 => -26358,
    42518 => -26360,
    42519 => -26362,
    42520 => -26364,
    42521 => -26365,
    42522 => -26367,
    42523 => -26369,
    42524 => -26371,
    42525 => -26373,
    42526 => -26375,
    42527 => -26377,
    42528 => -26378,
    42529 => -26380,
    42530 => -26382,
    42531 => -26384,
    42532 => -26386,
    42533 => -26388,
    42534 => -26390,
    42535 => -26392,
    42536 => -26393,
    42537 => -26395,
    42538 => -26397,
    42539 => -26399,
    42540 => -26401,
    42541 => -26403,
    42542 => -26405,
    42543 => -26406,
    42544 => -26408,
    42545 => -26410,
    42546 => -26412,
    42547 => -26414,
    42548 => -26416,
    42549 => -26418,
    42550 => -26419,
    42551 => -26421,
    42552 => -26423,
    42553 => -26425,
    42554 => -26427,
    42555 => -26429,
    42556 => -26431,
    42557 => -26432,
    42558 => -26434,
    42559 => -26436,
    42560 => -26438,
    42561 => -26440,
    42562 => -26442,
    42563 => -26444,
    42564 => -26445,
    42565 => -26447,
    42566 => -26449,
    42567 => -26451,
    42568 => -26453,
    42569 => -26455,
    42570 => -26457,
    42571 => -26458,
    42572 => -26460,
    42573 => -26462,
    42574 => -26464,
    42575 => -26466,
    42576 => -26468,
    42577 => -26469,
    42578 => -26471,
    42579 => -26473,
    42580 => -26475,
    42581 => -26477,
    42582 => -26479,
    42583 => -26481,
    42584 => -26482,
    42585 => -26484,
    42586 => -26486,
    42587 => -26488,
    42588 => -26490,
    42589 => -26492,
    42590 => -26494,
    42591 => -26495,
    42592 => -26497,
    42593 => -26499,
    42594 => -26501,
    42595 => -26503,
    42596 => -26505,
    42597 => -26506,
    42598 => -26508,
    42599 => -26510,
    42600 => -26512,
    42601 => -26514,
    42602 => -26516,
    42603 => -26518,
    42604 => -26519,
    42605 => -26521,
    42606 => -26523,
    42607 => -26525,
    42608 => -26527,
    42609 => -26529,
    42610 => -26530,
    42611 => -26532,
    42612 => -26534,
    42613 => -26536,
    42614 => -26538,
    42615 => -26540,
    42616 => -26542,
    42617 => -26543,
    42618 => -26545,
    42619 => -26547,
    42620 => -26549,
    42621 => -26551,
    42622 => -26553,
    42623 => -26554,
    42624 => -26556,
    42625 => -26558,
    42626 => -26560,
    42627 => -26562,
    42628 => -26564,
    42629 => -26565,
    42630 => -26567,
    42631 => -26569,
    42632 => -26571,
    42633 => -26573,
    42634 => -26575,
    42635 => -26576,
    42636 => -26578,
    42637 => -26580,
    42638 => -26582,
    42639 => -26584,
    42640 => -26586,
    42641 => -26588,
    42642 => -26589,
    42643 => -26591,
    42644 => -26593,
    42645 => -26595,
    42646 => -26597,
    42647 => -26599,
    42648 => -26600,
    42649 => -26602,
    42650 => -26604,
    42651 => -26606,
    42652 => -26608,
    42653 => -26610,
    42654 => -26611,
    42655 => -26613,
    42656 => -26615,
    42657 => -26617,
    42658 => -26619,
    42659 => -26621,
    42660 => -26622,
    42661 => -26624,
    42662 => -26626,
    42663 => -26628,
    42664 => -26630,
    42665 => -26631,
    42666 => -26633,
    42667 => -26635,
    42668 => -26637,
    42669 => -26639,
    42670 => -26641,
    42671 => -26642,
    42672 => -26644,
    42673 => -26646,
    42674 => -26648,
    42675 => -26650,
    42676 => -26652,
    42677 => -26653,
    42678 => -26655,
    42679 => -26657,
    42680 => -26659,
    42681 => -26661,
    42682 => -26663,
    42683 => -26664,
    42684 => -26666,
    42685 => -26668,
    42686 => -26670,
    42687 => -26672,
    42688 => -26674,
    42689 => -26675,
    42690 => -26677,
    42691 => -26679,
    42692 => -26681,
    42693 => -26683,
    42694 => -26684,
    42695 => -26686,
    42696 => -26688,
    42697 => -26690,
    42698 => -26692,
    42699 => -26694,
    42700 => -26695,
    42701 => -26697,
    42702 => -26699,
    42703 => -26701,
    42704 => -26703,
    42705 => -26705,
    42706 => -26706,
    42707 => -26708,
    42708 => -26710,
    42709 => -26712,
    42710 => -26714,
    42711 => -26715,
    42712 => -26717,
    42713 => -26719,
    42714 => -26721,
    42715 => -26723,
    42716 => -26725,
    42717 => -26726,
    42718 => -26728,
    42719 => -26730,
    42720 => -26732,
    42721 => -26734,
    42722 => -26735,
    42723 => -26737,
    42724 => -26739,
    42725 => -26741,
    42726 => -26743,
    42727 => -26745,
    42728 => -26746,
    42729 => -26748,
    42730 => -26750,
    42731 => -26752,
    42732 => -26754,
    42733 => -26755,
    42734 => -26757,
    42735 => -26759,
    42736 => -26761,
    42737 => -26763,
    42738 => -26764,
    42739 => -26766,
    42740 => -26768,
    42741 => -26770,
    42742 => -26772,
    42743 => -26774,
    42744 => -26775,
    42745 => -26777,
    42746 => -26779,
    42747 => -26781,
    42748 => -26783,
    42749 => -26784,
    42750 => -26786,
    42751 => -26788,
    42752 => -26790,
    42753 => -26792,
    42754 => -26793,
    42755 => -26795,
    42756 => -26797,
    42757 => -26799,
    42758 => -26801,
    42759 => -26802,
    42760 => -26804,
    42761 => -26806,
    42762 => -26808,
    42763 => -26810,
    42764 => -26811,
    42765 => -26813,
    42766 => -26815,
    42767 => -26817,
    42768 => -26819,
    42769 => -26821,
    42770 => -26822,
    42771 => -26824,
    42772 => -26826,
    42773 => -26828,
    42774 => -26830,
    42775 => -26831,
    42776 => -26833,
    42777 => -26835,
    42778 => -26837,
    42779 => -26839,
    42780 => -26840,
    42781 => -26842,
    42782 => -26844,
    42783 => -26846,
    42784 => -26848,
    42785 => -26849,
    42786 => -26851,
    42787 => -26853,
    42788 => -26855,
    42789 => -26857,
    42790 => -26858,
    42791 => -26860,
    42792 => -26862,
    42793 => -26864,
    42794 => -26866,
    42795 => -26867,
    42796 => -26869,
    42797 => -26871,
    42798 => -26873,
    42799 => -26875,
    42800 => -26876,
    42801 => -26878,
    42802 => -26880,
    42803 => -26882,
    42804 => -26884,
    42805 => -26885,
    42806 => -26887,
    42807 => -26889,
    42808 => -26891,
    42809 => -26893,
    42810 => -26894,
    42811 => -26896,
    42812 => -26898,
    42813 => -26900,
    42814 => -26901,
    42815 => -26903,
    42816 => -26905,
    42817 => -26907,
    42818 => -26909,
    42819 => -26910,
    42820 => -26912,
    42821 => -26914,
    42822 => -26916,
    42823 => -26918,
    42824 => -26919,
    42825 => -26921,
    42826 => -26923,
    42827 => -26925,
    42828 => -26927,
    42829 => -26928,
    42830 => -26930,
    42831 => -26932,
    42832 => -26934,
    42833 => -26936,
    42834 => -26937,
    42835 => -26939,
    42836 => -26941,
    42837 => -26943,
    42838 => -26944,
    42839 => -26946,
    42840 => -26948,
    42841 => -26950,
    42842 => -26952,
    42843 => -26953,
    42844 => -26955,
    42845 => -26957,
    42846 => -26959,
    42847 => -26961,
    42848 => -26962,
    42849 => -26964,
    42850 => -26966,
    42851 => -26968,
    42852 => -26969,
    42853 => -26971,
    42854 => -26973,
    42855 => -26975,
    42856 => -26977,
    42857 => -26978,
    42858 => -26980,
    42859 => -26982,
    42860 => -26984,
    42861 => -26986,
    42862 => -26987,
    42863 => -26989,
    42864 => -26991,
    42865 => -26993,
    42866 => -26994,
    42867 => -26996,
    42868 => -26998,
    42869 => -27000,
    42870 => -27002,
    42871 => -27003,
    42872 => -27005,
    42873 => -27007,
    42874 => -27009,
    42875 => -27010,
    42876 => -27012,
    42877 => -27014,
    42878 => -27016,
    42879 => -27018,
    42880 => -27019,
    42881 => -27021,
    42882 => -27023,
    42883 => -27025,
    42884 => -27026,
    42885 => -27028,
    42886 => -27030,
    42887 => -27032,
    42888 => -27034,
    42889 => -27035,
    42890 => -27037,
    42891 => -27039,
    42892 => -27041,
    42893 => -27042,
    42894 => -27044,
    42895 => -27046,
    42896 => -27048,
    42897 => -27049,
    42898 => -27051,
    42899 => -27053,
    42900 => -27055,
    42901 => -27057,
    42902 => -27058,
    42903 => -27060,
    42904 => -27062,
    42905 => -27064,
    42906 => -27065,
    42907 => -27067,
    42908 => -27069,
    42909 => -27071,
    42910 => -27073,
    42911 => -27074,
    42912 => -27076,
    42913 => -27078,
    42914 => -27080,
    42915 => -27081,
    42916 => -27083,
    42917 => -27085,
    42918 => -27087,
    42919 => -27088,
    42920 => -27090,
    42921 => -27092,
    42922 => -27094,
    42923 => -27096,
    42924 => -27097,
    42925 => -27099,
    42926 => -27101,
    42927 => -27103,
    42928 => -27104,
    42929 => -27106,
    42930 => -27108,
    42931 => -27110,
    42932 => -27111,
    42933 => -27113,
    42934 => -27115,
    42935 => -27117,
    42936 => -27118,
    42937 => -27120,
    42938 => -27122,
    42939 => -27124,
    42940 => -27126,
    42941 => -27127,
    42942 => -27129,
    42943 => -27131,
    42944 => -27133,
    42945 => -27134,
    42946 => -27136,
    42947 => -27138,
    42948 => -27140,
    42949 => -27141,
    42950 => -27143,
    42951 => -27145,
    42952 => -27147,
    42953 => -27148,
    42954 => -27150,
    42955 => -27152,
    42956 => -27154,
    42957 => -27155,
    42958 => -27157,
    42959 => -27159,
    42960 => -27161,
    42961 => -27162,
    42962 => -27164,
    42963 => -27166,
    42964 => -27168,
    42965 => -27169,
    42966 => -27171,
    42967 => -27173,
    42968 => -27175,
    42969 => -27177,
    42970 => -27178,
    42971 => -27180,
    42972 => -27182,
    42973 => -27184,
    42974 => -27185,
    42975 => -27187,
    42976 => -27189,
    42977 => -27191,
    42978 => -27192,
    42979 => -27194,
    42980 => -27196,
    42981 => -27198,
    42982 => -27199,
    42983 => -27201,
    42984 => -27203,
    42985 => -27205,
    42986 => -27206,
    42987 => -27208,
    42988 => -27210,
    42989 => -27212,
    42990 => -27213,
    42991 => -27215,
    42992 => -27217,
    42993 => -27219,
    42994 => -27220,
    42995 => -27222,
    42996 => -27224,
    42997 => -27226,
    42998 => -27227,
    42999 => -27229,
    43000 => -27231,
    43001 => -27233,
    43002 => -27234,
    43003 => -27236,
    43004 => -27238,
    43005 => -27240,
    43006 => -27241,
    43007 => -27243,
    43008 => -27245,
    43009 => -27247,
    43010 => -27248,
    43011 => -27250,
    43012 => -27252,
    43013 => -27253,
    43014 => -27255,
    43015 => -27257,
    43016 => -27259,
    43017 => -27260,
    43018 => -27262,
    43019 => -27264,
    43020 => -27266,
    43021 => -27267,
    43022 => -27269,
    43023 => -27271,
    43024 => -27273,
    43025 => -27274,
    43026 => -27276,
    43027 => -27278,
    43028 => -27280,
    43029 => -27281,
    43030 => -27283,
    43031 => -27285,
    43032 => -27287,
    43033 => -27288,
    43034 => -27290,
    43035 => -27292,
    43036 => -27294,
    43037 => -27295,
    43038 => -27297,
    43039 => -27299,
    43040 => -27300,
    43041 => -27302,
    43042 => -27304,
    43043 => -27306,
    43044 => -27307,
    43045 => -27309,
    43046 => -27311,
    43047 => -27313,
    43048 => -27314,
    43049 => -27316,
    43050 => -27318,
    43051 => -27320,
    43052 => -27321,
    43053 => -27323,
    43054 => -27325,
    43055 => -27327,
    43056 => -27328,
    43057 => -27330,
    43058 => -27332,
    43059 => -27333,
    43060 => -27335,
    43061 => -27337,
    43062 => -27339,
    43063 => -27340,
    43064 => -27342,
    43065 => -27344,
    43066 => -27346,
    43067 => -27347,
    43068 => -27349,
    43069 => -27351,
    43070 => -27352,
    43071 => -27354,
    43072 => -27356,
    43073 => -27358,
    43074 => -27359,
    43075 => -27361,
    43076 => -27363,
    43077 => -27365,
    43078 => -27366,
    43079 => -27368,
    43080 => -27370,
    43081 => -27372,
    43082 => -27373,
    43083 => -27375,
    43084 => -27377,
    43085 => -27378,
    43086 => -27380,
    43087 => -27382,
    43088 => -27384,
    43089 => -27385,
    43090 => -27387,
    43091 => -27389,
    43092 => -27390,
    43093 => -27392,
    43094 => -27394,
    43095 => -27396,
    43096 => -27397,
    43097 => -27399,
    43098 => -27401,
    43099 => -27403,
    43100 => -27404,
    43101 => -27406,
    43102 => -27408,
    43103 => -27409,
    43104 => -27411,
    43105 => -27413,
    43106 => -27415,
    43107 => -27416,
    43108 => -27418,
    43109 => -27420,
    43110 => -27421,
    43111 => -27423,
    43112 => -27425,
    43113 => -27427,
    43114 => -27428,
    43115 => -27430,
    43116 => -27432,
    43117 => -27434,
    43118 => -27435,
    43119 => -27437,
    43120 => -27439,
    43121 => -27440,
    43122 => -27442,
    43123 => -27444,
    43124 => -27446,
    43125 => -27447,
    43126 => -27449,
    43127 => -27451,
    43128 => -27452,
    43129 => -27454,
    43130 => -27456,
    43131 => -27458,
    43132 => -27459,
    43133 => -27461,
    43134 => -27463,
    43135 => -27464,
    43136 => -27466,
    43137 => -27468,
    43138 => -27470,
    43139 => -27471,
    43140 => -27473,
    43141 => -27475,
    43142 => -27476,
    43143 => -27478,
    43144 => -27480,
    43145 => -27482,
    43146 => -27483,
    43147 => -27485,
    43148 => -27487,
    43149 => -27488,
    43150 => -27490,
    43151 => -27492,
    43152 => -27493,
    43153 => -27495,
    43154 => -27497,
    43155 => -27499,
    43156 => -27500,
    43157 => -27502,
    43158 => -27504,
    43159 => -27505,
    43160 => -27507,
    43161 => -27509,
    43162 => -27511,
    43163 => -27512,
    43164 => -27514,
    43165 => -27516,
    43166 => -27517,
    43167 => -27519,
    43168 => -27521,
    43169 => -27523,
    43170 => -27524,
    43171 => -27526,
    43172 => -27528,
    43173 => -27529,
    43174 => -27531,
    43175 => -27533,
    43176 => -27534,
    43177 => -27536,
    43178 => -27538,
    43179 => -27540,
    43180 => -27541,
    43181 => -27543,
    43182 => -27545,
    43183 => -27546,
    43184 => -27548,
    43185 => -27550,
    43186 => -27551,
    43187 => -27553,
    43188 => -27555,
    43189 => -27557,
    43190 => -27558,
    43191 => -27560,
    43192 => -27562,
    43193 => -27563,
    43194 => -27565,
    43195 => -27567,
    43196 => -27568,
    43197 => -27570,
    43198 => -27572,
    43199 => -27574,
    43200 => -27575,
    43201 => -27577,
    43202 => -27579,
    43203 => -27580,
    43204 => -27582,
    43205 => -27584,
    43206 => -27585,
    43207 => -27587,
    43208 => -27589,
    43209 => -27590,
    43210 => -27592,
    43211 => -27594,
    43212 => -27596,
    43213 => -27597,
    43214 => -27599,
    43215 => -27601,
    43216 => -27602,
    43217 => -27604,
    43218 => -27606,
    43219 => -27607,
    43220 => -27609,
    43221 => -27611,
    43222 => -27613,
    43223 => -27614,
    43224 => -27616,
    43225 => -27618,
    43226 => -27619,
    43227 => -27621,
    43228 => -27623,
    43229 => -27624,
    43230 => -27626,
    43231 => -27628,
    43232 => -27629,
    43233 => -27631,
    43234 => -27633,
    43235 => -27634,
    43236 => -27636,
    43237 => -27638,
    43238 => -27640,
    43239 => -27641,
    43240 => -27643,
    43241 => -27645,
    43242 => -27646,
    43243 => -27648,
    43244 => -27650,
    43245 => -27651,
    43246 => -27653,
    43247 => -27655,
    43248 => -27656,
    43249 => -27658,
    43250 => -27660,
    43251 => -27661,
    43252 => -27663,
    43253 => -27665,
    43254 => -27666,
    43255 => -27668,
    43256 => -27670,
    43257 => -27672,
    43258 => -27673,
    43259 => -27675,
    43260 => -27677,
    43261 => -27678,
    43262 => -27680,
    43263 => -27682,
    43264 => -27683,
    43265 => -27685,
    43266 => -27687,
    43267 => -27688,
    43268 => -27690,
    43269 => -27692,
    43270 => -27693,
    43271 => -27695,
    43272 => -27697,
    43273 => -27698,
    43274 => -27700,
    43275 => -27702,
    43276 => -27703,
    43277 => -27705,
    43278 => -27707,
    43279 => -27708,
    43280 => -27710,
    43281 => -27712,
    43282 => -27714,
    43283 => -27715,
    43284 => -27717,
    43285 => -27719,
    43286 => -27720,
    43287 => -27722,
    43288 => -27724,
    43289 => -27725,
    43290 => -27727,
    43291 => -27729,
    43292 => -27730,
    43293 => -27732,
    43294 => -27734,
    43295 => -27735,
    43296 => -27737,
    43297 => -27739,
    43298 => -27740,
    43299 => -27742,
    43300 => -27744,
    43301 => -27745,
    43302 => -27747,
    43303 => -27749,
    43304 => -27750,
    43305 => -27752,
    43306 => -27754,
    43307 => -27755,
    43308 => -27757,
    43309 => -27759,
    43310 => -27760,
    43311 => -27762,
    43312 => -27764,
    43313 => -27765,
    43314 => -27767,
    43315 => -27769,
    43316 => -27770,
    43317 => -27772,
    43318 => -27774,
    43319 => -27775,
    43320 => -27777,
    43321 => -27779,
    43322 => -27780,
    43323 => -27782,
    43324 => -27784,
    43325 => -27785,
    43326 => -27787,
    43327 => -27789,
    43328 => -27790,
    43329 => -27792,
    43330 => -27794,
    43331 => -27795,
    43332 => -27797,
    43333 => -27799,
    43334 => -27800,
    43335 => -27802,
    43336 => -27804,
    43337 => -27805,
    43338 => -27807,
    43339 => -27809,
    43340 => -27810,
    43341 => -27812,
    43342 => -27814,
    43343 => -27815,
    43344 => -27817,
    43345 => -27819,
    43346 => -27820,
    43347 => -27822,
    43348 => -27824,
    43349 => -27825,
    43350 => -27827,
    43351 => -27829,
    43352 => -27830,
    43353 => -27832,
    43354 => -27834,
    43355 => -27835,
    43356 => -27837,
    43357 => -27839,
    43358 => -27840,
    43359 => -27842,
    43360 => -27843,
    43361 => -27845,
    43362 => -27847,
    43363 => -27848,
    43364 => -27850,
    43365 => -27852,
    43366 => -27853,
    43367 => -27855,
    43368 => -27857,
    43369 => -27858,
    43370 => -27860,
    43371 => -27862,
    43372 => -27863,
    43373 => -27865,
    43374 => -27867,
    43375 => -27868,
    43376 => -27870,
    43377 => -27872,
    43378 => -27873,
    43379 => -27875,
    43380 => -27877,
    43381 => -27878,
    43382 => -27880,
    43383 => -27882,
    43384 => -27883,
    43385 => -27885,
    43386 => -27886,
    43387 => -27888,
    43388 => -27890,
    43389 => -27891,
    43390 => -27893,
    43391 => -27895,
    43392 => -27896,
    43393 => -27898,
    43394 => -27900,
    43395 => -27901,
    43396 => -27903,
    43397 => -27905,
    43398 => -27906,
    43399 => -27908,
    43400 => -27910,
    43401 => -27911,
    43402 => -27913,
    43403 => -27914,
    43404 => -27916,
    43405 => -27918,
    43406 => -27919,
    43407 => -27921,
    43408 => -27923,
    43409 => -27924,
    43410 => -27926,
    43411 => -27928,
    43412 => -27929,
    43413 => -27931,
    43414 => -27933,
    43415 => -27934,
    43416 => -27936,
    43417 => -27937,
    43418 => -27939,
    43419 => -27941,
    43420 => -27942,
    43421 => -27944,
    43422 => -27946,
    43423 => -27947,
    43424 => -27949,
    43425 => -27951,
    43426 => -27952,
    43427 => -27954,
    43428 => -27956,
    43429 => -27957,
    43430 => -27959,
    43431 => -27960,
    43432 => -27962,
    43433 => -27964,
    43434 => -27965,
    43435 => -27967,
    43436 => -27969,
    43437 => -27970,
    43438 => -27972,
    43439 => -27974,
    43440 => -27975,
    43441 => -27977,
    43442 => -27978,
    43443 => -27980,
    43444 => -27982,
    43445 => -27983,
    43446 => -27985,
    43447 => -27987,
    43448 => -27988,
    43449 => -27990,
    43450 => -27992,
    43451 => -27993,
    43452 => -27995,
    43453 => -27996,
    43454 => -27998,
    43455 => -28000,
    43456 => -28001,
    43457 => -28003,
    43458 => -28005,
    43459 => -28006,
    43460 => -28008,
    43461 => -28009,
    43462 => -28011,
    43463 => -28013,
    43464 => -28014,
    43465 => -28016,
    43466 => -28018,
    43467 => -28019,
    43468 => -28021,
    43469 => -28022,
    43470 => -28024,
    43471 => -28026,
    43472 => -28027,
    43473 => -28029,
    43474 => -28031,
    43475 => -28032,
    43476 => -28034,
    43477 => -28036,
    43478 => -28037,
    43479 => -28039,
    43480 => -28040,
    43481 => -28042,
    43482 => -28044,
    43483 => -28045,
    43484 => -28047,
    43485 => -28049,
    43486 => -28050,
    43487 => -28052,
    43488 => -28053,
    43489 => -28055,
    43490 => -28057,
    43491 => -28058,
    43492 => -28060,
    43493 => -28061,
    43494 => -28063,
    43495 => -28065,
    43496 => -28066,
    43497 => -28068,
    43498 => -28070,
    43499 => -28071,
    43500 => -28073,
    43501 => -28074,
    43502 => -28076,
    43503 => -28078,
    43504 => -28079,
    43505 => -28081,
    43506 => -28083,
    43507 => -28084,
    43508 => -28086,
    43509 => -28087,
    43510 => -28089,
    43511 => -28091,
    43512 => -28092,
    43513 => -28094,
    43514 => -28095,
    43515 => -28097,
    43516 => -28099,
    43517 => -28100,
    43518 => -28102,
    43519 => -28104,
    43520 => -28105,
    43521 => -28107,
    43522 => -28108,
    43523 => -28110,
    43524 => -28112,
    43525 => -28113,
    43526 => -28115,
    43527 => -28116,
    43528 => -28118,
    43529 => -28120,
    43530 => -28121,
    43531 => -28123,
    43532 => -28125,
    43533 => -28126,
    43534 => -28128,
    43535 => -28129,
    43536 => -28131,
    43537 => -28133,
    43538 => -28134,
    43539 => -28136,
    43540 => -28137,
    43541 => -28139,
    43542 => -28141,
    43543 => -28142,
    43544 => -28144,
    43545 => -28145,
    43546 => -28147,
    43547 => -28149,
    43548 => -28150,
    43549 => -28152,
    43550 => -28154,
    43551 => -28155,
    43552 => -28157,
    43553 => -28158,
    43554 => -28160,
    43555 => -28162,
    43556 => -28163,
    43557 => -28165,
    43558 => -28166,
    43559 => -28168,
    43560 => -28170,
    43561 => -28171,
    43562 => -28173,
    43563 => -28174,
    43564 => -28176,
    43565 => -28178,
    43566 => -28179,
    43567 => -28181,
    43568 => -28182,
    43569 => -28184,
    43570 => -28186,
    43571 => -28187,
    43572 => -28189,
    43573 => -28190,
    43574 => -28192,
    43575 => -28194,
    43576 => -28195,
    43577 => -28197,
    43578 => -28198,
    43579 => -28200,
    43580 => -28202,
    43581 => -28203,
    43582 => -28205,
    43583 => -28206,
    43584 => -28208,
    43585 => -28210,
    43586 => -28211,
    43587 => -28213,
    43588 => -28214,
    43589 => -28216,
    43590 => -28218,
    43591 => -28219,
    43592 => -28221,
    43593 => -28222,
    43594 => -28224,
    43595 => -28226,
    43596 => -28227,
    43597 => -28229,
    43598 => -28230,
    43599 => -28232,
    43600 => -28234,
    43601 => -28235,
    43602 => -28237,
    43603 => -28238,
    43604 => -28240,
    43605 => -28242,
    43606 => -28243,
    43607 => -28245,
    43608 => -28246,
    43609 => -28248,
    43610 => -28249,
    43611 => -28251,
    43612 => -28253,
    43613 => -28254,
    43614 => -28256,
    43615 => -28257,
    43616 => -28259,
    43617 => -28261,
    43618 => -28262,
    43619 => -28264,
    43620 => -28265,
    43621 => -28267,
    43622 => -28269,
    43623 => -28270,
    43624 => -28272,
    43625 => -28273,
    43626 => -28275,
    43627 => -28277,
    43628 => -28278,
    43629 => -28280,
    43630 => -28281,
    43631 => -28283,
    43632 => -28284,
    43633 => -28286,
    43634 => -28288,
    43635 => -28289,
    43636 => -28291,
    43637 => -28292,
    43638 => -28294,
    43639 => -28296,
    43640 => -28297,
    43641 => -28299,
    43642 => -28300,
    43643 => -28302,
    43644 => -28303,
    43645 => -28305,
    43646 => -28307,
    43647 => -28308,
    43648 => -28310,
    43649 => -28311,
    43650 => -28313,
    43651 => -28315,
    43652 => -28316,
    43653 => -28318,
    43654 => -28319,
    43655 => -28321,
    43656 => -28322,
    43657 => -28324,
    43658 => -28326,
    43659 => -28327,
    43660 => -28329,
    43661 => -28330,
    43662 => -28332,
    43663 => -28333,
    43664 => -28335,
    43665 => -28337,
    43666 => -28338,
    43667 => -28340,
    43668 => -28341,
    43669 => -28343,
    43670 => -28345,
    43671 => -28346,
    43672 => -28348,
    43673 => -28349,
    43674 => -28351,
    43675 => -28352,
    43676 => -28354,
    43677 => -28356,
    43678 => -28357,
    43679 => -28359,
    43680 => -28360,
    43681 => -28362,
    43682 => -28363,
    43683 => -28365,
    43684 => -28367,
    43685 => -28368,
    43686 => -28370,
    43687 => -28371,
    43688 => -28373,
    43689 => -28374,
    43690 => -28376,
    43691 => -28378,
    43692 => -28379,
    43693 => -28381,
    43694 => -28382,
    43695 => -28384,
    43696 => -28385,
    43697 => -28387,
    43698 => -28389,
    43699 => -28390,
    43700 => -28392,
    43701 => -28393,
    43702 => -28395,
    43703 => -28396,
    43704 => -28398,
    43705 => -28400,
    43706 => -28401,
    43707 => -28403,
    43708 => -28404,
    43709 => -28406,
    43710 => -28407,
    43711 => -28409,
    43712 => -28411,
    43713 => -28412,
    43714 => -28414,
    43715 => -28415,
    43716 => -28417,
    43717 => -28418,
    43718 => -28420,
    43719 => -28421,
    43720 => -28423,
    43721 => -28425,
    43722 => -28426,
    43723 => -28428,
    43724 => -28429,
    43725 => -28431,
    43726 => -28432,
    43727 => -28434,
    43728 => -28436,
    43729 => -28437,
    43730 => -28439,
    43731 => -28440,
    43732 => -28442,
    43733 => -28443,
    43734 => -28445,
    43735 => -28446,
    43736 => -28448,
    43737 => -28450,
    43738 => -28451,
    43739 => -28453,
    43740 => -28454,
    43741 => -28456,
    43742 => -28457,
    43743 => -28459,
    43744 => -28460,
    43745 => -28462,
    43746 => -28464,
    43747 => -28465,
    43748 => -28467,
    43749 => -28468,
    43750 => -28470,
    43751 => -28471,
    43752 => -28473,
    43753 => -28474,
    43754 => -28476,
    43755 => -28478,
    43756 => -28479,
    43757 => -28481,
    43758 => -28482,
    43759 => -28484,
    43760 => -28485,
    43761 => -28487,
    43762 => -28488,
    43763 => -28490,
    43764 => -28492,
    43765 => -28493,
    43766 => -28495,
    43767 => -28496,
    43768 => -28498,
    43769 => -28499,
    43770 => -28501,
    43771 => -28502,
    43772 => -28504,
    43773 => -28505,
    43774 => -28507,
    43775 => -28509,
    43776 => -28510,
    43777 => -28512,
    43778 => -28513,
    43779 => -28515,
    43780 => -28516,
    43781 => -28518,
    43782 => -28519,
    43783 => -28521,
    43784 => -28523,
    43785 => -28524,
    43786 => -28526,
    43787 => -28527,
    43788 => -28529,
    43789 => -28530,
    43790 => -28532,
    43791 => -28533,
    43792 => -28535,
    43793 => -28536,
    43794 => -28538,
    43795 => -28540,
    43796 => -28541,
    43797 => -28543,
    43798 => -28544,
    43799 => -28546,
    43800 => -28547,
    43801 => -28549,
    43802 => -28550,
    43803 => -28552,
    43804 => -28553,
    43805 => -28555,
    43806 => -28556,
    43807 => -28558,
    43808 => -28560,
    43809 => -28561,
    43810 => -28563,
    43811 => -28564,
    43812 => -28566,
    43813 => -28567,
    43814 => -28569,
    43815 => -28570,
    43816 => -28572,
    43817 => -28573,
    43818 => -28575,
    43819 => -28576,
    43820 => -28578,
    43821 => -28580,
    43822 => -28581,
    43823 => -28583,
    43824 => -28584,
    43825 => -28586,
    43826 => -28587,
    43827 => -28589,
    43828 => -28590,
    43829 => -28592,
    43830 => -28593,
    43831 => -28595,
    43832 => -28596,
    43833 => -28598,
    43834 => -28600,
    43835 => -28601,
    43836 => -28603,
    43837 => -28604,
    43838 => -28606,
    43839 => -28607,
    43840 => -28609,
    43841 => -28610,
    43842 => -28612,
    43843 => -28613,
    43844 => -28615,
    43845 => -28616,
    43846 => -28618,
    43847 => -28619,
    43848 => -28621,
    43849 => -28622,
    43850 => -28624,
    43851 => -28626,
    43852 => -28627,
    43853 => -28629,
    43854 => -28630,
    43855 => -28632,
    43856 => -28633,
    43857 => -28635,
    43858 => -28636,
    43859 => -28638,
    43860 => -28639,
    43861 => -28641,
    43862 => -28642,
    43863 => -28644,
    43864 => -28645,
    43865 => -28647,
    43866 => -28648,
    43867 => -28650,
    43868 => -28651,
    43869 => -28653,
    43870 => -28655,
    43871 => -28656,
    43872 => -28658,
    43873 => -28659,
    43874 => -28661,
    43875 => -28662,
    43876 => -28664,
    43877 => -28665,
    43878 => -28667,
    43879 => -28668,
    43880 => -28670,
    43881 => -28671,
    43882 => -28673,
    43883 => -28674,
    43884 => -28676,
    43885 => -28677,
    43886 => -28679,
    43887 => -28680,
    43888 => -28682,
    43889 => -28683,
    43890 => -28685,
    43891 => -28686,
    43892 => -28688,
    43893 => -28690,
    43894 => -28691,
    43895 => -28693,
    43896 => -28694,
    43897 => -28696,
    43898 => -28697,
    43899 => -28699,
    43900 => -28700,
    43901 => -28702,
    43902 => -28703,
    43903 => -28705,
    43904 => -28706,
    43905 => -28708,
    43906 => -28709,
    43907 => -28711,
    43908 => -28712,
    43909 => -28714,
    43910 => -28715,
    43911 => -28717,
    43912 => -28718,
    43913 => -28720,
    43914 => -28721,
    43915 => -28723,
    43916 => -28724,
    43917 => -28726,
    43918 => -28727,
    43919 => -28729,
    43920 => -28730,
    43921 => -28732,
    43922 => -28733,
    43923 => -28735,
    43924 => -28736,
    43925 => -28738,
    43926 => -28739,
    43927 => -28741,
    43928 => -28742,
    43929 => -28744,
    43930 => -28745,
    43931 => -28747,
    43932 => -28748,
    43933 => -28750,
    43934 => -28752,
    43935 => -28753,
    43936 => -28755,
    43937 => -28756,
    43938 => -28758,
    43939 => -28759,
    43940 => -28761,
    43941 => -28762,
    43942 => -28764,
    43943 => -28765,
    43944 => -28767,
    43945 => -28768,
    43946 => -28770,
    43947 => -28771,
    43948 => -28773,
    43949 => -28774,
    43950 => -28776,
    43951 => -28777,
    43952 => -28779,
    43953 => -28780,
    43954 => -28782,
    43955 => -28783,
    43956 => -28785,
    43957 => -28786,
    43958 => -28788,
    43959 => -28789,
    43960 => -28791,
    43961 => -28792,
    43962 => -28794,
    43963 => -28795,
    43964 => -28797,
    43965 => -28798,
    43966 => -28800,
    43967 => -28801,
    43968 => -28803,
    43969 => -28804,
    43970 => -28806,
    43971 => -28807,
    43972 => -28809,
    43973 => -28810,
    43974 => -28812,
    43975 => -28813,
    43976 => -28815,
    43977 => -28816,
    43978 => -28818,
    43979 => -28819,
    43980 => -28821,
    43981 => -28822,
    43982 => -28824,
    43983 => -28825,
    43984 => -28827,
    43985 => -28828,
    43986 => -28830,
    43987 => -28831,
    43988 => -28832,
    43989 => -28834,
    43990 => -28835,
    43991 => -28837,
    43992 => -28838,
    43993 => -28840,
    43994 => -28841,
    43995 => -28843,
    43996 => -28844,
    43997 => -28846,
    43998 => -28847,
    43999 => -28849,
    44000 => -28850,
    44001 => -28852,
    44002 => -28853,
    44003 => -28855,
    44004 => -28856,
    44005 => -28858,
    44006 => -28859,
    44007 => -28861,
    44008 => -28862,
    44009 => -28864,
    44010 => -28865,
    44011 => -28867,
    44012 => -28868,
    44013 => -28870,
    44014 => -28871,
    44015 => -28873,
    44016 => -28874,
    44017 => -28876,
    44018 => -28877,
    44019 => -28879,
    44020 => -28880,
    44021 => -28882,
    44022 => -28883,
    44023 => -28885,
    44024 => -28886,
    44025 => -28888,
    44026 => -28889,
    44027 => -28891,
    44028 => -28892,
    44029 => -28893,
    44030 => -28895,
    44031 => -28896,
    44032 => -28898,
    44033 => -28899,
    44034 => -28901,
    44035 => -28902,
    44036 => -28904,
    44037 => -28905,
    44038 => -28907,
    44039 => -28908,
    44040 => -28910,
    44041 => -28911,
    44042 => -28913,
    44043 => -28914,
    44044 => -28916,
    44045 => -28917,
    44046 => -28919,
    44047 => -28920,
    44048 => -28922,
    44049 => -28923,
    44050 => -28925,
    44051 => -28926,
    44052 => -28927,
    44053 => -28929,
    44054 => -28930,
    44055 => -28932,
    44056 => -28933,
    44057 => -28935,
    44058 => -28936,
    44059 => -28938,
    44060 => -28939,
    44061 => -28941,
    44062 => -28942,
    44063 => -28944,
    44064 => -28945,
    44065 => -28947,
    44066 => -28948,
    44067 => -28950,
    44068 => -28951,
    44069 => -28953,
    44070 => -28954,
    44071 => -28955,
    44072 => -28957,
    44073 => -28958,
    44074 => -28960,
    44075 => -28961,
    44076 => -28963,
    44077 => -28964,
    44078 => -28966,
    44079 => -28967,
    44080 => -28969,
    44081 => -28970,
    44082 => -28972,
    44083 => -28973,
    44084 => -28975,
    44085 => -28976,
    44086 => -28977,
    44087 => -28979,
    44088 => -28980,
    44089 => -28982,
    44090 => -28983,
    44091 => -28985,
    44092 => -28986,
    44093 => -28988,
    44094 => -28989,
    44095 => -28991,
    44096 => -28992,
    44097 => -28994,
    44098 => -28995,
    44099 => -28997,
    44100 => -28998,
    44101 => -28999,
    44102 => -29001,
    44103 => -29002,
    44104 => -29004,
    44105 => -29005,
    44106 => -29007,
    44107 => -29008,
    44108 => -29010,
    44109 => -29011,
    44110 => -29013,
    44111 => -29014,
    44112 => -29016,
    44113 => -29017,
    44114 => -29018,
    44115 => -29020,
    44116 => -29021,
    44117 => -29023,
    44118 => -29024,
    44119 => -29026,
    44120 => -29027,
    44121 => -29029,
    44122 => -29030,
    44123 => -29032,
    44124 => -29033,
    44125 => -29034,
    44126 => -29036,
    44127 => -29037,
    44128 => -29039,
    44129 => -29040,
    44130 => -29042,
    44131 => -29043,
    44132 => -29045,
    44133 => -29046,
    44134 => -29048,
    44135 => -29049,
    44136 => -29050,
    44137 => -29052,
    44138 => -29053,
    44139 => -29055,
    44140 => -29056,
    44141 => -29058,
    44142 => -29059,
    44143 => -29061,
    44144 => -29062,
    44145 => -29064,
    44146 => -29065,
    44147 => -29066,
    44148 => -29068,
    44149 => -29069,
    44150 => -29071,
    44151 => -29072,
    44152 => -29074,
    44153 => -29075,
    44154 => -29077,
    44155 => -29078,
    44156 => -29079,
    44157 => -29081,
    44158 => -29082,
    44159 => -29084,
    44160 => -29085,
    44161 => -29087,
    44162 => -29088,
    44163 => -29090,
    44164 => -29091,
    44165 => -29093,
    44166 => -29094,
    44167 => -29095,
    44168 => -29097,
    44169 => -29098,
    44170 => -29100,
    44171 => -29101,
    44172 => -29103,
    44173 => -29104,
    44174 => -29106,
    44175 => -29107,
    44176 => -29108,
    44177 => -29110,
    44178 => -29111,
    44179 => -29113,
    44180 => -29114,
    44181 => -29116,
    44182 => -29117,
    44183 => -29118,
    44184 => -29120,
    44185 => -29121,
    44186 => -29123,
    44187 => -29124,
    44188 => -29126,
    44189 => -29127,
    44190 => -29129,
    44191 => -29130,
    44192 => -29131,
    44193 => -29133,
    44194 => -29134,
    44195 => -29136,
    44196 => -29137,
    44197 => -29139,
    44198 => -29140,
    44199 => -29142,
    44200 => -29143,
    44201 => -29144,
    44202 => -29146,
    44203 => -29147,
    44204 => -29149,
    44205 => -29150,
    44206 => -29152,
    44207 => -29153,
    44208 => -29154,
    44209 => -29156,
    44210 => -29157,
    44211 => -29159,
    44212 => -29160,
    44213 => -29162,
    44214 => -29163,
    44215 => -29164,
    44216 => -29166,
    44217 => -29167,
    44218 => -29169,
    44219 => -29170,
    44220 => -29172,
    44221 => -29173,
    44222 => -29174,
    44223 => -29176,
    44224 => -29177,
    44225 => -29179,
    44226 => -29180,
    44227 => -29182,
    44228 => -29183,
    44229 => -29184,
    44230 => -29186,
    44231 => -29187,
    44232 => -29189,
    44233 => -29190,
    44234 => -29192,
    44235 => -29193,
    44236 => -29194,
    44237 => -29196,
    44238 => -29197,
    44239 => -29199,
    44240 => -29200,
    44241 => -29202,
    44242 => -29203,
    44243 => -29204,
    44244 => -29206,
    44245 => -29207,
    44246 => -29209,
    44247 => -29210,
    44248 => -29212,
    44249 => -29213,
    44250 => -29214,
    44251 => -29216,
    44252 => -29217,
    44253 => -29219,
    44254 => -29220,
    44255 => -29222,
    44256 => -29223,
    44257 => -29224,
    44258 => -29226,
    44259 => -29227,
    44260 => -29229,
    44261 => -29230,
    44262 => -29231,
    44263 => -29233,
    44264 => -29234,
    44265 => -29236,
    44266 => -29237,
    44267 => -29239,
    44268 => -29240,
    44269 => -29241,
    44270 => -29243,
    44271 => -29244,
    44272 => -29246,
    44273 => -29247,
    44274 => -29248,
    44275 => -29250,
    44276 => -29251,
    44277 => -29253,
    44278 => -29254,
    44279 => -29256,
    44280 => -29257,
    44281 => -29258,
    44282 => -29260,
    44283 => -29261,
    44284 => -29263,
    44285 => -29264,
    44286 => -29265,
    44287 => -29267,
    44288 => -29268,
    44289 => -29270,
    44290 => -29271,
    44291 => -29273,
    44292 => -29274,
    44293 => -29275,
    44294 => -29277,
    44295 => -29278,
    44296 => -29280,
    44297 => -29281,
    44298 => -29282,
    44299 => -29284,
    44300 => -29285,
    44301 => -29287,
    44302 => -29288,
    44303 => -29289,
    44304 => -29291,
    44305 => -29292,
    44306 => -29294,
    44307 => -29295,
    44308 => -29296,
    44309 => -29298,
    44310 => -29299,
    44311 => -29301,
    44312 => -29302,
    44313 => -29304,
    44314 => -29305,
    44315 => -29306,
    44316 => -29308,
    44317 => -29309,
    44318 => -29311,
    44319 => -29312,
    44320 => -29313,
    44321 => -29315,
    44322 => -29316,
    44323 => -29318,
    44324 => -29319,
    44325 => -29320,
    44326 => -29322,
    44327 => -29323,
    44328 => -29325,
    44329 => -29326,
    44330 => -29327,
    44331 => -29329,
    44332 => -29330,
    44333 => -29332,
    44334 => -29333,
    44335 => -29334,
    44336 => -29336,
    44337 => -29337,
    44338 => -29339,
    44339 => -29340,
    44340 => -29341,
    44341 => -29343,
    44342 => -29344,
    44343 => -29346,
    44344 => -29347,
    44345 => -29348,
    44346 => -29350,
    44347 => -29351,
    44348 => -29353,
    44349 => -29354,
    44350 => -29355,
    44351 => -29357,
    44352 => -29358,
    44353 => -29360,
    44354 => -29361,
    44355 => -29362,
    44356 => -29364,
    44357 => -29365,
    44358 => -29366,
    44359 => -29368,
    44360 => -29369,
    44361 => -29371,
    44362 => -29372,
    44363 => -29373,
    44364 => -29375,
    44365 => -29376,
    44366 => -29378,
    44367 => -29379,
    44368 => -29380,
    44369 => -29382,
    44370 => -29383,
    44371 => -29385,
    44372 => -29386,
    44373 => -29387,
    44374 => -29389,
    44375 => -29390,
    44376 => -29392,
    44377 => -29393,
    44378 => -29394,
    44379 => -29396,
    44380 => -29397,
    44381 => -29398,
    44382 => -29400,
    44383 => -29401,
    44384 => -29403,
    44385 => -29404,
    44386 => -29405,
    44387 => -29407,
    44388 => -29408,
    44389 => -29410,
    44390 => -29411,
    44391 => -29412,
    44392 => -29414,
    44393 => -29415,
    44394 => -29416,
    44395 => -29418,
    44396 => -29419,
    44397 => -29421,
    44398 => -29422,
    44399 => -29423,
    44400 => -29425,
    44401 => -29426,
    44402 => -29428,
    44403 => -29429,
    44404 => -29430,
    44405 => -29432,
    44406 => -29433,
    44407 => -29434,
    44408 => -29436,
    44409 => -29437,
    44410 => -29439,
    44411 => -29440,
    44412 => -29441,
    44413 => -29443,
    44414 => -29444,
    44415 => -29445,
    44416 => -29447,
    44417 => -29448,
    44418 => -29450,
    44419 => -29451,
    44420 => -29452,
    44421 => -29454,
    44422 => -29455,
    44423 => -29457,
    44424 => -29458,
    44425 => -29459,
    44426 => -29461,
    44427 => -29462,
    44428 => -29463,
    44429 => -29465,
    44430 => -29466,
    44431 => -29468,
    44432 => -29469,
    44433 => -29470,
    44434 => -29472,
    44435 => -29473,
    44436 => -29474,
    44437 => -29476,
    44438 => -29477,
    44439 => -29478,
    44440 => -29480,
    44441 => -29481,
    44442 => -29483,
    44443 => -29484,
    44444 => -29485,
    44445 => -29487,
    44446 => -29488,
    44447 => -29489,
    44448 => -29491,
    44449 => -29492,
    44450 => -29494,
    44451 => -29495,
    44452 => -29496,
    44453 => -29498,
    44454 => -29499,
    44455 => -29500,
    44456 => -29502,
    44457 => -29503,
    44458 => -29504,
    44459 => -29506,
    44460 => -29507,
    44461 => -29509,
    44462 => -29510,
    44463 => -29511,
    44464 => -29513,
    44465 => -29514,
    44466 => -29515,
    44467 => -29517,
    44468 => -29518,
    44469 => -29520,
    44470 => -29521,
    44471 => -29522,
    44472 => -29524,
    44473 => -29525,
    44474 => -29526,
    44475 => -29528,
    44476 => -29529,
    44477 => -29530,
    44478 => -29532,
    44479 => -29533,
    44480 => -29534,
    44481 => -29536,
    44482 => -29537,
    44483 => -29539,
    44484 => -29540,
    44485 => -29541,
    44486 => -29543,
    44487 => -29544,
    44488 => -29545,
    44489 => -29547,
    44490 => -29548,
    44491 => -29549,
    44492 => -29551,
    44493 => -29552,
    44494 => -29554,
    44495 => -29555,
    44496 => -29556,
    44497 => -29558,
    44498 => -29559,
    44499 => -29560,
    44500 => -29562,
    44501 => -29563,
    44502 => -29564,
    44503 => -29566,
    44504 => -29567,
    44505 => -29568,
    44506 => -29570,
    44507 => -29571,
    44508 => -29572,
    44509 => -29574,
    44510 => -29575,
    44511 => -29577,
    44512 => -29578,
    44513 => -29579,
    44514 => -29581,
    44515 => -29582,
    44516 => -29583,
    44517 => -29585,
    44518 => -29586,
    44519 => -29587,
    44520 => -29589,
    44521 => -29590,
    44522 => -29591,
    44523 => -29593,
    44524 => -29594,
    44525 => -29595,
    44526 => -29597,
    44527 => -29598,
    44528 => -29599,
    44529 => -29601,
    44530 => -29602,
    44531 => -29604,
    44532 => -29605,
    44533 => -29606,
    44534 => -29608,
    44535 => -29609,
    44536 => -29610,
    44537 => -29612,
    44538 => -29613,
    44539 => -29614,
    44540 => -29616,
    44541 => -29617,
    44542 => -29618,
    44543 => -29620,
    44544 => -29621,
    44545 => -29622,
    44546 => -29624,
    44547 => -29625,
    44548 => -29626,
    44549 => -29628,
    44550 => -29629,
    44551 => -29630,
    44552 => -29632,
    44553 => -29633,
    44554 => -29634,
    44555 => -29636,
    44556 => -29637,
    44557 => -29638,
    44558 => -29640,
    44559 => -29641,
    44560 => -29642,
    44561 => -29644,
    44562 => -29645,
    44563 => -29646,
    44564 => -29648,
    44565 => -29649,
    44566 => -29651,
    44567 => -29652,
    44568 => -29653,
    44569 => -29655,
    44570 => -29656,
    44571 => -29657,
    44572 => -29659,
    44573 => -29660,
    44574 => -29661,
    44575 => -29663,
    44576 => -29664,
    44577 => -29665,
    44578 => -29667,
    44579 => -29668,
    44580 => -29669,
    44581 => -29671,
    44582 => -29672,
    44583 => -29673,
    44584 => -29675,
    44585 => -29676,
    44586 => -29677,
    44587 => -29679,
    44588 => -29680,
    44589 => -29681,
    44590 => -29683,
    44591 => -29684,
    44592 => -29685,
    44593 => -29687,
    44594 => -29688,
    44595 => -29689,
    44596 => -29690,
    44597 => -29692,
    44598 => -29693,
    44599 => -29694,
    44600 => -29696,
    44601 => -29697,
    44602 => -29698,
    44603 => -29700,
    44604 => -29701,
    44605 => -29702,
    44606 => -29704,
    44607 => -29705,
    44608 => -29706,
    44609 => -29708,
    44610 => -29709,
    44611 => -29710,
    44612 => -29712,
    44613 => -29713,
    44614 => -29714,
    44615 => -29716,
    44616 => -29717,
    44617 => -29718,
    44618 => -29720,
    44619 => -29721,
    44620 => -29722,
    44621 => -29724,
    44622 => -29725,
    44623 => -29726,
    44624 => -29728,
    44625 => -29729,
    44626 => -29730,
    44627 => -29732,
    44628 => -29733,
    44629 => -29734,
    44630 => -29736,
    44631 => -29737,
    44632 => -29738,
    44633 => -29739,
    44634 => -29741,
    44635 => -29742,
    44636 => -29743,
    44637 => -29745,
    44638 => -29746,
    44639 => -29747,
    44640 => -29749,
    44641 => -29750,
    44642 => -29751,
    44643 => -29753,
    44644 => -29754,
    44645 => -29755,
    44646 => -29757,
    44647 => -29758,
    44648 => -29759,
    44649 => -29761,
    44650 => -29762,
    44651 => -29763,
    44652 => -29764,
    44653 => -29766,
    44654 => -29767,
    44655 => -29768,
    44656 => -29770,
    44657 => -29771,
    44658 => -29772,
    44659 => -29774,
    44660 => -29775,
    44661 => -29776,
    44662 => -29778,
    44663 => -29779,
    44664 => -29780,
    44665 => -29782,
    44666 => -29783,
    44667 => -29784,
    44668 => -29785,
    44669 => -29787,
    44670 => -29788,
    44671 => -29789,
    44672 => -29791,
    44673 => -29792,
    44674 => -29793,
    44675 => -29795,
    44676 => -29796,
    44677 => -29797,
    44678 => -29799,
    44679 => -29800,
    44680 => -29801,
    44681 => -29802,
    44682 => -29804,
    44683 => -29805,
    44684 => -29806,
    44685 => -29808,
    44686 => -29809,
    44687 => -29810,
    44688 => -29812,
    44689 => -29813,
    44690 => -29814,
    44691 => -29816,
    44692 => -29817,
    44693 => -29818,
    44694 => -29819,
    44695 => -29821,
    44696 => -29822,
    44697 => -29823,
    44698 => -29825,
    44699 => -29826,
    44700 => -29827,
    44701 => -29829,
    44702 => -29830,
    44703 => -29831,
    44704 => -29832,
    44705 => -29834,
    44706 => -29835,
    44707 => -29836,
    44708 => -29838,
    44709 => -29839,
    44710 => -29840,
    44711 => -29842,
    44712 => -29843,
    44713 => -29844,
    44714 => -29845,
    44715 => -29847,
    44716 => -29848,
    44717 => -29849,
    44718 => -29851,
    44719 => -29852,
    44720 => -29853,
    44721 => -29854,
    44722 => -29856,
    44723 => -29857,
    44724 => -29858,
    44725 => -29860,
    44726 => -29861,
    44727 => -29862,
    44728 => -29864,
    44729 => -29865,
    44730 => -29866,
    44731 => -29867,
    44732 => -29869,
    44733 => -29870,
    44734 => -29871,
    44735 => -29873,
    44736 => -29874,
    44737 => -29875,
    44738 => -29876,
    44739 => -29878,
    44740 => -29879,
    44741 => -29880,
    44742 => -29882,
    44743 => -29883,
    44744 => -29884,
    44745 => -29885,
    44746 => -29887,
    44747 => -29888,
    44748 => -29889,
    44749 => -29891,
    44750 => -29892,
    44751 => -29893,
    44752 => -29894,
    44753 => -29896,
    44754 => -29897,
    44755 => -29898,
    44756 => -29900,
    44757 => -29901,
    44758 => -29902,
    44759 => -29903,
    44760 => -29905,
    44761 => -29906,
    44762 => -29907,
    44763 => -29909,
    44764 => -29910,
    44765 => -29911,
    44766 => -29912,
    44767 => -29914,
    44768 => -29915,
    44769 => -29916,
    44770 => -29918,
    44771 => -29919,
    44772 => -29920,
    44773 => -29921,
    44774 => -29923,
    44775 => -29924,
    44776 => -29925,
    44777 => -29927,
    44778 => -29928,
    44779 => -29929,
    44780 => -29930,
    44781 => -29932,
    44782 => -29933,
    44783 => -29934,
    44784 => -29936,
    44785 => -29937,
    44786 => -29938,
    44787 => -29939,
    44788 => -29941,
    44789 => -29942,
    44790 => -29943,
    44791 => -29944,
    44792 => -29946,
    44793 => -29947,
    44794 => -29948,
    44795 => -29950,
    44796 => -29951,
    44797 => -29952,
    44798 => -29953,
    44799 => -29955,
    44800 => -29956,
    44801 => -29957,
    44802 => -29958,
    44803 => -29960,
    44804 => -29961,
    44805 => -29962,
    44806 => -29964,
    44807 => -29965,
    44808 => -29966,
    44809 => -29967,
    44810 => -29969,
    44811 => -29970,
    44812 => -29971,
    44813 => -29972,
    44814 => -29974,
    44815 => -29975,
    44816 => -29976,
    44817 => -29978,
    44818 => -29979,
    44819 => -29980,
    44820 => -29981,
    44821 => -29983,
    44822 => -29984,
    44823 => -29985,
    44824 => -29986,
    44825 => -29988,
    44826 => -29989,
    44827 => -29990,
    44828 => -29991,
    44829 => -29993,
    44830 => -29994,
    44831 => -29995,
    44832 => -29997,
    44833 => -29998,
    44834 => -29999,
    44835 => -30000,
    44836 => -30002,
    44837 => -30003,
    44838 => -30004,
    44839 => -30005,
    44840 => -30007,
    44841 => -30008,
    44842 => -30009,
    44843 => -30010,
    44844 => -30012,
    44845 => -30013,
    44846 => -30014,
    44847 => -30015,
    44848 => -30017,
    44849 => -30018,
    44850 => -30019,
    44851 => -30020,
    44852 => -30022,
    44853 => -30023,
    44854 => -30024,
    44855 => -30026,
    44856 => -30027,
    44857 => -30028,
    44858 => -30029,
    44859 => -30031,
    44860 => -30032,
    44861 => -30033,
    44862 => -30034,
    44863 => -30036,
    44864 => -30037,
    44865 => -30038,
    44866 => -30039,
    44867 => -30041,
    44868 => -30042,
    44869 => -30043,
    44870 => -30044,
    44871 => -30046,
    44872 => -30047,
    44873 => -30048,
    44874 => -30049,
    44875 => -30051,
    44876 => -30052,
    44877 => -30053,
    44878 => -30054,
    44879 => -30056,
    44880 => -30057,
    44881 => -30058,
    44882 => -30059,
    44883 => -30061,
    44884 => -30062,
    44885 => -30063,
    44886 => -30064,
    44887 => -30066,
    44888 => -30067,
    44889 => -30068,
    44890 => -30069,
    44891 => -30071,
    44892 => -30072,
    44893 => -30073,
    44894 => -30074,
    44895 => -30076,
    44896 => -30077,
    44897 => -30078,
    44898 => -30079,
    44899 => -30081,
    44900 => -30082,
    44901 => -30083,
    44902 => -30084,
    44903 => -30086,
    44904 => -30087,
    44905 => -30088,
    44906 => -30089,
    44907 => -30091,
    44908 => -30092,
    44909 => -30093,
    44910 => -30094,
    44911 => -30096,
    44912 => -30097,
    44913 => -30098,
    44914 => -30099,
    44915 => -30100,
    44916 => -30102,
    44917 => -30103,
    44918 => -30104,
    44919 => -30105,
    44920 => -30107,
    44921 => -30108,
    44922 => -30109,
    44923 => -30110,
    44924 => -30112,
    44925 => -30113,
    44926 => -30114,
    44927 => -30115,
    44928 => -30117,
    44929 => -30118,
    44930 => -30119,
    44931 => -30120,
    44932 => -30122,
    44933 => -30123,
    44934 => -30124,
    44935 => -30125,
    44936 => -30126,
    44937 => -30128,
    44938 => -30129,
    44939 => -30130,
    44940 => -30131,
    44941 => -30133,
    44942 => -30134,
    44943 => -30135,
    44944 => -30136,
    44945 => -30138,
    44946 => -30139,
    44947 => -30140,
    44948 => -30141,
    44949 => -30143,
    44950 => -30144,
    44951 => -30145,
    44952 => -30146,
    44953 => -30147,
    44954 => -30149,
    44955 => -30150,
    44956 => -30151,
    44957 => -30152,
    44958 => -30154,
    44959 => -30155,
    44960 => -30156,
    44961 => -30157,
    44962 => -30159,
    44963 => -30160,
    44964 => -30161,
    44965 => -30162,
    44966 => -30163,
    44967 => -30165,
    44968 => -30166,
    44969 => -30167,
    44970 => -30168,
    44971 => -30170,
    44972 => -30171,
    44973 => -30172,
    44974 => -30173,
    44975 => -30174,
    44976 => -30176,
    44977 => -30177,
    44978 => -30178,
    44979 => -30179,
    44980 => -30181,
    44981 => -30182,
    44982 => -30183,
    44983 => -30184,
    44984 => -30185,
    44985 => -30187,
    44986 => -30188,
    44987 => -30189,
    44988 => -30190,
    44989 => -30192,
    44990 => -30193,
    44991 => -30194,
    44992 => -30195,
    44993 => -30196,
    44994 => -30198,
    44995 => -30199,
    44996 => -30200,
    44997 => -30201,
    44998 => -30203,
    44999 => -30204,
    45000 => -30205,
    45001 => -30206,
    45002 => -30207,
    45003 => -30209,
    45004 => -30210,
    45005 => -30211,
    45006 => -30212,
    45007 => -30214,
    45008 => -30215,
    45009 => -30216,
    45010 => -30217,
    45011 => -30218,
    45012 => -30220,
    45013 => -30221,
    45014 => -30222,
    45015 => -30223,
    45016 => -30224,
    45017 => -30226,
    45018 => -30227,
    45019 => -30228,
    45020 => -30229,
    45021 => -30231,
    45022 => -30232,
    45023 => -30233,
    45024 => -30234,
    45025 => -30235,
    45026 => -30237,
    45027 => -30238,
    45028 => -30239,
    45029 => -30240,
    45030 => -30241,
    45031 => -30243,
    45032 => -30244,
    45033 => -30245,
    45034 => -30246,
    45035 => -30247,
    45036 => -30249,
    45037 => -30250,
    45038 => -30251,
    45039 => -30252,
    45040 => -30253,
    45041 => -30255,
    45042 => -30256,
    45043 => -30257,
    45044 => -30258,
    45045 => -30260,
    45046 => -30261,
    45047 => -30262,
    45048 => -30263,
    45049 => -30264,
    45050 => -30266,
    45051 => -30267,
    45052 => -30268,
    45053 => -30269,
    45054 => -30270,
    45055 => -30272,
    45056 => -30273,
    45057 => -30274,
    45058 => -30275,
    45059 => -30276,
    45060 => -30278,
    45061 => -30279,
    45062 => -30280,
    45063 => -30281,
    45064 => -30282,
    45065 => -30284,
    45066 => -30285,
    45067 => -30286,
    45068 => -30287,
    45069 => -30288,
    45070 => -30290,
    45071 => -30291,
    45072 => -30292,
    45073 => -30293,
    45074 => -30294,
    45075 => -30296,
    45076 => -30297,
    45077 => -30298,
    45078 => -30299,
    45079 => -30300,
    45080 => -30302,
    45081 => -30303,
    45082 => -30304,
    45083 => -30305,
    45084 => -30306,
    45085 => -30308,
    45086 => -30309,
    45087 => -30310,
    45088 => -30311,
    45089 => -30312,
    45090 => -30313,
    45091 => -30315,
    45092 => -30316,
    45093 => -30317,
    45094 => -30318,
    45095 => -30319,
    45096 => -30321,
    45097 => -30322,
    45098 => -30323,
    45099 => -30324,
    45100 => -30325,
    45101 => -30327,
    45102 => -30328,
    45103 => -30329,
    45104 => -30330,
    45105 => -30331,
    45106 => -30333,
    45107 => -30334,
    45108 => -30335,
    45109 => -30336,
    45110 => -30337,
    45111 => -30338,
    45112 => -30340,
    45113 => -30341,
    45114 => -30342,
    45115 => -30343,
    45116 => -30344,
    45117 => -30346,
    45118 => -30347,
    45119 => -30348,
    45120 => -30349,
    45121 => -30350,
    45122 => -30351,
    45123 => -30353,
    45124 => -30354,
    45125 => -30355,
    45126 => -30356,
    45127 => -30357,
    45128 => -30359,
    45129 => -30360,
    45130 => -30361,
    45131 => -30362,
    45132 => -30363,
    45133 => -30365,
    45134 => -30366,
    45135 => -30367,
    45136 => -30368,
    45137 => -30369,
    45138 => -30370,
    45139 => -30372,
    45140 => -30373,
    45141 => -30374,
    45142 => -30375,
    45143 => -30376,
    45144 => -30377,
    45145 => -30379,
    45146 => -30380,
    45147 => -30381,
    45148 => -30382,
    45149 => -30383,
    45150 => -30385,
    45151 => -30386,
    45152 => -30387,
    45153 => -30388,
    45154 => -30389,
    45155 => -30390,
    45156 => -30392,
    45157 => -30393,
    45158 => -30394,
    45159 => -30395,
    45160 => -30396,
    45161 => -30397,
    45162 => -30399,
    45163 => -30400,
    45164 => -30401,
    45165 => -30402,
    45166 => -30403,
    45167 => -30404,
    45168 => -30406,
    45169 => -30407,
    45170 => -30408,
    45171 => -30409,
    45172 => -30410,
    45173 => -30412,
    45174 => -30413,
    45175 => -30414,
    45176 => -30415,
    45177 => -30416,
    45178 => -30417,
    45179 => -30419,
    45180 => -30420,
    45181 => -30421,
    45182 => -30422,
    45183 => -30423,
    45184 => -30424,
    45185 => -30426,
    45186 => -30427,
    45187 => -30428,
    45188 => -30429,
    45189 => -30430,
    45190 => -30431,
    45191 => -30433,
    45192 => -30434,
    45193 => -30435,
    45194 => -30436,
    45195 => -30437,
    45196 => -30438,
    45197 => -30439,
    45198 => -30441,
    45199 => -30442,
    45200 => -30443,
    45201 => -30444,
    45202 => -30445,
    45203 => -30446,
    45204 => -30448,
    45205 => -30449,
    45206 => -30450,
    45207 => -30451,
    45208 => -30452,
    45209 => -30453,
    45210 => -30455,
    45211 => -30456,
    45212 => -30457,
    45213 => -30458,
    45214 => -30459,
    45215 => -30460,
    45216 => -30462,
    45217 => -30463,
    45218 => -30464,
    45219 => -30465,
    45220 => -30466,
    45221 => -30467,
    45222 => -30468,
    45223 => -30470,
    45224 => -30471,
    45225 => -30472,
    45226 => -30473,
    45227 => -30474,
    45228 => -30475,
    45229 => -30477,
    45230 => -30478,
    45231 => -30479,
    45232 => -30480,
    45233 => -30481,
    45234 => -30482,
    45235 => -30483,
    45236 => -30485,
    45237 => -30486,
    45238 => -30487,
    45239 => -30488,
    45240 => -30489,
    45241 => -30490,
    45242 => -30492,
    45243 => -30493,
    45244 => -30494,
    45245 => -30495,
    45246 => -30496,
    45247 => -30497,
    45248 => -30498,
    45249 => -30500,
    45250 => -30501,
    45251 => -30502,
    45252 => -30503,
    45253 => -30504,
    45254 => -30505,
    45255 => -30506,
    45256 => -30508,
    45257 => -30509,
    45258 => -30510,
    45259 => -30511,
    45260 => -30512,
    45261 => -30513,
    45262 => -30514,
    45263 => -30516,
    45264 => -30517,
    45265 => -30518,
    45266 => -30519,
    45267 => -30520,
    45268 => -30521,
    45269 => -30522,
    45270 => -30524,
    45271 => -30525,
    45272 => -30526,
    45273 => -30527,
    45274 => -30528,
    45275 => -30529,
    45276 => -30530,
    45277 => -30532,
    45278 => -30533,
    45279 => -30534,
    45280 => -30535,
    45281 => -30536,
    45282 => -30537,
    45283 => -30538,
    45284 => -30540,
    45285 => -30541,
    45286 => -30542,
    45287 => -30543,
    45288 => -30544,
    45289 => -30545,
    45290 => -30546,
    45291 => -30548,
    45292 => -30549,
    45293 => -30550,
    45294 => -30551,
    45295 => -30552,
    45296 => -30553,
    45297 => -30554,
    45298 => -30556,
    45299 => -30557,
    45300 => -30558,
    45301 => -30559,
    45302 => -30560,
    45303 => -30561,
    45304 => -30562,
    45305 => -30563,
    45306 => -30565,
    45307 => -30566,
    45308 => -30567,
    45309 => -30568,
    45310 => -30569,
    45311 => -30570,
    45312 => -30571,
    45313 => -30573,
    45314 => -30574,
    45315 => -30575,
    45316 => -30576,
    45317 => -30577,
    45318 => -30578,
    45319 => -30579,
    45320 => -30580,
    45321 => -30582,
    45322 => -30583,
    45323 => -30584,
    45324 => -30585,
    45325 => -30586,
    45326 => -30587,
    45327 => -30588,
    45328 => -30589,
    45329 => -30591,
    45330 => -30592,
    45331 => -30593,
    45332 => -30594,
    45333 => -30595,
    45334 => -30596,
    45335 => -30597,
    45336 => -30598,
    45337 => -30600,
    45338 => -30601,
    45339 => -30602,
    45340 => -30603,
    45341 => -30604,
    45342 => -30605,
    45343 => -30606,
    45344 => -30607,
    45345 => -30609,
    45346 => -30610,
    45347 => -30611,
    45348 => -30612,
    45349 => -30613,
    45350 => -30614,
    45351 => -30615,
    45352 => -30616,
    45353 => -30617,
    45354 => -30619,
    45355 => -30620,
    45356 => -30621,
    45357 => -30622,
    45358 => -30623,
    45359 => -30624,
    45360 => -30625,
    45361 => -30626,
    45362 => -30628,
    45363 => -30629,
    45364 => -30630,
    45365 => -30631,
    45366 => -30632,
    45367 => -30633,
    45368 => -30634,
    45369 => -30635,
    45370 => -30636,
    45371 => -30638,
    45372 => -30639,
    45373 => -30640,
    45374 => -30641,
    45375 => -30642,
    45376 => -30643,
    45377 => -30644,
    45378 => -30645,
    45379 => -30646,
    45380 => -30648,
    45381 => -30649,
    45382 => -30650,
    45383 => -30651,
    45384 => -30652,
    45385 => -30653,
    45386 => -30654,
    45387 => -30655,
    45388 => -30656,
    45389 => -30658,
    45390 => -30659,
    45391 => -30660,
    45392 => -30661,
    45393 => -30662,
    45394 => -30663,
    45395 => -30664,
    45396 => -30665,
    45397 => -30666,
    45398 => -30668,
    45399 => -30669,
    45400 => -30670,
    45401 => -30671,
    45402 => -30672,
    45403 => -30673,
    45404 => -30674,
    45405 => -30675,
    45406 => -30676,
    45407 => -30678,
    45408 => -30679,
    45409 => -30680,
    45410 => -30681,
    45411 => -30682,
    45412 => -30683,
    45413 => -30684,
    45414 => -30685,
    45415 => -30686,
    45416 => -30687,
    45417 => -30689,
    45418 => -30690,
    45419 => -30691,
    45420 => -30692,
    45421 => -30693,
    45422 => -30694,
    45423 => -30695,
    45424 => -30696,
    45425 => -30697,
    45426 => -30698,
    45427 => -30700,
    45428 => -30701,
    45429 => -30702,
    45430 => -30703,
    45431 => -30704,
    45432 => -30705,
    45433 => -30706,
    45434 => -30707,
    45435 => -30708,
    45436 => -30709,
    45437 => -30711,
    45438 => -30712,
    45439 => -30713,
    45440 => -30714,
    45441 => -30715,
    45442 => -30716,
    45443 => -30717,
    45444 => -30718,
    45445 => -30719,
    45446 => -30720,
    45447 => -30721,
    45448 => -30723,
    45449 => -30724,
    45450 => -30725,
    45451 => -30726,
    45452 => -30727,
    45453 => -30728,
    45454 => -30729,
    45455 => -30730,
    45456 => -30731,
    45457 => -30732,
    45458 => -30733,
    45459 => -30735,
    45460 => -30736,
    45461 => -30737,
    45462 => -30738,
    45463 => -30739,
    45464 => -30740,
    45465 => -30741,
    45466 => -30742,
    45467 => -30743,
    45468 => -30744,
    45469 => -30745,
    45470 => -30746,
    45471 => -30748,
    45472 => -30749,
    45473 => -30750,
    45474 => -30751,
    45475 => -30752,
    45476 => -30753,
    45477 => -30754,
    45478 => -30755,
    45479 => -30756,
    45480 => -30757,
    45481 => -30758,
    45482 => -30760,
    45483 => -30761,
    45484 => -30762,
    45485 => -30763,
    45486 => -30764,
    45487 => -30765,
    45488 => -30766,
    45489 => -30767,
    45490 => -30768,
    45491 => -30769,
    45492 => -30770,
    45493 => -30771,
    45494 => -30772,
    45495 => -30774,
    45496 => -30775,
    45497 => -30776,
    45498 => -30777,
    45499 => -30778,
    45500 => -30779,
    45501 => -30780,
    45502 => -30781,
    45503 => -30782,
    45504 => -30783,
    45505 => -30784,
    45506 => -30785,
    45507 => -30786,
    45508 => -30788,
    45509 => -30789,
    45510 => -30790,
    45511 => -30791,
    45512 => -30792,
    45513 => -30793,
    45514 => -30794,
    45515 => -30795,
    45516 => -30796,
    45517 => -30797,
    45518 => -30798,
    45519 => -30799,
    45520 => -30800,
    45521 => -30802,
    45522 => -30803,
    45523 => -30804,
    45524 => -30805,
    45525 => -30806,
    45526 => -30807,
    45527 => -30808,
    45528 => -30809,
    45529 => -30810,
    45530 => -30811,
    45531 => -30812,
    45532 => -30813,
    45533 => -30814,
    45534 => -30815,
    45535 => -30816,
    45536 => -30818,
    45537 => -30819,
    45538 => -30820,
    45539 => -30821,
    45540 => -30822,
    45541 => -30823,
    45542 => -30824,
    45543 => -30825,
    45544 => -30826,
    45545 => -30827,
    45546 => -30828,
    45547 => -30829,
    45548 => -30830,
    45549 => -30831,
    45550 => -30832,
    45551 => -30834,
    45552 => -30835,
    45553 => -30836,
    45554 => -30837,
    45555 => -30838,
    45556 => -30839,
    45557 => -30840,
    45558 => -30841,
    45559 => -30842,
    45560 => -30843,
    45561 => -30844,
    45562 => -30845,
    45563 => -30846,
    45564 => -30847,
    45565 => -30848,
    45566 => -30849,
    45567 => -30851,
    45568 => -30852,
    45569 => -30853,
    45570 => -30854,
    45571 => -30855,
    45572 => -30856,
    45573 => -30857,
    45574 => -30858,
    45575 => -30859,
    45576 => -30860,
    45577 => -30861,
    45578 => -30862,
    45579 => -30863,
    45580 => -30864,
    45581 => -30865,
    45582 => -30866,
    45583 => -30867,
    45584 => -30868,
    45585 => -30870,
    45586 => -30871,
    45587 => -30872,
    45588 => -30873,
    45589 => -30874,
    45590 => -30875,
    45591 => -30876,
    45592 => -30877,
    45593 => -30878,
    45594 => -30879,
    45595 => -30880,
    45596 => -30881,
    45597 => -30882,
    45598 => -30883,
    45599 => -30884,
    45600 => -30885,
    45601 => -30886,
    45602 => -30887,
    45603 => -30888,
    45604 => -30889,
    45605 => -30891,
    45606 => -30892,
    45607 => -30893,
    45608 => -30894,
    45609 => -30895,
    45610 => -30896,
    45611 => -30897,
    45612 => -30898,
    45613 => -30899,
    45614 => -30900,
    45615 => -30901,
    45616 => -30902,
    45617 => -30903,
    45618 => -30904,
    45619 => -30905,
    45620 => -30906,
    45621 => -30907,
    45622 => -30908,
    45623 => -30909,
    45624 => -30910,
    45625 => -30911,
    45626 => -30912,
    45627 => -30914,
    45628 => -30915,
    45629 => -30916,
    45630 => -30917,
    45631 => -30918,
    45632 => -30919,
    45633 => -30920,
    45634 => -30921,
    45635 => -30922,
    45636 => -30923,
    45637 => -30924,
    45638 => -30925,
    45639 => -30926,
    45640 => -30927,
    45641 => -30928,
    45642 => -30929,
    45643 => -30930,
    45644 => -30931,
    45645 => -30932,
    45646 => -30933,
    45647 => -30934,
    45648 => -30935,
    45649 => -30936,
    45650 => -30937,
    45651 => -30938,
    45652 => -30939,
    45653 => -30941,
    45654 => -30942,
    45655 => -30943,
    45656 => -30944,
    45657 => -30945,
    45658 => -30946,
    45659 => -30947,
    45660 => -30948,
    45661 => -30949,
    45662 => -30950,
    45663 => -30951,
    45664 => -30952,
    45665 => -30953,
    45666 => -30954,
    45667 => -30955,
    45668 => -30956,
    45669 => -30957,
    45670 => -30958,
    45671 => -30959,
    45672 => -30960,
    45673 => -30961,
    45674 => -30962,
    45675 => -30963,
    45676 => -30964,
    45677 => -30965,
    45678 => -30966,
    45679 => -30967,
    45680 => -30968,
    45681 => -30969,
    45682 => -30970,
    45683 => -30971,
    45684 => -30972,
    45685 => -30973,
    45686 => -30974,
    45687 => -30976,
    45688 => -30977,
    45689 => -30978,
    45690 => -30979,
    45691 => -30980,
    45692 => -30981,
    45693 => -30982,
    45694 => -30983,
    45695 => -30984,
    45696 => -30985,
    45697 => -30986,
    45698 => -30987,
    45699 => -30988,
    45700 => -30989,
    45701 => -30990,
    45702 => -30991,
    45703 => -30992,
    45704 => -30993,
    45705 => -30994,
    45706 => -30995,
    45707 => -30996,
    45708 => -30997,
    45709 => -30998,
    45710 => -30999,
    45711 => -31000,
    45712 => -31001,
    45713 => -31002,
    45714 => -31003,
    45715 => -31004,
    45716 => -31005,
    45717 => -31006,
    45718 => -31007,
    45719 => -31008,
    45720 => -31009,
    45721 => -31010,
    45722 => -31011,
    45723 => -31012,
    45724 => -31013,
    45725 => -31014,
    45726 => -31015,
    45727 => -31016,
    45728 => -31017,
    45729 => -31018,
    45730 => -31019,
    45731 => -31020,
    45732 => -31021,
    45733 => -31022,
    45734 => -31023,
    45735 => -31024,
    45736 => -31025,
    45737 => -31026,
    45738 => -31027,
    45739 => -31028,
    45740 => -31029,
    45741 => -31030,
    45742 => -31031,
    45743 => -31032,
    45744 => -31033,
    45745 => -31034,
    45746 => -31035,
    45747 => -31036,
    45748 => -31037,
    45749 => -31038,
    45750 => -31039,
    45751 => -31040,
    45752 => -31041,
    45753 => -31043,
    45754 => -31044,
    45755 => -31045,
    45756 => -31046,
    45757 => -31047,
    45758 => -31048,
    45759 => -31049,
    45760 => -31050,
    45761 => -31051,
    45762 => -31052,
    45763 => -31053,
    45764 => -31054,
    45765 => -31055,
    45766 => -31056,
    45767 => -31057,
    45768 => -31058,
    45769 => -31059,
    45770 => -31060,
    45771 => -31061,
    45772 => -31062,
    45773 => -31063,
    45774 => -31064,
    45775 => -31065,
    45776 => -31066,
    45777 => -31067,
    45778 => -31068,
    45779 => -31069,
    45780 => -31070,
    45781 => -31071,
    45782 => -31072,
    45783 => -31073,
    45784 => -31074,
    45785 => -31075,
    45786 => -31076,
    45787 => -31077,
    45788 => -31078,
    45789 => -31079,
    45790 => -31080,
    45791 => -31081,
    45792 => -31082,
    45793 => -31083,
    45794 => -31083,
    45795 => -31084,
    45796 => -31085,
    45797 => -31086,
    45798 => -31087,
    45799 => -31088,
    45800 => -31089,
    45801 => -31090,
    45802 => -31091,
    45803 => -31092,
    45804 => -31093,
    45805 => -31094,
    45806 => -31095,
    45807 => -31096,
    45808 => -31097,
    45809 => -31098,
    45810 => -31099,
    45811 => -31100,
    45812 => -31101,
    45813 => -31102,
    45814 => -31103,
    45815 => -31104,
    45816 => -31105,
    45817 => -31106,
    45818 => -31107,
    45819 => -31108,
    45820 => -31109,
    45821 => -31110,
    45822 => -31111,
    45823 => -31112,
    45824 => -31113,
    45825 => -31114,
    45826 => -31115,
    45827 => -31116,
    45828 => -31117,
    45829 => -31118,
    45830 => -31119,
    45831 => -31120,
    45832 => -31121,
    45833 => -31122,
    45834 => -31123,
    45835 => -31124,
    45836 => -31125,
    45837 => -31126,
    45838 => -31127,
    45839 => -31128,
    45840 => -31129,
    45841 => -31130,
    45842 => -31131,
    45843 => -31132,
    45844 => -31133,
    45845 => -31134,
    45846 => -31135,
    45847 => -31136,
    45848 => -31137,
    45849 => -31138,
    45850 => -31139,
    45851 => -31140,
    45852 => -31141,
    45853 => -31142,
    45854 => -31143,
    45855 => -31144,
    45856 => -31145,
    45857 => -31146,
    45858 => -31147,
    45859 => -31148,
    45860 => -31148,
    45861 => -31149,
    45862 => -31150,
    45863 => -31151,
    45864 => -31152,
    45865 => -31153,
    45866 => -31154,
    45867 => -31155,
    45868 => -31156,
    45869 => -31157,
    45870 => -31158,
    45871 => -31159,
    45872 => -31160,
    45873 => -31161,
    45874 => -31162,
    45875 => -31163,
    45876 => -31164,
    45877 => -31165,
    45878 => -31166,
    45879 => -31167,
    45880 => -31168,
    45881 => -31169,
    45882 => -31170,
    45883 => -31171,
    45884 => -31172,
    45885 => -31173,
    45886 => -31174,
    45887 => -31175,
    45888 => -31176,
    45889 => -31177,
    45890 => -31178,
    45891 => -31179,
    45892 => -31180,
    45893 => -31181,
    45894 => -31181,
    45895 => -31182,
    45896 => -31183,
    45897 => -31184,
    45898 => -31185,
    45899 => -31186,
    45900 => -31187,
    45901 => -31188,
    45902 => -31189,
    45903 => -31190,
    45904 => -31191,
    45905 => -31192,
    45906 => -31193,
    45907 => -31194,
    45908 => -31195,
    45909 => -31196,
    45910 => -31197,
    45911 => -31198,
    45912 => -31199,
    45913 => -31200,
    45914 => -31201,
    45915 => -31202,
    45916 => -31203,
    45917 => -31204,
    45918 => -31205,
    45919 => -31206,
    45920 => -31206,
    45921 => -31207,
    45922 => -31208,
    45923 => -31209,
    45924 => -31210,
    45925 => -31211,
    45926 => -31212,
    45927 => -31213,
    45928 => -31214,
    45929 => -31215,
    45930 => -31216,
    45931 => -31217,
    45932 => -31218,
    45933 => -31219,
    45934 => -31220,
    45935 => -31221,
    45936 => -31222,
    45937 => -31223,
    45938 => -31224,
    45939 => -31225,
    45940 => -31226,
    45941 => -31227,
    45942 => -31227,
    45943 => -31228,
    45944 => -31229,
    45945 => -31230,
    45946 => -31231,
    45947 => -31232,
    45948 => -31233,
    45949 => -31234,
    45950 => -31235,
    45951 => -31236,
    45952 => -31237,
    45953 => -31238,
    45954 => -31239,
    45955 => -31240,
    45956 => -31241,
    45957 => -31242,
    45958 => -31243,
    45959 => -31244,
    45960 => -31245,
    45961 => -31246,
    45962 => -31246,
    45963 => -31247,
    45964 => -31248,
    45965 => -31249,
    45966 => -31250,
    45967 => -31251,
    45968 => -31252,
    45969 => -31253,
    45970 => -31254,
    45971 => -31255,
    45972 => -31256,
    45973 => -31257,
    45974 => -31258,
    45975 => -31259,
    45976 => -31260,
    45977 => -31261,
    45978 => -31262,
    45979 => -31262,
    45980 => -31263,
    45981 => -31264,
    45982 => -31265,
    45983 => -31266,
    45984 => -31267,
    45985 => -31268,
    45986 => -31269,
    45987 => -31270,
    45988 => -31271,
    45989 => -31272,
    45990 => -31273,
    45991 => -31274,
    45992 => -31275,
    45993 => -31276,
    45994 => -31277,
    45995 => -31278,
    45996 => -31278,
    45997 => -31279,
    45998 => -31280,
    45999 => -31281,
    46000 => -31282,
    46001 => -31283,
    46002 => -31284,
    46003 => -31285,
    46004 => -31286,
    46005 => -31287,
    46006 => -31288,
    46007 => -31289,
    46008 => -31290,
    46009 => -31291,
    46010 => -31292,
    46011 => -31292,
    46012 => -31293,
    46013 => -31294,
    46014 => -31295,
    46015 => -31296,
    46016 => -31297,
    46017 => -31298,
    46018 => -31299,
    46019 => -31300,
    46020 => -31301,
    46021 => -31302,
    46022 => -31303,
    46023 => -31304,
    46024 => -31305,
    46025 => -31305,
    46026 => -31306,
    46027 => -31307,
    46028 => -31308,
    46029 => -31309,
    46030 => -31310,
    46031 => -31311,
    46032 => -31312,
    46033 => -31313,
    46034 => -31314,
    46035 => -31315,
    46036 => -31316,
    46037 => -31317,
    46038 => -31318,
    46039 => -31318,
    46040 => -31319,
    46041 => -31320,
    46042 => -31321,
    46043 => -31322,
    46044 => -31323,
    46045 => -31324,
    46046 => -31325,
    46047 => -31326,
    46048 => -31327,
    46049 => -31328,
    46050 => -31329,
    46051 => -31329,
    46052 => -31330,
    46053 => -31331,
    46054 => -31332,
    46055 => -31333,
    46056 => -31334,
    46057 => -31335,
    46058 => -31336,
    46059 => -31337,
    46060 => -31338,
    46061 => -31339,
    46062 => -31340,
    46063 => -31341,
    46064 => -31341,
    46065 => -31342,
    46066 => -31343,
    46067 => -31344,
    46068 => -31345,
    46069 => -31346,
    46070 => -31347,
    46071 => -31348,
    46072 => -31349,
    46073 => -31350,
    46074 => -31351,
    46075 => -31352,
    46076 => -31352,
    46077 => -31353,
    46078 => -31354,
    46079 => -31355,
    46080 => -31356,
    46081 => -31357,
    46082 => -31358,
    46083 => -31359,
    46084 => -31360,
    46085 => -31361,
    46086 => -31362,
    46087 => -31362,
    46088 => -31363,
    46089 => -31364,
    46090 => -31365,
    46091 => -31366,
    46092 => -31367,
    46093 => -31368,
    46094 => -31369,
    46095 => -31370,
    46096 => -31371,
    46097 => -31372,
    46098 => -31372,
    46099 => -31373,
    46100 => -31374,
    46101 => -31375,
    46102 => -31376,
    46103 => -31377,
    46104 => -31378,
    46105 => -31379,
    46106 => -31380,
    46107 => -31381,
    46108 => -31381,
    46109 => -31382,
    46110 => -31383,
    46111 => -31384,
    46112 => -31385,
    46113 => -31386,
    46114 => -31387,
    46115 => -31388,
    46116 => -31389,
    46117 => -31390,
    46118 => -31391,
    46119 => -31391,
    46120 => -31392,
    46121 => -31393,
    46122 => -31394,
    46123 => -31395,
    46124 => -31396,
    46125 => -31397,
    46126 => -31398,
    46127 => -31399,
    46128 => -31400,
    46129 => -31400,
    46130 => -31401,
    46131 => -31402,
    46132 => -31403,
    46133 => -31404,
    46134 => -31405,
    46135 => -31406,
    46136 => -31407,
    46137 => -31408,
    46138 => -31408,
    46139 => -31409,
    46140 => -31410,
    46141 => -31411,
    46142 => -31412,
    46143 => -31413,
    46144 => -31414,
    46145 => -31415,
    46146 => -31416,
    46147 => -31417,
    46148 => -31417,
    46149 => -31418,
    46150 => -31419,
    46151 => -31420,
    46152 => -31421,
    46153 => -31422,
    46154 => -31423,
    46155 => -31424,
    46156 => -31425,
    46157 => -31425,
    46158 => -31426,
    46159 => -31427,
    46160 => -31428,
    46161 => -31429,
    46162 => -31430,
    46163 => -31431,
    46164 => -31432,
    46165 => -31433,
    46166 => -31433,
    46167 => -31434,
    46168 => -31435,
    46169 => -31436,
    46170 => -31437,
    46171 => -31438,
    46172 => -31439,
    46173 => -31440,
    46174 => -31441,
    46175 => -31441,
    46176 => -31442,
    46177 => -31443,
    46178 => -31444,
    46179 => -31445,
    46180 => -31446,
    46181 => -31447,
    46182 => -31448,
    46183 => -31448,
    46184 => -31449,
    46185 => -31450,
    46186 => -31451,
    46187 => -31452,
    46188 => -31453,
    46189 => -31454,
    46190 => -31455,
    46191 => -31456,
    46192 => -31456,
    46193 => -31457,
    46194 => -31458,
    46195 => -31459,
    46196 => -31460,
    46197 => -31461,
    46198 => -31462,
    46199 => -31463,
    46200 => -31463,
    46201 => -31464,
    46202 => -31465,
    46203 => -31466,
    46204 => -31467,
    46205 => -31468,
    46206 => -31469,
    46207 => -31470,
    46208 => -31470,
    46209 => -31471,
    46210 => -31472,
    46211 => -31473,
    46212 => -31474,
    46213 => -31475,
    46214 => -31476,
    46215 => -31477,
    46216 => -31477,
    46217 => -31478,
    46218 => -31479,
    46219 => -31480,
    46220 => -31481,
    46221 => -31482,
    46222 => -31483,
    46223 => -31484,
    46224 => -31484,
    46225 => -31485,
    46226 => -31486,
    46227 => -31487,
    46228 => -31488,
    46229 => -31489,
    46230 => -31490,
    46231 => -31490,
    46232 => -31491,
    46233 => -31492,
    46234 => -31493,
    46235 => -31494,
    46236 => -31495,
    46237 => -31496,
    46238 => -31497,
    46239 => -31497,
    46240 => -31498,
    46241 => -31499,
    46242 => -31500,
    46243 => -31501,
    46244 => -31502,
    46245 => -31503,
    46246 => -31503,
    46247 => -31504,
    46248 => -31505,
    46249 => -31506,
    46250 => -31507,
    46251 => -31508,
    46252 => -31509,
    46253 => -31510,
    46254 => -31510,
    46255 => -31511,
    46256 => -31512,
    46257 => -31513,
    46258 => -31514,
    46259 => -31515,
    46260 => -31516,
    46261 => -31516,
    46262 => -31517,
    46263 => -31518,
    46264 => -31519,
    46265 => -31520,
    46266 => -31521,
    46267 => -31522,
    46268 => -31522,
    46269 => -31523,
    46270 => -31524,
    46271 => -31525,
    46272 => -31526,
    46273 => -31527,
    46274 => -31528,
    46275 => -31528,
    46276 => -31529,
    46277 => -31530,
    46278 => -31531,
    46279 => -31532,
    46280 => -31533,
    46281 => -31534,
    46282 => -31534,
    46283 => -31535,
    46284 => -31536,
    46285 => -31537,
    46286 => -31538,
    46287 => -31539,
    46288 => -31539,
    46289 => -31540,
    46290 => -31541,
    46291 => -31542,
    46292 => -31543,
    46293 => -31544,
    46294 => -31545,
    46295 => -31545,
    46296 => -31546,
    46297 => -31547,
    46298 => -31548,
    46299 => -31549,
    46300 => -31550,
    46301 => -31551,
    46302 => -31551,
    46303 => -31552,
    46304 => -31553,
    46305 => -31554,
    46306 => -31555,
    46307 => -31556,
    46308 => -31556,
    46309 => -31557,
    46310 => -31558,
    46311 => -31559,
    46312 => -31560,
    46313 => -31561,
    46314 => -31562,
    46315 => -31562,
    46316 => -31563,
    46317 => -31564,
    46318 => -31565,
    46319 => -31566,
    46320 => -31567,
    46321 => -31567,
    46322 => -31568,
    46323 => -31569,
    46324 => -31570,
    46325 => -31571,
    46326 => -31572,
    46327 => -31572,
    46328 => -31573,
    46329 => -31574,
    46330 => -31575,
    46331 => -31576,
    46332 => -31577,
    46333 => -31578,
    46334 => -31578,
    46335 => -31579,
    46336 => -31580,
    46337 => -31581,
    46338 => -31582,
    46339 => -31583,
    46340 => -31583,
    46341 => -31584,
    46342 => -31585,
    46343 => -31586,
    46344 => -31587,
    46345 => -31588,
    46346 => -31588,
    46347 => -31589,
    46348 => -31590,
    46349 => -31591,
    46350 => -31592,
    46351 => -31593,
    46352 => -31593,
    46353 => -31594,
    46354 => -31595,
    46355 => -31596,
    46356 => -31597,
    46357 => -31598,
    46358 => -31598,
    46359 => -31599,
    46360 => -31600,
    46361 => -31601,
    46362 => -31602,
    46363 => -31603,
    46364 => -31603,
    46365 => -31604,
    46366 => -31605,
    46367 => -31606,
    46368 => -31607,
    46369 => -31608,
    46370 => -31608,
    46371 => -31609,
    46372 => -31610,
    46373 => -31611,
    46374 => -31612,
    46375 => -31613,
    46376 => -31613,
    46377 => -31614,
    46378 => -31615,
    46379 => -31616,
    46380 => -31617,
    46381 => -31617,
    46382 => -31618,
    46383 => -31619,
    46384 => -31620,
    46385 => -31621,
    46386 => -31622,
    46387 => -31622,
    46388 => -31623,
    46389 => -31624,
    46390 => -31625,
    46391 => -31626,
    46392 => -31627,
    46393 => -31627,
    46394 => -31628,
    46395 => -31629,
    46396 => -31630,
    46397 => -31631,
    46398 => -31631,
    46399 => -31632,
    46400 => -31633,
    46401 => -31634,
    46402 => -31635,
    46403 => -31636,
    46404 => -31636,
    46405 => -31637,
    46406 => -31638,
    46407 => -31639,
    46408 => -31640,
    46409 => -31640,
    46410 => -31641,
    46411 => -31642,
    46412 => -31643,
    46413 => -31644,
    46414 => -31645,
    46415 => -31645,
    46416 => -31646,
    46417 => -31647,
    46418 => -31648,
    46419 => -31649,
    46420 => -31649,
    46421 => -31650,
    46422 => -31651,
    46423 => -31652,
    46424 => -31653,
    46425 => -31653,
    46426 => -31654,
    46427 => -31655,
    46428 => -31656,
    46429 => -31657,
    46430 => -31658,
    46431 => -31658,
    46432 => -31659,
    46433 => -31660,
    46434 => -31661,
    46435 => -31662,
    46436 => -31662,
    46437 => -31663,
    46438 => -31664,
    46439 => -31665,
    46440 => -31666,
    46441 => -31666,
    46442 => -31667,
    46443 => -31668,
    46444 => -31669,
    46445 => -31670,
    46446 => -31670,
    46447 => -31671,
    46448 => -31672,
    46449 => -31673,
    46450 => -31674,
    46451 => -31674,
    46452 => -31675,
    46453 => -31676,
    46454 => -31677,
    46455 => -31678,
    46456 => -31679,
    46457 => -31679,
    46458 => -31680,
    46459 => -31681,
    46460 => -31682,
    46461 => -31683,
    46462 => -31683,
    46463 => -31684,
    46464 => -31685,
    46465 => -31686,
    46466 => -31687,
    46467 => -31687,
    46468 => -31688,
    46469 => -31689,
    46470 => -31690,
    46471 => -31691,
    46472 => -31691,
    46473 => -31692,
    46474 => -31693,
    46475 => -31694,
    46476 => -31695,
    46477 => -31695,
    46478 => -31696,
    46479 => -31697,
    46480 => -31698,
    46481 => -31698,
    46482 => -31699,
    46483 => -31700,
    46484 => -31701,
    46485 => -31702,
    46486 => -31702,
    46487 => -31703,
    46488 => -31704,
    46489 => -31705,
    46490 => -31706,
    46491 => -31706,
    46492 => -31707,
    46493 => -31708,
    46494 => -31709,
    46495 => -31710,
    46496 => -31710,
    46497 => -31711,
    46498 => -31712,
    46499 => -31713,
    46500 => -31714,
    46501 => -31714,
    46502 => -31715,
    46503 => -31716,
    46504 => -31717,
    46505 => -31718,
    46506 => -31718,
    46507 => -31719,
    46508 => -31720,
    46509 => -31721,
    46510 => -31721,
    46511 => -31722,
    46512 => -31723,
    46513 => -31724,
    46514 => -31725,
    46515 => -31725,
    46516 => -31726,
    46517 => -31727,
    46518 => -31728,
    46519 => -31729,
    46520 => -31729,
    46521 => -31730,
    46522 => -31731,
    46523 => -31732,
    46524 => -31732,
    46525 => -31733,
    46526 => -31734,
    46527 => -31735,
    46528 => -31736,
    46529 => -31736,
    46530 => -31737,
    46531 => -31738,
    46532 => -31739,
    46533 => -31739,
    46534 => -31740,
    46535 => -31741,
    46536 => -31742,
    46537 => -31743,
    46538 => -31743,
    46539 => -31744,
    46540 => -31745,
    46541 => -31746,
    46542 => -31746,
    46543 => -31747,
    46544 => -31748,
    46545 => -31749,
    46546 => -31750,
    46547 => -31750,
    46548 => -31751,
    46549 => -31752,
    46550 => -31753,
    46551 => -31753,
    46552 => -31754,
    46553 => -31755,
    46554 => -31756,
    46555 => -31757,
    46556 => -31757,
    46557 => -31758,
    46558 => -31759,
    46559 => -31760,
    46560 => -31760,
    46561 => -31761,
    46562 => -31762,
    46563 => -31763,
    46564 => -31764,
    46565 => -31764,
    46566 => -31765,
    46567 => -31766,
    46568 => -31767,
    46569 => -31767,
    46570 => -31768,
    46571 => -31769,
    46572 => -31770,
    46573 => -31770,
    46574 => -31771,
    46575 => -31772,
    46576 => -31773,
    46577 => -31774,
    46578 => -31774,
    46579 => -31775,
    46580 => -31776,
    46581 => -31777,
    46582 => -31777,
    46583 => -31778,
    46584 => -31779,
    46585 => -31780,
    46586 => -31780,
    46587 => -31781,
    46588 => -31782,
    46589 => -31783,
    46590 => -31783,
    46591 => -31784,
    46592 => -31785,
    46593 => -31786,
    46594 => -31787,
    46595 => -31787,
    46596 => -31788,
    46597 => -31789,
    46598 => -31790,
    46599 => -31790,
    46600 => -31791,
    46601 => -31792,
    46602 => -31793,
    46603 => -31793,
    46604 => -31794,
    46605 => -31795,
    46606 => -31796,
    46607 => -31796,
    46608 => -31797,
    46609 => -31798,
    46610 => -31799,
    46611 => -31799,
    46612 => -31800,
    46613 => -31801,
    46614 => -31802,
    46615 => -31802,
    46616 => -31803,
    46617 => -31804,
    46618 => -31805,
    46619 => -31806,
    46620 => -31806,
    46621 => -31807,
    46622 => -31808,
    46623 => -31809,
    46624 => -31809,
    46625 => -31810,
    46626 => -31811,
    46627 => -31812,
    46628 => -31812,
    46629 => -31813,
    46630 => -31814,
    46631 => -31815,
    46632 => -31815,
    46633 => -31816,
    46634 => -31817,
    46635 => -31818,
    46636 => -31818,
    46637 => -31819,
    46638 => -31820,
    46639 => -31821,
    46640 => -31821,
    46641 => -31822,
    46642 => -31823,
    46643 => -31824,
    46644 => -31824,
    46645 => -31825,
    46646 => -31826,
    46647 => -31827,
    46648 => -31827,
    46649 => -31828,
    46650 => -31829,
    46651 => -31830,
    46652 => -31830,
    46653 => -31831,
    46654 => -31832,
    46655 => -31833,
    46656 => -31833,
    46657 => -31834,
    46658 => -31835,
    46659 => -31836,
    46660 => -31836,
    46661 => -31837,
    46662 => -31838,
    46663 => -31838,
    46664 => -31839,
    46665 => -31840,
    46666 => -31841,
    46667 => -31841,
    46668 => -31842,
    46669 => -31843,
    46670 => -31844,
    46671 => -31844,
    46672 => -31845,
    46673 => -31846,
    46674 => -31847,
    46675 => -31847,
    46676 => -31848,
    46677 => -31849,
    46678 => -31850,
    46679 => -31850,
    46680 => -31851,
    46681 => -31852,
    46682 => -31853,
    46683 => -31853,
    46684 => -31854,
    46685 => -31855,
    46686 => -31855,
    46687 => -31856,
    46688 => -31857,
    46689 => -31858,
    46690 => -31858,
    46691 => -31859,
    46692 => -31860,
    46693 => -31861,
    46694 => -31861,
    46695 => -31862,
    46696 => -31863,
    46697 => -31864,
    46698 => -31864,
    46699 => -31865,
    46700 => -31866,
    46701 => -31866,
    46702 => -31867,
    46703 => -31868,
    46704 => -31869,
    46705 => -31869,
    46706 => -31870,
    46707 => -31871,
    46708 => -31872,
    46709 => -31872,
    46710 => -31873,
    46711 => -31874,
    46712 => -31875,
    46713 => -31875,
    46714 => -31876,
    46715 => -31877,
    46716 => -31877,
    46717 => -31878,
    46718 => -31879,
    46719 => -31880,
    46720 => -31880,
    46721 => -31881,
    46722 => -31882,
    46723 => -31882,
    46724 => -31883,
    46725 => -31884,
    46726 => -31885,
    46727 => -31885,
    46728 => -31886,
    46729 => -31887,
    46730 => -31888,
    46731 => -31888,
    46732 => -31889,
    46733 => -31890,
    46734 => -31890,
    46735 => -31891,
    46736 => -31892,
    46737 => -31893,
    46738 => -31893,
    46739 => -31894,
    46740 => -31895,
    46741 => -31896,
    46742 => -31896,
    46743 => -31897,
    46744 => -31898,
    46745 => -31898,
    46746 => -31899,
    46747 => -31900,
    46748 => -31901,
    46749 => -31901,
    46750 => -31902,
    46751 => -31903,
    46752 => -31903,
    46753 => -31904,
    46754 => -31905,
    46755 => -31906,
    46756 => -31906,
    46757 => -31907,
    46758 => -31908,
    46759 => -31908,
    46760 => -31909,
    46761 => -31910,
    46762 => -31911,
    46763 => -31911,
    46764 => -31912,
    46765 => -31913,
    46766 => -31913,
    46767 => -31914,
    46768 => -31915,
    46769 => -31916,
    46770 => -31916,
    46771 => -31917,
    46772 => -31918,
    46773 => -31918,
    46774 => -31919,
    46775 => -31920,
    46776 => -31921,
    46777 => -31921,
    46778 => -31922,
    46779 => -31923,
    46780 => -31923,
    46781 => -31924,
    46782 => -31925,
    46783 => -31925,
    46784 => -31926,
    46785 => -31927,
    46786 => -31928,
    46787 => -31928,
    46788 => -31929,
    46789 => -31930,
    46790 => -31930,
    46791 => -31931,
    46792 => -31932,
    46793 => -31933,
    46794 => -31933,
    46795 => -31934,
    46796 => -31935,
    46797 => -31935,
    46798 => -31936,
    46799 => -31937,
    46800 => -31937,
    46801 => -31938,
    46802 => -31939,
    46803 => -31940,
    46804 => -31940,
    46805 => -31941,
    46806 => -31942,
    46807 => -31942,
    46808 => -31943,
    46809 => -31944,
    46810 => -31944,
    46811 => -31945,
    46812 => -31946,
    46813 => -31947,
    46814 => -31947,
    46815 => -31948,
    46816 => -31949,
    46817 => -31949,
    46818 => -31950,
    46819 => -31951,
    46820 => -31951,
    46821 => -31952,
    46822 => -31953,
    46823 => -31954,
    46824 => -31954,
    46825 => -31955,
    46826 => -31956,
    46827 => -31956,
    46828 => -31957,
    46829 => -31958,
    46830 => -31958,
    46831 => -31959,
    46832 => -31960,
    46833 => -31960,
    46834 => -31961,
    46835 => -31962,
    46836 => -31963,
    46837 => -31963,
    46838 => -31964,
    46839 => -31965,
    46840 => -31965,
    46841 => -31966,
    46842 => -31967,
    46843 => -31967,
    46844 => -31968,
    46845 => -31969,
    46846 => -31969,
    46847 => -31970,
    46848 => -31971,
    46849 => -31972,
    46850 => -31972,
    46851 => -31973,
    46852 => -31974,
    46853 => -31974,
    46854 => -31975,
    46855 => -31976,
    46856 => -31976,
    46857 => -31977,
    46858 => -31978,
    46859 => -31978,
    46860 => -31979,
    46861 => -31980,
    46862 => -31980,
    46863 => -31981,
    46864 => -31982,
    46865 => -31982,
    46866 => -31983,
    46867 => -31984,
    46868 => -31985,
    46869 => -31985,
    46870 => -31986,
    46871 => -31987,
    46872 => -31987,
    46873 => -31988,
    46874 => -31989,
    46875 => -31989,
    46876 => -31990,
    46877 => -31991,
    46878 => -31991,
    46879 => -31992,
    46880 => -31993,
    46881 => -31993,
    46882 => -31994,
    46883 => -31995,
    46884 => -31995,
    46885 => -31996,
    46886 => -31997,
    46887 => -31997,
    46888 => -31998,
    46889 => -31999,
    46890 => -31999,
    46891 => -32000,
    46892 => -32001,
    46893 => -32002,
    46894 => -32002,
    46895 => -32003,
    46896 => -32004,
    46897 => -32004,
    46898 => -32005,
    46899 => -32006,
    46900 => -32006,
    46901 => -32007,
    46902 => -32008,
    46903 => -32008,
    46904 => -32009,
    46905 => -32010,
    46906 => -32010,
    46907 => -32011,
    46908 => -32012,
    46909 => -32012,
    46910 => -32013,
    46911 => -32014,
    46912 => -32014,
    46913 => -32015,
    46914 => -32016,
    46915 => -32016,
    46916 => -32017,
    46917 => -32018,
    46918 => -32018,
    46919 => -32019,
    46920 => -32020,
    46921 => -32020,
    46922 => -32021,
    46923 => -32022,
    46924 => -32022,
    46925 => -32023,
    46926 => -32024,
    46927 => -32024,
    46928 => -32025,
    46929 => -32026,
    46930 => -32026,
    46931 => -32027,
    46932 => -32028,
    46933 => -32028,
    46934 => -32029,
    46935 => -32030,
    46936 => -32030,
    46937 => -32031,
    46938 => -32032,
    46939 => -32032,
    46940 => -32033,
    46941 => -32034,
    46942 => -32034,
    46943 => -32035,
    46944 => -32036,
    46945 => -32036,
    46946 => -32037,
    46947 => -32038,
    46948 => -32038,
    46949 => -32039,
    46950 => -32040,
    46951 => -32040,
    46952 => -32041,
    46953 => -32041,
    46954 => -32042,
    46955 => -32043,
    46956 => -32043,
    46957 => -32044,
    46958 => -32045,
    46959 => -32045,
    46960 => -32046,
    46961 => -32047,
    46962 => -32047,
    46963 => -32048,
    46964 => -32049,
    46965 => -32049,
    46966 => -32050,
    46967 => -32051,
    46968 => -32051,
    46969 => -32052,
    46970 => -32053,
    46971 => -32053,
    46972 => -32054,
    46973 => -32055,
    46974 => -32055,
    46975 => -32056,
    46976 => -32057,
    46977 => -32057,
    46978 => -32058,
    46979 => -32058,
    46980 => -32059,
    46981 => -32060,
    46982 => -32060,
    46983 => -32061,
    46984 => -32062,
    46985 => -32062,
    46986 => -32063,
    46987 => -32064,
    46988 => -32064,
    46989 => -32065,
    46990 => -32066,
    46991 => -32066,
    46992 => -32067,
    46993 => -32068,
    46994 => -32068,
    46995 => -32069,
    46996 => -32069,
    46997 => -32070,
    46998 => -32071,
    46999 => -32071,
    47000 => -32072,
    47001 => -32073,
    47002 => -32073,
    47003 => -32074,
    47004 => -32075,
    47005 => -32075,
    47006 => -32076,
    47007 => -32077,
    47008 => -32077,
    47009 => -32078,
    47010 => -32078,
    47011 => -32079,
    47012 => -32080,
    47013 => -32080,
    47014 => -32081,
    47015 => -32082,
    47016 => -32082,
    47017 => -32083,
    47018 => -32084,
    47019 => -32084,
    47020 => -32085,
    47021 => -32086,
    47022 => -32086,
    47023 => -32087,
    47024 => -32087,
    47025 => -32088,
    47026 => -32089,
    47027 => -32089,
    47028 => -32090,
    47029 => -32091,
    47030 => -32091,
    47031 => -32092,
    47032 => -32092,
    47033 => -32093,
    47034 => -32094,
    47035 => -32094,
    47036 => -32095,
    47037 => -32096,
    47038 => -32096,
    47039 => -32097,
    47040 => -32098,
    47041 => -32098,
    47042 => -32099,
    47043 => -32099,
    47044 => -32100,
    47045 => -32101,
    47046 => -32101,
    47047 => -32102,
    47048 => -32103,
    47049 => -32103,
    47050 => -32104,
    47051 => -32104,
    47052 => -32105,
    47053 => -32106,
    47054 => -32106,
    47055 => -32107,
    47056 => -32108,
    47057 => -32108,
    47058 => -32109,
    47059 => -32110,
    47060 => -32110,
    47061 => -32111,
    47062 => -32111,
    47063 => -32112,
    47064 => -32113,
    47065 => -32113,
    47066 => -32114,
    47067 => -32115,
    47068 => -32115,
    47069 => -32116,
    47070 => -32116,
    47071 => -32117,
    47072 => -32118,
    47073 => -32118,
    47074 => -32119,
    47075 => -32119,
    47076 => -32120,
    47077 => -32121,
    47078 => -32121,
    47079 => -32122,
    47080 => -32123,
    47081 => -32123,
    47082 => -32124,
    47083 => -32124,
    47084 => -32125,
    47085 => -32126,
    47086 => -32126,
    47087 => -32127,
    47088 => -32128,
    47089 => -32128,
    47090 => -32129,
    47091 => -32129,
    47092 => -32130,
    47093 => -32131,
    47094 => -32131,
    47095 => -32132,
    47096 => -32132,
    47097 => -32133,
    47098 => -32134,
    47099 => -32134,
    47100 => -32135,
    47101 => -32136,
    47102 => -32136,
    47103 => -32137,
    47104 => -32137,
    47105 => -32138,
    47106 => -32139,
    47107 => -32139,
    47108 => -32140,
    47109 => -32140,
    47110 => -32141,
    47111 => -32142,
    47112 => -32142,
    47113 => -32143,
    47114 => -32144,
    47115 => -32144,
    47116 => -32145,
    47117 => -32145,
    47118 => -32146,
    47119 => -32147,
    47120 => -32147,
    47121 => -32148,
    47122 => -32148,
    47123 => -32149,
    47124 => -32150,
    47125 => -32150,
    47126 => -32151,
    47127 => -32151,
    47128 => -32152,
    47129 => -32153,
    47130 => -32153,
    47131 => -32154,
    47132 => -32154,
    47133 => -32155,
    47134 => -32156,
    47135 => -32156,
    47136 => -32157,
    47137 => -32157,
    47138 => -32158,
    47139 => -32159,
    47140 => -32159,
    47141 => -32160,
    47142 => -32160,
    47143 => -32161,
    47144 => -32162,
    47145 => -32162,
    47146 => -32163,
    47147 => -32163,
    47148 => -32164,
    47149 => -32165,
    47150 => -32165,
    47151 => -32166,
    47152 => -32166,
    47153 => -32167,
    47154 => -32168,
    47155 => -32168,
    47156 => -32169,
    47157 => -32169,
    47158 => -32170,
    47159 => -32171,
    47160 => -32171,
    47161 => -32172,
    47162 => -32172,
    47163 => -32173,
    47164 => -32174,
    47165 => -32174,
    47166 => -32175,
    47167 => -32175,
    47168 => -32176,
    47169 => -32177,
    47170 => -32177,
    47171 => -32178,
    47172 => -32178,
    47173 => -32179,
    47174 => -32180,
    47175 => -32180,
    47176 => -32181,
    47177 => -32181,
    47178 => -32182,
    47179 => -32183,
    47180 => -32183,
    47181 => -32184,
    47182 => -32184,
    47183 => -32185,
    47184 => -32185,
    47185 => -32186,
    47186 => -32187,
    47187 => -32187,
    47188 => -32188,
    47189 => -32188,
    47190 => -32189,
    47191 => -32190,
    47192 => -32190,
    47193 => -32191,
    47194 => -32191,
    47195 => -32192,
    47196 => -32193,
    47197 => -32193,
    47198 => -32194,
    47199 => -32194,
    47200 => -32195,
    47201 => -32195,
    47202 => -32196,
    47203 => -32197,
    47204 => -32197,
    47205 => -32198,
    47206 => -32198,
    47207 => -32199,
    47208 => -32200,
    47209 => -32200,
    47210 => -32201,
    47211 => -32201,
    47212 => -32202,
    47213 => -32202,
    47214 => -32203,
    47215 => -32204,
    47216 => -32204,
    47217 => -32205,
    47218 => -32205,
    47219 => -32206,
    47220 => -32206,
    47221 => -32207,
    47222 => -32208,
    47223 => -32208,
    47224 => -32209,
    47225 => -32209,
    47226 => -32210,
    47227 => -32211,
    47228 => -32211,
    47229 => -32212,
    47230 => -32212,
    47231 => -32213,
    47232 => -32213,
    47233 => -32214,
    47234 => -32215,
    47235 => -32215,
    47236 => -32216,
    47237 => -32216,
    47238 => -32217,
    47239 => -32217,
    47240 => -32218,
    47241 => -32219,
    47242 => -32219,
    47243 => -32220,
    47244 => -32220,
    47245 => -32221,
    47246 => -32221,
    47247 => -32222,
    47248 => -32223,
    47249 => -32223,
    47250 => -32224,
    47251 => -32224,
    47252 => -32225,
    47253 => -32225,
    47254 => -32226,
    47255 => -32227,
    47256 => -32227,
    47257 => -32228,
    47258 => -32228,
    47259 => -32229,
    47260 => -32229,
    47261 => -32230,
    47262 => -32231,
    47263 => -32231,
    47264 => -32232,
    47265 => -32232,
    47266 => -32233,
    47267 => -32233,
    47268 => -32234,
    47269 => -32234,
    47270 => -32235,
    47271 => -32236,
    47272 => -32236,
    47273 => -32237,
    47274 => -32237,
    47275 => -32238,
    47276 => -32238,
    47277 => -32239,
    47278 => -32240,
    47279 => -32240,
    47280 => -32241,
    47281 => -32241,
    47282 => -32242,
    47283 => -32242,
    47284 => -32243,
    47285 => -32243,
    47286 => -32244,
    47287 => -32245,
    47288 => -32245,
    47289 => -32246,
    47290 => -32246,
    47291 => -32247,
    47292 => -32247,
    47293 => -32248,
    47294 => -32248,
    47295 => -32249,
    47296 => -32250,
    47297 => -32250,
    47298 => -32251,
    47299 => -32251,
    47300 => -32252,
    47301 => -32252,
    47302 => -32253,
    47303 => -32253,
    47304 => -32254,
    47305 => -32255,
    47306 => -32255,
    47307 => -32256,
    47308 => -32256,
    47309 => -32257,
    47310 => -32257,
    47311 => -32258,
    47312 => -32258,
    47313 => -32259,
    47314 => -32260,
    47315 => -32260,
    47316 => -32261,
    47317 => -32261,
    47318 => -32262,
    47319 => -32262,
    47320 => -32263,
    47321 => -32263,
    47322 => -32264,
    47323 => -32265,
    47324 => -32265,
    47325 => -32266,
    47326 => -32266,
    47327 => -32267,
    47328 => -32267,
    47329 => -32268,
    47330 => -32268,
    47331 => -32269,
    47332 => -32269,
    47333 => -32270,
    47334 => -32271,
    47335 => -32271,
    47336 => -32272,
    47337 => -32272,
    47338 => -32273,
    47339 => -32273,
    47340 => -32274,
    47341 => -32274,
    47342 => -32275,
    47343 => -32275,
    47344 => -32276,
    47345 => -32277,
    47346 => -32277,
    47347 => -32278,
    47348 => -32278,
    47349 => -32279,
    47350 => -32279,
    47351 => -32280,
    47352 => -32280,
    47353 => -32281,
    47354 => -32281,
    47355 => -32282,
    47356 => -32282,
    47357 => -32283,
    47358 => -32284,
    47359 => -32284,
    47360 => -32285,
    47361 => -32285,
    47362 => -32286,
    47363 => -32286,
    47364 => -32287,
    47365 => -32287,
    47366 => -32288,
    47367 => -32288,
    47368 => -32289,
    47369 => -32289,
    47370 => -32290,
    47371 => -32290,
    47372 => -32291,
    47373 => -32292,
    47374 => -32292,
    47375 => -32293,
    47376 => -32293,
    47377 => -32294,
    47378 => -32294,
    47379 => -32295,
    47380 => -32295,
    47381 => -32296,
    47382 => -32296,
    47383 => -32297,
    47384 => -32297,
    47385 => -32298,
    47386 => -32298,
    47387 => -32299,
    47388 => -32300,
    47389 => -32300,
    47390 => -32301,
    47391 => -32301,
    47392 => -32302,
    47393 => -32302,
    47394 => -32303,
    47395 => -32303,
    47396 => -32304,
    47397 => -32304,
    47398 => -32305,
    47399 => -32305,
    47400 => -32306,
    47401 => -32306,
    47402 => -32307,
    47403 => -32307,
    47404 => -32308,
    47405 => -32308,
    47406 => -32309,
    47407 => -32310,
    47408 => -32310,
    47409 => -32311,
    47410 => -32311,
    47411 => -32312,
    47412 => -32312,
    47413 => -32313,
    47414 => -32313,
    47415 => -32314,
    47416 => -32314,
    47417 => -32315,
    47418 => -32315,
    47419 => -32316,
    47420 => -32316,
    47421 => -32317,
    47422 => -32317,
    47423 => -32318,
    47424 => -32318,
    47425 => -32319,
    47426 => -32319,
    47427 => -32320,
    47428 => -32320,
    47429 => -32321,
    47430 => -32321,
    47431 => -32322,
    47432 => -32322,
    47433 => -32323,
    47434 => -32324,
    47435 => -32324,
    47436 => -32325,
    47437 => -32325,
    47438 => -32326,
    47439 => -32326,
    47440 => -32327,
    47441 => -32327,
    47442 => -32328,
    47443 => -32328,
    47444 => -32329,
    47445 => -32329,
    47446 => -32330,
    47447 => -32330,
    47448 => -32331,
    47449 => -32331,
    47450 => -32332,
    47451 => -32332,
    47452 => -32333,
    47453 => -32333,
    47454 => -32334,
    47455 => -32334,
    47456 => -32335,
    47457 => -32335,
    47458 => -32336,
    47459 => -32336,
    47460 => -32337,
    47461 => -32337,
    47462 => -32338,
    47463 => -32338,
    47464 => -32339,
    47465 => -32339,
    47466 => -32340,
    47467 => -32340,
    47468 => -32341,
    47469 => -32341,
    47470 => -32342,
    47471 => -32342,
    47472 => -32343,
    47473 => -32343,
    47474 => -32344,
    47475 => -32344,
    47476 => -32345,
    47477 => -32345,
    47478 => -32346,
    47479 => -32346,
    47480 => -32347,
    47481 => -32347,
    47482 => -32348,
    47483 => -32348,
    47484 => -32349,
    47485 => -32349,
    47486 => -32350,
    47487 => -32350,
    47488 => -32351,
    47489 => -32351,
    47490 => -32352,
    47491 => -32352,
    47492 => -32353,
    47493 => -32353,
    47494 => -32354,
    47495 => -32354,
    47496 => -32355,
    47497 => -32355,
    47498 => -32356,
    47499 => -32356,
    47500 => -32357,
    47501 => -32357,
    47502 => -32358,
    47503 => -32358,
    47504 => -32359,
    47505 => -32359,
    47506 => -32360,
    47507 => -32360,
    47508 => -32361,
    47509 => -32361,
    47510 => -32362,
    47511 => -32362,
    47512 => -32363,
    47513 => -32363,
    47514 => -32364,
    47515 => -32364,
    47516 => -32365,
    47517 => -32365,
    47518 => -32366,
    47519 => -32366,
    47520 => -32367,
    47521 => -32367,
    47522 => -32368,
    47523 => -32368,
    47524 => -32369,
    47525 => -32369,
    47526 => -32370,
    47527 => -32370,
    47528 => -32371,
    47529 => -32371,
    47530 => -32372,
    47531 => -32372,
    47532 => -32373,
    47533 => -32373,
    47534 => -32374,
    47535 => -32374,
    47536 => -32375,
    47537 => -32375,
    47538 => -32375,
    47539 => -32376,
    47540 => -32376,
    47541 => -32377,
    47542 => -32377,
    47543 => -32378,
    47544 => -32378,
    47545 => -32379,
    47546 => -32379,
    47547 => -32380,
    47548 => -32380,
    47549 => -32381,
    47550 => -32381,
    47551 => -32382,
    47552 => -32382,
    47553 => -32383,
    47554 => -32383,
    47555 => -32384,
    47556 => -32384,
    47557 => -32385,
    47558 => -32385,
    47559 => -32386,
    47560 => -32386,
    47561 => -32387,
    47562 => -32387,
    47563 => -32387,
    47564 => -32388,
    47565 => -32388,
    47566 => -32389,
    47567 => -32389,
    47568 => -32390,
    47569 => -32390,
    47570 => -32391,
    47571 => -32391,
    47572 => -32392,
    47573 => -32392,
    47574 => -32393,
    47575 => -32393,
    47576 => -32394,
    47577 => -32394,
    47578 => -32395,
    47579 => -32395,
    47580 => -32396,
    47581 => -32396,
    47582 => -32397,
    47583 => -32397,
    47584 => -32397,
    47585 => -32398,
    47586 => -32398,
    47587 => -32399,
    47588 => -32399,
    47589 => -32400,
    47590 => -32400,
    47591 => -32401,
    47592 => -32401,
    47593 => -32402,
    47594 => -32402,
    47595 => -32403,
    47596 => -32403,
    47597 => -32404,
    47598 => -32404,
    47599 => -32404,
    47600 => -32405,
    47601 => -32405,
    47602 => -32406,
    47603 => -32406,
    47604 => -32407,
    47605 => -32407,
    47606 => -32408,
    47607 => -32408,
    47608 => -32409,
    47609 => -32409,
    47610 => -32410,
    47611 => -32410,
    47612 => -32411,
    47613 => -32411,
    47614 => -32411,
    47615 => -32412,
    47616 => -32412,
    47617 => -32413,
    47618 => -32413,
    47619 => -32414,
    47620 => -32414,
    47621 => -32415,
    47622 => -32415,
    47623 => -32416,
    47624 => -32416,
    47625 => -32416,
    47626 => -32417,
    47627 => -32417,
    47628 => -32418,
    47629 => -32418,
    47630 => -32419,
    47631 => -32419,
    47632 => -32420,
    47633 => -32420,
    47634 => -32421,
    47635 => -32421,
    47636 => -32422,
    47637 => -32422,
    47638 => -32422,
    47639 => -32423,
    47640 => -32423,
    47641 => -32424,
    47642 => -32424,
    47643 => -32425,
    47644 => -32425,
    47645 => -32426,
    47646 => -32426,
    47647 => -32426,
    47648 => -32427,
    47649 => -32427,
    47650 => -32428,
    47651 => -32428,
    47652 => -32429,
    47653 => -32429,
    47654 => -32430,
    47655 => -32430,
    47656 => -32431,
    47657 => -32431,
    47658 => -32431,
    47659 => -32432,
    47660 => -32432,
    47661 => -32433,
    47662 => -32433,
    47663 => -32434,
    47664 => -32434,
    47665 => -32435,
    47666 => -32435,
    47667 => -32435,
    47668 => -32436,
    47669 => -32436,
    47670 => -32437,
    47671 => -32437,
    47672 => -32438,
    47673 => -32438,
    47674 => -32439,
    47675 => -32439,
    47676 => -32439,
    47677 => -32440,
    47678 => -32440,
    47679 => -32441,
    47680 => -32441,
    47681 => -32442,
    47682 => -32442,
    47683 => -32443,
    47684 => -32443,
    47685 => -32443,
    47686 => -32444,
    47687 => -32444,
    47688 => -32445,
    47689 => -32445,
    47690 => -32446,
    47691 => -32446,
    47692 => -32447,
    47693 => -32447,
    47694 => -32447,
    47695 => -32448,
    47696 => -32448,
    47697 => -32449,
    47698 => -32449,
    47699 => -32450,
    47700 => -32450,
    47701 => -32450,
    47702 => -32451,
    47703 => -32451,
    47704 => -32452,
    47705 => -32452,
    47706 => -32453,
    47707 => -32453,
    47708 => -32453,
    47709 => -32454,
    47710 => -32454,
    47711 => -32455,
    47712 => -32455,
    47713 => -32456,
    47714 => -32456,
    47715 => -32457,
    47716 => -32457,
    47717 => -32457,
    47718 => -32458,
    47719 => -32458,
    47720 => -32459,
    47721 => -32459,
    47722 => -32460,
    47723 => -32460,
    47724 => -32460,
    47725 => -32461,
    47726 => -32461,
    47727 => -32462,
    47728 => -32462,
    47729 => -32463,
    47730 => -32463,
    47731 => -32463,
    47732 => -32464,
    47733 => -32464,
    47734 => -32465,
    47735 => -32465,
    47736 => -32466,
    47737 => -32466,
    47738 => -32466,
    47739 => -32467,
    47740 => -32467,
    47741 => -32468,
    47742 => -32468,
    47743 => -32468,
    47744 => -32469,
    47745 => -32469,
    47746 => -32470,
    47747 => -32470,
    47748 => -32471,
    47749 => -32471,
    47750 => -32471,
    47751 => -32472,
    47752 => -32472,
    47753 => -32473,
    47754 => -32473,
    47755 => -32474,
    47756 => -32474,
    47757 => -32474,
    47758 => -32475,
    47759 => -32475,
    47760 => -32476,
    47761 => -32476,
    47762 => -32476,
    47763 => -32477,
    47764 => -32477,
    47765 => -32478,
    47766 => -32478,
    47767 => -32479,
    47768 => -32479,
    47769 => -32479,
    47770 => -32480,
    47771 => -32480,
    47772 => -32481,
    47773 => -32481,
    47774 => -32481,
    47775 => -32482,
    47776 => -32482,
    47777 => -32483,
    47778 => -32483,
    47779 => -32484,
    47780 => -32484,
    47781 => -32484,
    47782 => -32485,
    47783 => -32485,
    47784 => -32486,
    47785 => -32486,
    47786 => -32486,
    47787 => -32487,
    47788 => -32487,
    47789 => -32488,
    47790 => -32488,
    47791 => -32488,
    47792 => -32489,
    47793 => -32489,
    47794 => -32490,
    47795 => -32490,
    47796 => -32490,
    47797 => -32491,
    47798 => -32491,
    47799 => -32492,
    47800 => -32492,
    47801 => -32493,
    47802 => -32493,
    47803 => -32493,
    47804 => -32494,
    47805 => -32494,
    47806 => -32495,
    47807 => -32495,
    47808 => -32495,
    47809 => -32496,
    47810 => -32496,
    47811 => -32497,
    47812 => -32497,
    47813 => -32497,
    47814 => -32498,
    47815 => -32498,
    47816 => -32499,
    47817 => -32499,
    47818 => -32499,
    47819 => -32500,
    47820 => -32500,
    47821 => -32501,
    47822 => -32501,
    47823 => -32501,
    47824 => -32502,
    47825 => -32502,
    47826 => -32503,
    47827 => -32503,
    47828 => -32503,
    47829 => -32504,
    47830 => -32504,
    47831 => -32505,
    47832 => -32505,
    47833 => -32505,
    47834 => -32506,
    47835 => -32506,
    47836 => -32507,
    47837 => -32507,
    47838 => -32507,
    47839 => -32508,
    47840 => -32508,
    47841 => -32509,
    47842 => -32509,
    47843 => -32509,
    47844 => -32510,
    47845 => -32510,
    47846 => -32510,
    47847 => -32511,
    47848 => -32511,
    47849 => -32512,
    47850 => -32512,
    47851 => -32512,
    47852 => -32513,
    47853 => -32513,
    47854 => -32514,
    47855 => -32514,
    47856 => -32514,
    47857 => -32515,
    47858 => -32515,
    47859 => -32516,
    47860 => -32516,
    47861 => -32516,
    47862 => -32517,
    47863 => -32517,
    47864 => -32517,
    47865 => -32518,
    47866 => -32518,
    47867 => -32519,
    47868 => -32519,
    47869 => -32519,
    47870 => -32520,
    47871 => -32520,
    47872 => -32521,
    47873 => -32521,
    47874 => -32521,
    47875 => -32522,
    47876 => -32522,
    47877 => -32522,
    47878 => -32523,
    47879 => -32523,
    47880 => -32524,
    47881 => -32524,
    47882 => -32524,
    47883 => -32525,
    47884 => -32525,
    47885 => -32526,
    47886 => -32526,
    47887 => -32526,
    47888 => -32527,
    47889 => -32527,
    47890 => -32527,
    47891 => -32528,
    47892 => -32528,
    47893 => -32529,
    47894 => -32529,
    47895 => -32529,
    47896 => -32530,
    47897 => -32530,
    47898 => -32530,
    47899 => -32531,
    47900 => -32531,
    47901 => -32532,
    47902 => -32532,
    47903 => -32532,
    47904 => -32533,
    47905 => -32533,
    47906 => -32533,
    47907 => -32534,
    47908 => -32534,
    47909 => -32535,
    47910 => -32535,
    47911 => -32535,
    47912 => -32536,
    47913 => -32536,
    47914 => -32536,
    47915 => -32537,
    47916 => -32537,
    47917 => -32538,
    47918 => -32538,
    47919 => -32538,
    47920 => -32539,
    47921 => -32539,
    47922 => -32539,
    47923 => -32540,
    47924 => -32540,
    47925 => -32541,
    47926 => -32541,
    47927 => -32541,
    47928 => -32542,
    47929 => -32542,
    47930 => -32542,
    47931 => -32543,
    47932 => -32543,
    47933 => -32543,
    47934 => -32544,
    47935 => -32544,
    47936 => -32545,
    47937 => -32545,
    47938 => -32545,
    47939 => -32546,
    47940 => -32546,
    47941 => -32546,
    47942 => -32547,
    47943 => -32547,
    47944 => -32547,
    47945 => -32548,
    47946 => -32548,
    47947 => -32549,
    47948 => -32549,
    47949 => -32549,
    47950 => -32550,
    47951 => -32550,
    47952 => -32550,
    47953 => -32551,
    47954 => -32551,
    47955 => -32551,
    47956 => -32552,
    47957 => -32552,
    47958 => -32553,
    47959 => -32553,
    47960 => -32553,
    47961 => -32554,
    47962 => -32554,
    47963 => -32554,
    47964 => -32555,
    47965 => -32555,
    47966 => -32555,
    47967 => -32556,
    47968 => -32556,
    47969 => -32556,
    47970 => -32557,
    47971 => -32557,
    47972 => -32558,
    47973 => -32558,
    47974 => -32558,
    47975 => -32559,
    47976 => -32559,
    47977 => -32559,
    47978 => -32560,
    47979 => -32560,
    47980 => -32560,
    47981 => -32561,
    47982 => -32561,
    47983 => -32561,
    47984 => -32562,
    47985 => -32562,
    47986 => -32562,
    47987 => -32563,
    47988 => -32563,
    47989 => -32564,
    47990 => -32564,
    47991 => -32564,
    47992 => -32565,
    47993 => -32565,
    47994 => -32565,
    47995 => -32566,
    47996 => -32566,
    47997 => -32566,
    47998 => -32567,
    47999 => -32567,
    48000 => -32567,
    48001 => -32568,
    48002 => -32568,
    48003 => -32568,
    48004 => -32569,
    48005 => -32569,
    48006 => -32569,
    48007 => -32570,
    48008 => -32570,
    48009 => -32570,
    48010 => -32571,
    48011 => -32571,
    48012 => -32571,
    48013 => -32572,
    48014 => -32572,
    48015 => -32573,
    48016 => -32573,
    48017 => -32573,
    48018 => -32574,
    48019 => -32574,
    48020 => -32574,
    48021 => -32575,
    48022 => -32575,
    48023 => -32575,
    48024 => -32576,
    48025 => -32576,
    48026 => -32576,
    48027 => -32577,
    48028 => -32577,
    48029 => -32577,
    48030 => -32578,
    48031 => -32578,
    48032 => -32578,
    48033 => -32579,
    48034 => -32579,
    48035 => -32579,
    48036 => -32580,
    48037 => -32580,
    48038 => -32580,
    48039 => -32581,
    48040 => -32581,
    48041 => -32581,
    48042 => -32582,
    48043 => -32582,
    48044 => -32582,
    48045 => -32583,
    48046 => -32583,
    48047 => -32583,
    48048 => -32584,
    48049 => -32584,
    48050 => -32584,
    48051 => -32585,
    48052 => -32585,
    48053 => -32585,
    48054 => -32586,
    48055 => -32586,
    48056 => -32586,
    48057 => -32587,
    48058 => -32587,
    48059 => -32587,
    48060 => -32588,
    48061 => -32588,
    48062 => -32588,
    48063 => -32589,
    48064 => -32589,
    48065 => -32589,
    48066 => -32590,
    48067 => -32590,
    48068 => -32590,
    48069 => -32591,
    48070 => -32591,
    48071 => -32591,
    48072 => -32592,
    48073 => -32592,
    48074 => -32592,
    48075 => -32592,
    48076 => -32593,
    48077 => -32593,
    48078 => -32593,
    48079 => -32594,
    48080 => -32594,
    48081 => -32594,
    48082 => -32595,
    48083 => -32595,
    48084 => -32595,
    48085 => -32596,
    48086 => -32596,
    48087 => -32596,
    48088 => -32597,
    48089 => -32597,
    48090 => -32597,
    48091 => -32598,
    48092 => -32598,
    48093 => -32598,
    48094 => -32599,
    48095 => -32599,
    48096 => -32599,
    48097 => -32600,
    48098 => -32600,
    48099 => -32600,
    48100 => -32600,
    48101 => -32601,
    48102 => -32601,
    48103 => -32601,
    48104 => -32602,
    48105 => -32602,
    48106 => -32602,
    48107 => -32603,
    48108 => -32603,
    48109 => -32603,
    48110 => -32604,
    48111 => -32604,
    48112 => -32604,
    48113 => -32605,
    48114 => -32605,
    48115 => -32605,
    48116 => -32606,
    48117 => -32606,
    48118 => -32606,
    48119 => -32606,
    48120 => -32607,
    48121 => -32607,
    48122 => -32607,
    48123 => -32608,
    48124 => -32608,
    48125 => -32608,
    48126 => -32609,
    48127 => -32609,
    48128 => -32609,
    48129 => -32610,
    48130 => -32610,
    48131 => -32610,
    48132 => -32610,
    48133 => -32611,
    48134 => -32611,
    48135 => -32611,
    48136 => -32612,
    48137 => -32612,
    48138 => -32612,
    48139 => -32613,
    48140 => -32613,
    48141 => -32613,
    48142 => -32613,
    48143 => -32614,
    48144 => -32614,
    48145 => -32614,
    48146 => -32615,
    48147 => -32615,
    48148 => -32615,
    48149 => -32616,
    48150 => -32616,
    48151 => -32616,
    48152 => -32617,
    48153 => -32617,
    48154 => -32617,
    48155 => -32617,
    48156 => -32618,
    48157 => -32618,
    48158 => -32618,
    48159 => -32619,
    48160 => -32619,
    48161 => -32619,
    48162 => -32620,
    48163 => -32620,
    48164 => -32620,
    48165 => -32620,
    48166 => -32621,
    48167 => -32621,
    48168 => -32621,
    48169 => -32622,
    48170 => -32622,
    48171 => -32622,
    48172 => -32622,
    48173 => -32623,
    48174 => -32623,
    48175 => -32623,
    48176 => -32624,
    48177 => -32624,
    48178 => -32624,
    48179 => -32625,
    48180 => -32625,
    48181 => -32625,
    48182 => -32625,
    48183 => -32626,
    48184 => -32626,
    48185 => -32626,
    48186 => -32627,
    48187 => -32627,
    48188 => -32627,
    48189 => -32627,
    48190 => -32628,
    48191 => -32628,
    48192 => -32628,
    48193 => -32629,
    48194 => -32629,
    48195 => -32629,
    48196 => -32629,
    48197 => -32630,
    48198 => -32630,
    48199 => -32630,
    48200 => -32631,
    48201 => -32631,
    48202 => -32631,
    48203 => -32631,
    48204 => -32632,
    48205 => -32632,
    48206 => -32632,
    48207 => -32633,
    48208 => -32633,
    48209 => -32633,
    48210 => -32633,
    48211 => -32634,
    48212 => -32634,
    48213 => -32634,
    48214 => -32635,
    48215 => -32635,
    48216 => -32635,
    48217 => -32635,
    48218 => -32636,
    48219 => -32636,
    48220 => -32636,
    48221 => -32637,
    48222 => -32637,
    48223 => -32637,
    48224 => -32637,
    48225 => -32638,
    48226 => -32638,
    48227 => -32638,
    48228 => -32639,
    48229 => -32639,
    48230 => -32639,
    48231 => -32639,
    48232 => -32640,
    48233 => -32640,
    48234 => -32640,
    48235 => -32640,
    48236 => -32641,
    48237 => -32641,
    48238 => -32641,
    48239 => -32642,
    48240 => -32642,
    48241 => -32642,
    48242 => -32642,
    48243 => -32643,
    48244 => -32643,
    48245 => -32643,
    48246 => -32643,
    48247 => -32644,
    48248 => -32644,
    48249 => -32644,
    48250 => -32645,
    48251 => -32645,
    48252 => -32645,
    48253 => -32645,
    48254 => -32646,
    48255 => -32646,
    48256 => -32646,
    48257 => -32646,
    48258 => -32647,
    48259 => -32647,
    48260 => -32647,
    48261 => -32648,
    48262 => -32648,
    48263 => -32648,
    48264 => -32648,
    48265 => -32649,
    48266 => -32649,
    48267 => -32649,
    48268 => -32649,
    48269 => -32650,
    48270 => -32650,
    48271 => -32650,
    48272 => -32650,
    48273 => -32651,
    48274 => -32651,
    48275 => -32651,
    48276 => -32652,
    48277 => -32652,
    48278 => -32652,
    48279 => -32652,
    48280 => -32653,
    48281 => -32653,
    48282 => -32653,
    48283 => -32653,
    48284 => -32654,
    48285 => -32654,
    48286 => -32654,
    48287 => -32654,
    48288 => -32655,
    48289 => -32655,
    48290 => -32655,
    48291 => -32655,
    48292 => -32656,
    48293 => -32656,
    48294 => -32656,
    48295 => -32656,
    48296 => -32657,
    48297 => -32657,
    48298 => -32657,
    48299 => -32657,
    48300 => -32658,
    48301 => -32658,
    48302 => -32658,
    48303 => -32659,
    48304 => -32659,
    48305 => -32659,
    48306 => -32659,
    48307 => -32660,
    48308 => -32660,
    48309 => -32660,
    48310 => -32660,
    48311 => -32661,
    48312 => -32661,
    48313 => -32661,
    48314 => -32661,
    48315 => -32662,
    48316 => -32662,
    48317 => -32662,
    48318 => -32662,
    48319 => -32663,
    48320 => -32663,
    48321 => -32663,
    48322 => -32663,
    48323 => -32664,
    48324 => -32664,
    48325 => -32664,
    48326 => -32664,
    48327 => -32665,
    48328 => -32665,
    48329 => -32665,
    48330 => -32665,
    48331 => -32666,
    48332 => -32666,
    48333 => -32666,
    48334 => -32666,
    48335 => -32667,
    48336 => -32667,
    48337 => -32667,
    48338 => -32667,
    48339 => -32668,
    48340 => -32668,
    48341 => -32668,
    48342 => -32668,
    48343 => -32668,
    48344 => -32669,
    48345 => -32669,
    48346 => -32669,
    48347 => -32669,
    48348 => -32670,
    48349 => -32670,
    48350 => -32670,
    48351 => -32670,
    48352 => -32671,
    48353 => -32671,
    48354 => -32671,
    48355 => -32671,
    48356 => -32672,
    48357 => -32672,
    48358 => -32672,
    48359 => -32672,
    48360 => -32673,
    48361 => -32673,
    48362 => -32673,
    48363 => -32673,
    48364 => -32674,
    48365 => -32674,
    48366 => -32674,
    48367 => -32674,
    48368 => -32674,
    48369 => -32675,
    48370 => -32675,
    48371 => -32675,
    48372 => -32675,
    48373 => -32676,
    48374 => -32676,
    48375 => -32676,
    48376 => -32676,
    48377 => -32677,
    48378 => -32677,
    48379 => -32677,
    48380 => -32677,
    48381 => -32678,
    48382 => -32678,
    48383 => -32678,
    48384 => -32678,
    48385 => -32678,
    48386 => -32679,
    48387 => -32679,
    48388 => -32679,
    48389 => -32679,
    48390 => -32680,
    48391 => -32680,
    48392 => -32680,
    48393 => -32680,
    48394 => -32681,
    48395 => -32681,
    48396 => -32681,
    48397 => -32681,
    48398 => -32681,
    48399 => -32682,
    48400 => -32682,
    48401 => -32682,
    48402 => -32682,
    48403 => -32683,
    48404 => -32683,
    48405 => -32683,
    48406 => -32683,
    48407 => -32683,
    48408 => -32684,
    48409 => -32684,
    48410 => -32684,
    48411 => -32684,
    48412 => -32685,
    48413 => -32685,
    48414 => -32685,
    48415 => -32685,
    48416 => -32685,
    48417 => -32686,
    48418 => -32686,
    48419 => -32686,
    48420 => -32686,
    48421 => -32687,
    48422 => -32687,
    48423 => -32687,
    48424 => -32687,
    48425 => -32687,
    48426 => -32688,
    48427 => -32688,
    48428 => -32688,
    48429 => -32688,
    48430 => -32689,
    48431 => -32689,
    48432 => -32689,
    48433 => -32689,
    48434 => -32689,
    48435 => -32690,
    48436 => -32690,
    48437 => -32690,
    48438 => -32690,
    48439 => -32690,
    48440 => -32691,
    48441 => -32691,
    48442 => -32691,
    48443 => -32691,
    48444 => -32692,
    48445 => -32692,
    48446 => -32692,
    48447 => -32692,
    48448 => -32692,
    48449 => -32693,
    48450 => -32693,
    48451 => -32693,
    48452 => -32693,
    48453 => -32693,
    48454 => -32694,
    48455 => -32694,
    48456 => -32694,
    48457 => -32694,
    48458 => -32694,
    48459 => -32695,
    48460 => -32695,
    48461 => -32695,
    48462 => -32695,
    48463 => -32696,
    48464 => -32696,
    48465 => -32696,
    48466 => -32696,
    48467 => -32696,
    48468 => -32697,
    48469 => -32697,
    48470 => -32697,
    48471 => -32697,
    48472 => -32697,
    48473 => -32698,
    48474 => -32698,
    48475 => -32698,
    48476 => -32698,
    48477 => -32698,
    48478 => -32699,
    48479 => -32699,
    48480 => -32699,
    48481 => -32699,
    48482 => -32699,
    48483 => -32700,
    48484 => -32700,
    48485 => -32700,
    48486 => -32700,
    48487 => -32700,
    48488 => -32701,
    48489 => -32701,
    48490 => -32701,
    48491 => -32701,
    48492 => -32701,
    48493 => -32702,
    48494 => -32702,
    48495 => -32702,
    48496 => -32702,
    48497 => -32702,
    48498 => -32703,
    48499 => -32703,
    48500 => -32703,
    48501 => -32703,
    48502 => -32703,
    48503 => -32704,
    48504 => -32704,
    48505 => -32704,
    48506 => -32704,
    48507 => -32704,
    48508 => -32705,
    48509 => -32705,
    48510 => -32705,
    48511 => -32705,
    48512 => -32705,
    48513 => -32706,
    48514 => -32706,
    48515 => -32706,
    48516 => -32706,
    48517 => -32706,
    48518 => -32706,
    48519 => -32707,
    48520 => -32707,
    48521 => -32707,
    48522 => -32707,
    48523 => -32707,
    48524 => -32708,
    48525 => -32708,
    48526 => -32708,
    48527 => -32708,
    48528 => -32708,
    48529 => -32709,
    48530 => -32709,
    48531 => -32709,
    48532 => -32709,
    48533 => -32709,
    48534 => -32710,
    48535 => -32710,
    48536 => -32710,
    48537 => -32710,
    48538 => -32710,
    48539 => -32710,
    48540 => -32711,
    48541 => -32711,
    48542 => -32711,
    48543 => -32711,
    48544 => -32711,
    48545 => -32712,
    48546 => -32712,
    48547 => -32712,
    48548 => -32712,
    48549 => -32712,
    48550 => -32712,
    48551 => -32713,
    48552 => -32713,
    48553 => -32713,
    48554 => -32713,
    48555 => -32713,
    48556 => -32714,
    48557 => -32714,
    48558 => -32714,
    48559 => -32714,
    48560 => -32714,
    48561 => -32714,
    48562 => -32715,
    48563 => -32715,
    48564 => -32715,
    48565 => -32715,
    48566 => -32715,
    48567 => -32715,
    48568 => -32716,
    48569 => -32716,
    48570 => -32716,
    48571 => -32716,
    48572 => -32716,
    48573 => -32717,
    48574 => -32717,
    48575 => -32717,
    48576 => -32717,
    48577 => -32717,
    48578 => -32717,
    48579 => -32718,
    48580 => -32718,
    48581 => -32718,
    48582 => -32718,
    48583 => -32718,
    48584 => -32718,
    48585 => -32719,
    48586 => -32719,
    48587 => -32719,
    48588 => -32719,
    48589 => -32719,
    48590 => -32719,
    48591 => -32720,
    48592 => -32720,
    48593 => -32720,
    48594 => -32720,
    48595 => -32720,
    48596 => -32720,
    48597 => -32721,
    48598 => -32721,
    48599 => -32721,
    48600 => -32721,
    48601 => -32721,
    48602 => -32721,
    48603 => -32722,
    48604 => -32722,
    48605 => -32722,
    48606 => -32722,
    48607 => -32722,
    48608 => -32722,
    48609 => -32723,
    48610 => -32723,
    48611 => -32723,
    48612 => -32723,
    48613 => -32723,
    48614 => -32723,
    48615 => -32724,
    48616 => -32724,
    48617 => -32724,
    48618 => -32724,
    48619 => -32724,
    48620 => -32724,
    48621 => -32725,
    48622 => -32725,
    48623 => -32725,
    48624 => -32725,
    48625 => -32725,
    48626 => -32725,
    48627 => -32726,
    48628 => -32726,
    48629 => -32726,
    48630 => -32726,
    48631 => -32726,
    48632 => -32726,
    48633 => -32726,
    48634 => -32727,
    48635 => -32727,
    48636 => -32727,
    48637 => -32727,
    48638 => -32727,
    48639 => -32727,
    48640 => -32728,
    48641 => -32728,
    48642 => -32728,
    48643 => -32728,
    48644 => -32728,
    48645 => -32728,
    48646 => -32728,
    48647 => -32729,
    48648 => -32729,
    48649 => -32729,
    48650 => -32729,
    48651 => -32729,
    48652 => -32729,
    48653 => -32730,
    48654 => -32730,
    48655 => -32730,
    48656 => -32730,
    48657 => -32730,
    48658 => -32730,
    48659 => -32730,
    48660 => -32731,
    48661 => -32731,
    48662 => -32731,
    48663 => -32731,
    48664 => -32731,
    48665 => -32731,
    48666 => -32731,
    48667 => -32732,
    48668 => -32732,
    48669 => -32732,
    48670 => -32732,
    48671 => -32732,
    48672 => -32732,
    48673 => -32732,
    48674 => -32733,
    48675 => -32733,
    48676 => -32733,
    48677 => -32733,
    48678 => -32733,
    48679 => -32733,
    48680 => -32733,
    48681 => -32734,
    48682 => -32734,
    48683 => -32734,
    48684 => -32734,
    48685 => -32734,
    48686 => -32734,
    48687 => -32734,
    48688 => -32735,
    48689 => -32735,
    48690 => -32735,
    48691 => -32735,
    48692 => -32735,
    48693 => -32735,
    48694 => -32735,
    48695 => -32736,
    48696 => -32736,
    48697 => -32736,
    48698 => -32736,
    48699 => -32736,
    48700 => -32736,
    48701 => -32736,
    48702 => -32737,
    48703 => -32737,
    48704 => -32737,
    48705 => -32737,
    48706 => -32737,
    48707 => -32737,
    48708 => -32737,
    48709 => -32737,
    48710 => -32738,
    48711 => -32738,
    48712 => -32738,
    48713 => -32738,
    48714 => -32738,
    48715 => -32738,
    48716 => -32738,
    48717 => -32739,
    48718 => -32739,
    48719 => -32739,
    48720 => -32739,
    48721 => -32739,
    48722 => -32739,
    48723 => -32739,
    48724 => -32739,
    48725 => -32740,
    48726 => -32740,
    48727 => -32740,
    48728 => -32740,
    48729 => -32740,
    48730 => -32740,
    48731 => -32740,
    48732 => -32740,
    48733 => -32741,
    48734 => -32741,
    48735 => -32741,
    48736 => -32741,
    48737 => -32741,
    48738 => -32741,
    48739 => -32741,
    48740 => -32741,
    48741 => -32742,
    48742 => -32742,
    48743 => -32742,
    48744 => -32742,
    48745 => -32742,
    48746 => -32742,
    48747 => -32742,
    48748 => -32742,
    48749 => -32743,
    48750 => -32743,
    48751 => -32743,
    48752 => -32743,
    48753 => -32743,
    48754 => -32743,
    48755 => -32743,
    48756 => -32743,
    48757 => -32744,
    48758 => -32744,
    48759 => -32744,
    48760 => -32744,
    48761 => -32744,
    48762 => -32744,
    48763 => -32744,
    48764 => -32744,
    48765 => -32744,
    48766 => -32745,
    48767 => -32745,
    48768 => -32745,
    48769 => -32745,
    48770 => -32745,
    48771 => -32745,
    48772 => -32745,
    48773 => -32745,
    48774 => -32745,
    48775 => -32746,
    48776 => -32746,
    48777 => -32746,
    48778 => -32746,
    48779 => -32746,
    48780 => -32746,
    48781 => -32746,
    48782 => -32746,
    48783 => -32746,
    48784 => -32747,
    48785 => -32747,
    48786 => -32747,
    48787 => -32747,
    48788 => -32747,
    48789 => -32747,
    48790 => -32747,
    48791 => -32747,
    48792 => -32747,
    48793 => -32748,
    48794 => -32748,
    48795 => -32748,
    48796 => -32748,
    48797 => -32748,
    48798 => -32748,
    48799 => -32748,
    48800 => -32748,
    48801 => -32748,
    48802 => -32749,
    48803 => -32749,
    48804 => -32749,
    48805 => -32749,
    48806 => -32749,
    48807 => -32749,
    48808 => -32749,
    48809 => -32749,
    48810 => -32749,
    48811 => -32749,
    48812 => -32750,
    48813 => -32750,
    48814 => -32750,
    48815 => -32750,
    48816 => -32750,
    48817 => -32750,
    48818 => -32750,
    48819 => -32750,
    48820 => -32750,
    48821 => -32751,
    48822 => -32751,
    48823 => -32751,
    48824 => -32751,
    48825 => -32751,
    48826 => -32751,
    48827 => -32751,
    48828 => -32751,
    48829 => -32751,
    48830 => -32751,
    48831 => -32751,
    48832 => -32752,
    48833 => -32752,
    48834 => -32752,
    48835 => -32752,
    48836 => -32752,
    48837 => -32752,
    48838 => -32752,
    48839 => -32752,
    48840 => -32752,
    48841 => -32752,
    48842 => -32753,
    48843 => -32753,
    48844 => -32753,
    48845 => -32753,
    48846 => -32753,
    48847 => -32753,
    48848 => -32753,
    48849 => -32753,
    48850 => -32753,
    48851 => -32753,
    48852 => -32753,
    48853 => -32754,
    48854 => -32754,
    48855 => -32754,
    48856 => -32754,
    48857 => -32754,
    48858 => -32754,
    48859 => -32754,
    48860 => -32754,
    48861 => -32754,
    48862 => -32754,
    48863 => -32754,
    48864 => -32755,
    48865 => -32755,
    48866 => -32755,
    48867 => -32755,
    48868 => -32755,
    48869 => -32755,
    48870 => -32755,
    48871 => -32755,
    48872 => -32755,
    48873 => -32755,
    48874 => -32755,
    48875 => -32755,
    48876 => -32756,
    48877 => -32756,
    48878 => -32756,
    48879 => -32756,
    48880 => -32756,
    48881 => -32756,
    48882 => -32756,
    48883 => -32756,
    48884 => -32756,
    48885 => -32756,
    48886 => -32756,
    48887 => -32756,
    48888 => -32757,
    48889 => -32757,
    48890 => -32757,
    48891 => -32757,
    48892 => -32757,
    48893 => -32757,
    48894 => -32757,
    48895 => -32757,
    48896 => -32757,
    48897 => -32757,
    48898 => -32757,
    48899 => -32757,
    48900 => -32757,
    48901 => -32758,
    48902 => -32758,
    48903 => -32758,
    48904 => -32758,
    48905 => -32758,
    48906 => -32758,
    48907 => -32758,
    48908 => -32758,
    48909 => -32758,
    48910 => -32758,
    48911 => -32758,
    48912 => -32758,
    48913 => -32758,
    48914 => -32758,
    48915 => -32759,
    48916 => -32759,
    48917 => -32759,
    48918 => -32759,
    48919 => -32759,
    48920 => -32759,
    48921 => -32759,
    48922 => -32759,
    48923 => -32759,
    48924 => -32759,
    48925 => -32759,
    48926 => -32759,
    48927 => -32759,
    48928 => -32759,
    48929 => -32760,
    48930 => -32760,
    48931 => -32760,
    48932 => -32760,
    48933 => -32760,
    48934 => -32760,
    48935 => -32760,
    48936 => -32760,
    48937 => -32760,
    48938 => -32760,
    48939 => -32760,
    48940 => -32760,
    48941 => -32760,
    48942 => -32760,
    48943 => -32760,
    48944 => -32760,
    48945 => -32761,
    48946 => -32761,
    48947 => -32761,
    48948 => -32761,
    48949 => -32761,
    48950 => -32761,
    48951 => -32761,
    48952 => -32761,
    48953 => -32761,
    48954 => -32761,
    48955 => -32761,
    48956 => -32761,
    48957 => -32761,
    48958 => -32761,
    48959 => -32761,
    48960 => -32761,
    48961 => -32762,
    48962 => -32762,
    48963 => -32762,
    48964 => -32762,
    48965 => -32762,
    48966 => -32762,
    48967 => -32762,
    48968 => -32762,
    48969 => -32762,
    48970 => -32762,
    48971 => -32762,
    48972 => -32762,
    48973 => -32762,
    48974 => -32762,
    48975 => -32762,
    48976 => -32762,
    48977 => -32762,
    48978 => -32762,
    48979 => -32762,
    48980 => -32763,
    48981 => -32763,
    48982 => -32763,
    48983 => -32763,
    48984 => -32763,
    48985 => -32763,
    48986 => -32763,
    48987 => -32763,
    48988 => -32763,
    48989 => -32763,
    48990 => -32763,
    48991 => -32763,
    48992 => -32763,
    48993 => -32763,
    48994 => -32763,
    48995 => -32763,
    48996 => -32763,
    48997 => -32763,
    48998 => -32763,
    48999 => -32763,
    49000 => -32764,
    49001 => -32764,
    49002 => -32764,
    49003 => -32764,
    49004 => -32764,
    49005 => -32764,
    49006 => -32764,
    49007 => -32764,
    49008 => -32764,
    49009 => -32764,
    49010 => -32764,
    49011 => -32764,
    49012 => -32764,
    49013 => -32764,
    49014 => -32764,
    49015 => -32764,
    49016 => -32764,
    49017 => -32764,
    49018 => -32764,
    49019 => -32764,
    49020 => -32764,
    49021 => -32764,
    49022 => -32764,
    49023 => -32764,
    49024 => -32765,
    49025 => -32765,
    49026 => -32765,
    49027 => -32765,
    49028 => -32765,
    49029 => -32765,
    49030 => -32765,
    49031 => -32765,
    49032 => -32765,
    49033 => -32765,
    49034 => -32765,
    49035 => -32765,
    49036 => -32765,
    49037 => -32765,
    49038 => -32765,
    49039 => -32765,
    49040 => -32765,
    49041 => -32765,
    49042 => -32765,
    49043 => -32765,
    49044 => -32765,
    49045 => -32765,
    49046 => -32765,
    49047 => -32765,
    49048 => -32765,
    49049 => -32765,
    49050 => -32765,
    49051 => -32765,
    49052 => -32765,
    49053 => -32766,
    49054 => -32766,
    49055 => -32766,
    49056 => -32766,
    49057 => -32766,
    49058 => -32766,
    49059 => -32766,
    49060 => -32766,
    49061 => -32766,
    49062 => -32766,
    49063 => -32766,
    49064 => -32766,
    49065 => -32766,
    49066 => -32766,
    49067 => -32766,
    49068 => -32766,
    49069 => -32766,
    49070 => -32766,
    49071 => -32766,
    49072 => -32766,
    49073 => -32766,
    49074 => -32766,
    49075 => -32766,
    49076 => -32766,
    49077 => -32766,
    49078 => -32766,
    49079 => -32766,
    49080 => -32766,
    49081 => -32766,
    49082 => -32766,
    49083 => -32766,
    49084 => -32766,
    49085 => -32766,
    49086 => -32766,
    49087 => -32766,
    49088 => -32766,
    49089 => -32766,
    49090 => -32766,
    49091 => -32766,
    49092 => -32766,
    49093 => -32766,
    49094 => -32766,
    49095 => -32767,
    49096 => -32767,
    49097 => -32767,
    49098 => -32767,
    49099 => -32767,
    49100 => -32767,
    49101 => -32767,
    49102 => -32767,
    49103 => -32767,
    49104 => -32767,
    49105 => -32767,
    49106 => -32767,
    49107 => -32767,
    49108 => -32767,
    49109 => -32767,
    49110 => -32767,
    49111 => -32767,
    49112 => -32767,
    49113 => -32767,
    49114 => -32767,
    49115 => -32767,
    49116 => -32767,
    49117 => -32767,
    49118 => -32767,
    49119 => -32767,
    49120 => -32767,
    49121 => -32767,
    49122 => -32767,
    49123 => -32767,
    49124 => -32767,
    49125 => -32767,
    49126 => -32767,
    49127 => -32767,
    49128 => -32767,
    49129 => -32767,
    49130 => -32767,
    49131 => -32767,
    49132 => -32767,
    49133 => -32767,
    49134 => -32767,
    49135 => -32767,
    49136 => -32767,
    49137 => -32767,
    49138 => -32767,
    49139 => -32767,
    49140 => -32767,
    49141 => -32767,
    49142 => -32767,
    49143 => -32767,
    49144 => -32767,
    49145 => -32767,
    49146 => -32767,
    49147 => -32767,
    49148 => -32767,
    49149 => -32767,
    49150 => -32767,
    49151 => -32767,
    49152 => -32767,
    49153 => -32767,
    49154 => -32767,
    49155 => -32767,
    49156 => -32767,
    49157 => -32767,
    49158 => -32767,
    49159 => -32767,
    49160 => -32767,
    49161 => -32767,
    49162 => -32767,
    49163 => -32767,
    49164 => -32767,
    49165 => -32767,
    49166 => -32767,
    49167 => -32767,
    49168 => -32767,
    49169 => -32767,
    49170 => -32767,
    49171 => -32767,
    49172 => -32767,
    49173 => -32767,
    49174 => -32767,
    49175 => -32767,
    49176 => -32767,
    49177 => -32767,
    49178 => -32767,
    49179 => -32767,
    49180 => -32767,
    49181 => -32767,
    49182 => -32767,
    49183 => -32767,
    49184 => -32767,
    49185 => -32767,
    49186 => -32767,
    49187 => -32767,
    49188 => -32767,
    49189 => -32767,
    49190 => -32767,
    49191 => -32767,
    49192 => -32767,
    49193 => -32767,
    49194 => -32767,
    49195 => -32767,
    49196 => -32767,
    49197 => -32767,
    49198 => -32767,
    49199 => -32767,
    49200 => -32767,
    49201 => -32767,
    49202 => -32767,
    49203 => -32767,
    49204 => -32767,
    49205 => -32767,
    49206 => -32767,
    49207 => -32767,
    49208 => -32767,
    49209 => -32767,
    49210 => -32766,
    49211 => -32766,
    49212 => -32766,
    49213 => -32766,
    49214 => -32766,
    49215 => -32766,
    49216 => -32766,
    49217 => -32766,
    49218 => -32766,
    49219 => -32766,
    49220 => -32766,
    49221 => -32766,
    49222 => -32766,
    49223 => -32766,
    49224 => -32766,
    49225 => -32766,
    49226 => -32766,
    49227 => -32766,
    49228 => -32766,
    49229 => -32766,
    49230 => -32766,
    49231 => -32766,
    49232 => -32766,
    49233 => -32766,
    49234 => -32766,
    49235 => -32766,
    49236 => -32766,
    49237 => -32766,
    49238 => -32766,
    49239 => -32766,
    49240 => -32766,
    49241 => -32766,
    49242 => -32766,
    49243 => -32766,
    49244 => -32766,
    49245 => -32766,
    49246 => -32766,
    49247 => -32766,
    49248 => -32766,
    49249 => -32766,
    49250 => -32766,
    49251 => -32766,
    49252 => -32765,
    49253 => -32765,
    49254 => -32765,
    49255 => -32765,
    49256 => -32765,
    49257 => -32765,
    49258 => -32765,
    49259 => -32765,
    49260 => -32765,
    49261 => -32765,
    49262 => -32765,
    49263 => -32765,
    49264 => -32765,
    49265 => -32765,
    49266 => -32765,
    49267 => -32765,
    49268 => -32765,
    49269 => -32765,
    49270 => -32765,
    49271 => -32765,
    49272 => -32765,
    49273 => -32765,
    49274 => -32765,
    49275 => -32765,
    49276 => -32765,
    49277 => -32765,
    49278 => -32765,
    49279 => -32765,
    49280 => -32765,
    49281 => -32764,
    49282 => -32764,
    49283 => -32764,
    49284 => -32764,
    49285 => -32764,
    49286 => -32764,
    49287 => -32764,
    49288 => -32764,
    49289 => -32764,
    49290 => -32764,
    49291 => -32764,
    49292 => -32764,
    49293 => -32764,
    49294 => -32764,
    49295 => -32764,
    49296 => -32764,
    49297 => -32764,
    49298 => -32764,
    49299 => -32764,
    49300 => -32764,
    49301 => -32764,
    49302 => -32764,
    49303 => -32764,
    49304 => -32764,
    49305 => -32763,
    49306 => -32763,
    49307 => -32763,
    49308 => -32763,
    49309 => -32763,
    49310 => -32763,
    49311 => -32763,
    49312 => -32763,
    49313 => -32763,
    49314 => -32763,
    49315 => -32763,
    49316 => -32763,
    49317 => -32763,
    49318 => -32763,
    49319 => -32763,
    49320 => -32763,
    49321 => -32763,
    49322 => -32763,
    49323 => -32763,
    49324 => -32763,
    49325 => -32762,
    49326 => -32762,
    49327 => -32762,
    49328 => -32762,
    49329 => -32762,
    49330 => -32762,
    49331 => -32762,
    49332 => -32762,
    49333 => -32762,
    49334 => -32762,
    49335 => -32762,
    49336 => -32762,
    49337 => -32762,
    49338 => -32762,
    49339 => -32762,
    49340 => -32762,
    49341 => -32762,
    49342 => -32762,
    49343 => -32762,
    49344 => -32761,
    49345 => -32761,
    49346 => -32761,
    49347 => -32761,
    49348 => -32761,
    49349 => -32761,
    49350 => -32761,
    49351 => -32761,
    49352 => -32761,
    49353 => -32761,
    49354 => -32761,
    49355 => -32761,
    49356 => -32761,
    49357 => -32761,
    49358 => -32761,
    49359 => -32761,
    49360 => -32760,
    49361 => -32760,
    49362 => -32760,
    49363 => -32760,
    49364 => -32760,
    49365 => -32760,
    49366 => -32760,
    49367 => -32760,
    49368 => -32760,
    49369 => -32760,
    49370 => -32760,
    49371 => -32760,
    49372 => -32760,
    49373 => -32760,
    49374 => -32760,
    49375 => -32760,
    49376 => -32759,
    49377 => -32759,
    49378 => -32759,
    49379 => -32759,
    49380 => -32759,
    49381 => -32759,
    49382 => -32759,
    49383 => -32759,
    49384 => -32759,
    49385 => -32759,
    49386 => -32759,
    49387 => -32759,
    49388 => -32759,
    49389 => -32759,
    49390 => -32758,
    49391 => -32758,
    49392 => -32758,
    49393 => -32758,
    49394 => -32758,
    49395 => -32758,
    49396 => -32758,
    49397 => -32758,
    49398 => -32758,
    49399 => -32758,
    49400 => -32758,
    49401 => -32758,
    49402 => -32758,
    49403 => -32758,
    49404 => -32757,
    49405 => -32757,
    49406 => -32757,
    49407 => -32757,
    49408 => -32757,
    49409 => -32757,
    49410 => -32757,
    49411 => -32757,
    49412 => -32757,
    49413 => -32757,
    49414 => -32757,
    49415 => -32757,
    49416 => -32757,
    49417 => -32756,
    49418 => -32756,
    49419 => -32756,
    49420 => -32756,
    49421 => -32756,
    49422 => -32756,
    49423 => -32756,
    49424 => -32756,
    49425 => -32756,
    49426 => -32756,
    49427 => -32756,
    49428 => -32756,
    49429 => -32755,
    49430 => -32755,
    49431 => -32755,
    49432 => -32755,
    49433 => -32755,
    49434 => -32755,
    49435 => -32755,
    49436 => -32755,
    49437 => -32755,
    49438 => -32755,
    49439 => -32755,
    49440 => -32755,
    49441 => -32754,
    49442 => -32754,
    49443 => -32754,
    49444 => -32754,
    49445 => -32754,
    49446 => -32754,
    49447 => -32754,
    49448 => -32754,
    49449 => -32754,
    49450 => -32754,
    49451 => -32754,
    49452 => -32753,
    49453 => -32753,
    49454 => -32753,
    49455 => -32753,
    49456 => -32753,
    49457 => -32753,
    49458 => -32753,
    49459 => -32753,
    49460 => -32753,
    49461 => -32753,
    49462 => -32753,
    49463 => -32752,
    49464 => -32752,
    49465 => -32752,
    49466 => -32752,
    49467 => -32752,
    49468 => -32752,
    49469 => -32752,
    49470 => -32752,
    49471 => -32752,
    49472 => -32752,
    49473 => -32751,
    49474 => -32751,
    49475 => -32751,
    49476 => -32751,
    49477 => -32751,
    49478 => -32751,
    49479 => -32751,
    49480 => -32751,
    49481 => -32751,
    49482 => -32751,
    49483 => -32751,
    49484 => -32750,
    49485 => -32750,
    49486 => -32750,
    49487 => -32750,
    49488 => -32750,
    49489 => -32750,
    49490 => -32750,
    49491 => -32750,
    49492 => -32750,
    49493 => -32749,
    49494 => -32749,
    49495 => -32749,
    49496 => -32749,
    49497 => -32749,
    49498 => -32749,
    49499 => -32749,
    49500 => -32749,
    49501 => -32749,
    49502 => -32749,
    49503 => -32748,
    49504 => -32748,
    49505 => -32748,
    49506 => -32748,
    49507 => -32748,
    49508 => -32748,
    49509 => -32748,
    49510 => -32748,
    49511 => -32748,
    49512 => -32747,
    49513 => -32747,
    49514 => -32747,
    49515 => -32747,
    49516 => -32747,
    49517 => -32747,
    49518 => -32747,
    49519 => -32747,
    49520 => -32747,
    49521 => -32746,
    49522 => -32746,
    49523 => -32746,
    49524 => -32746,
    49525 => -32746,
    49526 => -32746,
    49527 => -32746,
    49528 => -32746,
    49529 => -32746,
    49530 => -32745,
    49531 => -32745,
    49532 => -32745,
    49533 => -32745,
    49534 => -32745,
    49535 => -32745,
    49536 => -32745,
    49537 => -32745,
    49538 => -32745,
    49539 => -32744,
    49540 => -32744,
    49541 => -32744,
    49542 => -32744,
    49543 => -32744,
    49544 => -32744,
    49545 => -32744,
    49546 => -32744,
    49547 => -32744,
    49548 => -32743,
    49549 => -32743,
    49550 => -32743,
    49551 => -32743,
    49552 => -32743,
    49553 => -32743,
    49554 => -32743,
    49555 => -32743,
    49556 => -32742,
    49557 => -32742,
    49558 => -32742,
    49559 => -32742,
    49560 => -32742,
    49561 => -32742,
    49562 => -32742,
    49563 => -32742,
    49564 => -32741,
    49565 => -32741,
    49566 => -32741,
    49567 => -32741,
    49568 => -32741,
    49569 => -32741,
    49570 => -32741,
    49571 => -32741,
    49572 => -32740,
    49573 => -32740,
    49574 => -32740,
    49575 => -32740,
    49576 => -32740,
    49577 => -32740,
    49578 => -32740,
    49579 => -32740,
    49580 => -32739,
    49581 => -32739,
    49582 => -32739,
    49583 => -32739,
    49584 => -32739,
    49585 => -32739,
    49586 => -32739,
    49587 => -32739,
    49588 => -32738,
    49589 => -32738,
    49590 => -32738,
    49591 => -32738,
    49592 => -32738,
    49593 => -32738,
    49594 => -32738,
    49595 => -32737,
    49596 => -32737,
    49597 => -32737,
    49598 => -32737,
    49599 => -32737,
    49600 => -32737,
    49601 => -32737,
    49602 => -32737,
    49603 => -32736,
    49604 => -32736,
    49605 => -32736,
    49606 => -32736,
    49607 => -32736,
    49608 => -32736,
    49609 => -32736,
    49610 => -32735,
    49611 => -32735,
    49612 => -32735,
    49613 => -32735,
    49614 => -32735,
    49615 => -32735,
    49616 => -32735,
    49617 => -32734,
    49618 => -32734,
    49619 => -32734,
    49620 => -32734,
    49621 => -32734,
    49622 => -32734,
    49623 => -32734,
    49624 => -32733,
    49625 => -32733,
    49626 => -32733,
    49627 => -32733,
    49628 => -32733,
    49629 => -32733,
    49630 => -32733,
    49631 => -32732,
    49632 => -32732,
    49633 => -32732,
    49634 => -32732,
    49635 => -32732,
    49636 => -32732,
    49637 => -32732,
    49638 => -32731,
    49639 => -32731,
    49640 => -32731,
    49641 => -32731,
    49642 => -32731,
    49643 => -32731,
    49644 => -32731,
    49645 => -32730,
    49646 => -32730,
    49647 => -32730,
    49648 => -32730,
    49649 => -32730,
    49650 => -32730,
    49651 => -32730,
    49652 => -32729,
    49653 => -32729,
    49654 => -32729,
    49655 => -32729,
    49656 => -32729,
    49657 => -32729,
    49658 => -32728,
    49659 => -32728,
    49660 => -32728,
    49661 => -32728,
    49662 => -32728,
    49663 => -32728,
    49664 => -32728,
    49665 => -32727,
    49666 => -32727,
    49667 => -32727,
    49668 => -32727,
    49669 => -32727,
    49670 => -32727,
    49671 => -32726,
    49672 => -32726,
    49673 => -32726,
    49674 => -32726,
    49675 => -32726,
    49676 => -32726,
    49677 => -32726,
    49678 => -32725,
    49679 => -32725,
    49680 => -32725,
    49681 => -32725,
    49682 => -32725,
    49683 => -32725,
    49684 => -32724,
    49685 => -32724,
    49686 => -32724,
    49687 => -32724,
    49688 => -32724,
    49689 => -32724,
    49690 => -32723,
    49691 => -32723,
    49692 => -32723,
    49693 => -32723,
    49694 => -32723,
    49695 => -32723,
    49696 => -32722,
    49697 => -32722,
    49698 => -32722,
    49699 => -32722,
    49700 => -32722,
    49701 => -32722,
    49702 => -32721,
    49703 => -32721,
    49704 => -32721,
    49705 => -32721,
    49706 => -32721,
    49707 => -32721,
    49708 => -32720,
    49709 => -32720,
    49710 => -32720,
    49711 => -32720,
    49712 => -32720,
    49713 => -32720,
    49714 => -32719,
    49715 => -32719,
    49716 => -32719,
    49717 => -32719,
    49718 => -32719,
    49719 => -32719,
    49720 => -32718,
    49721 => -32718,
    49722 => -32718,
    49723 => -32718,
    49724 => -32718,
    49725 => -32718,
    49726 => -32717,
    49727 => -32717,
    49728 => -32717,
    49729 => -32717,
    49730 => -32717,
    49731 => -32717,
    49732 => -32716,
    49733 => -32716,
    49734 => -32716,
    49735 => -32716,
    49736 => -32716,
    49737 => -32715,
    49738 => -32715,
    49739 => -32715,
    49740 => -32715,
    49741 => -32715,
    49742 => -32715,
    49743 => -32714,
    49744 => -32714,
    49745 => -32714,
    49746 => -32714,
    49747 => -32714,
    49748 => -32714,
    49749 => -32713,
    49750 => -32713,
    49751 => -32713,
    49752 => -32713,
    49753 => -32713,
    49754 => -32712,
    49755 => -32712,
    49756 => -32712,
    49757 => -32712,
    49758 => -32712,
    49759 => -32712,
    49760 => -32711,
    49761 => -32711,
    49762 => -32711,
    49763 => -32711,
    49764 => -32711,
    49765 => -32710,
    49766 => -32710,
    49767 => -32710,
    49768 => -32710,
    49769 => -32710,
    49770 => -32710,
    49771 => -32709,
    49772 => -32709,
    49773 => -32709,
    49774 => -32709,
    49775 => -32709,
    49776 => -32708,
    49777 => -32708,
    49778 => -32708,
    49779 => -32708,
    49780 => -32708,
    49781 => -32707,
    49782 => -32707,
    49783 => -32707,
    49784 => -32707,
    49785 => -32707,
    49786 => -32706,
    49787 => -32706,
    49788 => -32706,
    49789 => -32706,
    49790 => -32706,
    49791 => -32706,
    49792 => -32705,
    49793 => -32705,
    49794 => -32705,
    49795 => -32705,
    49796 => -32705,
    49797 => -32704,
    49798 => -32704,
    49799 => -32704,
    49800 => -32704,
    49801 => -32704,
    49802 => -32703,
    49803 => -32703,
    49804 => -32703,
    49805 => -32703,
    49806 => -32703,
    49807 => -32702,
    49808 => -32702,
    49809 => -32702,
    49810 => -32702,
    49811 => -32702,
    49812 => -32701,
    49813 => -32701,
    49814 => -32701,
    49815 => -32701,
    49816 => -32701,
    49817 => -32700,
    49818 => -32700,
    49819 => -32700,
    49820 => -32700,
    49821 => -32700,
    49822 => -32699,
    49823 => -32699,
    49824 => -32699,
    49825 => -32699,
    49826 => -32699,
    49827 => -32698,
    49828 => -32698,
    49829 => -32698,
    49830 => -32698,
    49831 => -32698,
    49832 => -32697,
    49833 => -32697,
    49834 => -32697,
    49835 => -32697,
    49836 => -32697,
    49837 => -32696,
    49838 => -32696,
    49839 => -32696,
    49840 => -32696,
    49841 => -32696,
    49842 => -32695,
    49843 => -32695,
    49844 => -32695,
    49845 => -32695,
    49846 => -32694,
    49847 => -32694,
    49848 => -32694,
    49849 => -32694,
    49850 => -32694,
    49851 => -32693,
    49852 => -32693,
    49853 => -32693,
    49854 => -32693,
    49855 => -32693,
    49856 => -32692,
    49857 => -32692,
    49858 => -32692,
    49859 => -32692,
    49860 => -32692,
    49861 => -32691,
    49862 => -32691,
    49863 => -32691,
    49864 => -32691,
    49865 => -32690,
    49866 => -32690,
    49867 => -32690,
    49868 => -32690,
    49869 => -32690,
    49870 => -32689,
    49871 => -32689,
    49872 => -32689,
    49873 => -32689,
    49874 => -32689,
    49875 => -32688,
    49876 => -32688,
    49877 => -32688,
    49878 => -32688,
    49879 => -32687,
    49880 => -32687,
    49881 => -32687,
    49882 => -32687,
    49883 => -32687,
    49884 => -32686,
    49885 => -32686,
    49886 => -32686,
    49887 => -32686,
    49888 => -32685,
    49889 => -32685,
    49890 => -32685,
    49891 => -32685,
    49892 => -32685,
    49893 => -32684,
    49894 => -32684,
    49895 => -32684,
    49896 => -32684,
    49897 => -32683,
    49898 => -32683,
    49899 => -32683,
    49900 => -32683,
    49901 => -32683,
    49902 => -32682,
    49903 => -32682,
    49904 => -32682,
    49905 => -32682,
    49906 => -32681,
    49907 => -32681,
    49908 => -32681,
    49909 => -32681,
    49910 => -32681,
    49911 => -32680,
    49912 => -32680,
    49913 => -32680,
    49914 => -32680,
    49915 => -32679,
    49916 => -32679,
    49917 => -32679,
    49918 => -32679,
    49919 => -32678,
    49920 => -32678,
    49921 => -32678,
    49922 => -32678,
    49923 => -32678,
    49924 => -32677,
    49925 => -32677,
    49926 => -32677,
    49927 => -32677,
    49928 => -32676,
    49929 => -32676,
    49930 => -32676,
    49931 => -32676,
    49932 => -32675,
    49933 => -32675,
    49934 => -32675,
    49935 => -32675,
    49936 => -32674,
    49937 => -32674,
    49938 => -32674,
    49939 => -32674,
    49940 => -32674,
    49941 => -32673,
    49942 => -32673,
    49943 => -32673,
    49944 => -32673,
    49945 => -32672,
    49946 => -32672,
    49947 => -32672,
    49948 => -32672,
    49949 => -32671,
    49950 => -32671,
    49951 => -32671,
    49952 => -32671,
    49953 => -32670,
    49954 => -32670,
    49955 => -32670,
    49956 => -32670,
    49957 => -32669,
    49958 => -32669,
    49959 => -32669,
    49960 => -32669,
    49961 => -32668,
    49962 => -32668,
    49963 => -32668,
    49964 => -32668,
    49965 => -32668,
    49966 => -32667,
    49967 => -32667,
    49968 => -32667,
    49969 => -32667,
    49970 => -32666,
    49971 => -32666,
    49972 => -32666,
    49973 => -32666,
    49974 => -32665,
    49975 => -32665,
    49976 => -32665,
    49977 => -32665,
    49978 => -32664,
    49979 => -32664,
    49980 => -32664,
    49981 => -32664,
    49982 => -32663,
    49983 => -32663,
    49984 => -32663,
    49985 => -32663,
    49986 => -32662,
    49987 => -32662,
    49988 => -32662,
    49989 => -32662,
    49990 => -32661,
    49991 => -32661,
    49992 => -32661,
    49993 => -32661,
    49994 => -32660,
    49995 => -32660,
    49996 => -32660,
    49997 => -32660,
    49998 => -32659,
    49999 => -32659,
    50000 => -32659,
    50001 => -32659,
    50002 => -32658,
    50003 => -32658,
    50004 => -32658,
    50005 => -32657,
    50006 => -32657,
    50007 => -32657,
    50008 => -32657,
    50009 => -32656,
    50010 => -32656,
    50011 => -32656,
    50012 => -32656,
    50013 => -32655,
    50014 => -32655,
    50015 => -32655,
    50016 => -32655,
    50017 => -32654,
    50018 => -32654,
    50019 => -32654,
    50020 => -32654,
    50021 => -32653,
    50022 => -32653,
    50023 => -32653,
    50024 => -32653,
    50025 => -32652,
    50026 => -32652,
    50027 => -32652,
    50028 => -32652,
    50029 => -32651,
    50030 => -32651,
    50031 => -32651,
    50032 => -32650,
    50033 => -32650,
    50034 => -32650,
    50035 => -32650,
    50036 => -32649,
    50037 => -32649,
    50038 => -32649,
    50039 => -32649,
    50040 => -32648,
    50041 => -32648,
    50042 => -32648,
    50043 => -32648,
    50044 => -32647,
    50045 => -32647,
    50046 => -32647,
    50047 => -32646,
    50048 => -32646,
    50049 => -32646,
    50050 => -32646,
    50051 => -32645,
    50052 => -32645,
    50053 => -32645,
    50054 => -32645,
    50055 => -32644,
    50056 => -32644,
    50057 => -32644,
    50058 => -32643,
    50059 => -32643,
    50060 => -32643,
    50061 => -32643,
    50062 => -32642,
    50063 => -32642,
    50064 => -32642,
    50065 => -32642,
    50066 => -32641,
    50067 => -32641,
    50068 => -32641,
    50069 => -32640,
    50070 => -32640,
    50071 => -32640,
    50072 => -32640,
    50073 => -32639,
    50074 => -32639,
    50075 => -32639,
    50076 => -32639,
    50077 => -32638,
    50078 => -32638,
    50079 => -32638,
    50080 => -32637,
    50081 => -32637,
    50082 => -32637,
    50083 => -32637,
    50084 => -32636,
    50085 => -32636,
    50086 => -32636,
    50087 => -32635,
    50088 => -32635,
    50089 => -32635,
    50090 => -32635,
    50091 => -32634,
    50092 => -32634,
    50093 => -32634,
    50094 => -32633,
    50095 => -32633,
    50096 => -32633,
    50097 => -32633,
    50098 => -32632,
    50099 => -32632,
    50100 => -32632,
    50101 => -32631,
    50102 => -32631,
    50103 => -32631,
    50104 => -32631,
    50105 => -32630,
    50106 => -32630,
    50107 => -32630,
    50108 => -32629,
    50109 => -32629,
    50110 => -32629,
    50111 => -32629,
    50112 => -32628,
    50113 => -32628,
    50114 => -32628,
    50115 => -32627,
    50116 => -32627,
    50117 => -32627,
    50118 => -32627,
    50119 => -32626,
    50120 => -32626,
    50121 => -32626,
    50122 => -32625,
    50123 => -32625,
    50124 => -32625,
    50125 => -32625,
    50126 => -32624,
    50127 => -32624,
    50128 => -32624,
    50129 => -32623,
    50130 => -32623,
    50131 => -32623,
    50132 => -32622,
    50133 => -32622,
    50134 => -32622,
    50135 => -32622,
    50136 => -32621,
    50137 => -32621,
    50138 => -32621,
    50139 => -32620,
    50140 => -32620,
    50141 => -32620,
    50142 => -32620,
    50143 => -32619,
    50144 => -32619,
    50145 => -32619,
    50146 => -32618,
    50147 => -32618,
    50148 => -32618,
    50149 => -32617,
    50150 => -32617,
    50151 => -32617,
    50152 => -32617,
    50153 => -32616,
    50154 => -32616,
    50155 => -32616,
    50156 => -32615,
    50157 => -32615,
    50158 => -32615,
    50159 => -32614,
    50160 => -32614,
    50161 => -32614,
    50162 => -32613,
    50163 => -32613,
    50164 => -32613,
    50165 => -32613,
    50166 => -32612,
    50167 => -32612,
    50168 => -32612,
    50169 => -32611,
    50170 => -32611,
    50171 => -32611,
    50172 => -32610,
    50173 => -32610,
    50174 => -32610,
    50175 => -32610,
    50176 => -32609,
    50177 => -32609,
    50178 => -32609,
    50179 => -32608,
    50180 => -32608,
    50181 => -32608,
    50182 => -32607,
    50183 => -32607,
    50184 => -32607,
    50185 => -32606,
    50186 => -32606,
    50187 => -32606,
    50188 => -32606,
    50189 => -32605,
    50190 => -32605,
    50191 => -32605,
    50192 => -32604,
    50193 => -32604,
    50194 => -32604,
    50195 => -32603,
    50196 => -32603,
    50197 => -32603,
    50198 => -32602,
    50199 => -32602,
    50200 => -32602,
    50201 => -32601,
    50202 => -32601,
    50203 => -32601,
    50204 => -32600,
    50205 => -32600,
    50206 => -32600,
    50207 => -32600,
    50208 => -32599,
    50209 => -32599,
    50210 => -32599,
    50211 => -32598,
    50212 => -32598,
    50213 => -32598,
    50214 => -32597,
    50215 => -32597,
    50216 => -32597,
    50217 => -32596,
    50218 => -32596,
    50219 => -32596,
    50220 => -32595,
    50221 => -32595,
    50222 => -32595,
    50223 => -32594,
    50224 => -32594,
    50225 => -32594,
    50226 => -32593,
    50227 => -32593,
    50228 => -32593,
    50229 => -32592,
    50230 => -32592,
    50231 => -32592,
    50232 => -32592,
    50233 => -32591,
    50234 => -32591,
    50235 => -32591,
    50236 => -32590,
    50237 => -32590,
    50238 => -32590,
    50239 => -32589,
    50240 => -32589,
    50241 => -32589,
    50242 => -32588,
    50243 => -32588,
    50244 => -32588,
    50245 => -32587,
    50246 => -32587,
    50247 => -32587,
    50248 => -32586,
    50249 => -32586,
    50250 => -32586,
    50251 => -32585,
    50252 => -32585,
    50253 => -32585,
    50254 => -32584,
    50255 => -32584,
    50256 => -32584,
    50257 => -32583,
    50258 => -32583,
    50259 => -32583,
    50260 => -32582,
    50261 => -32582,
    50262 => -32582,
    50263 => -32581,
    50264 => -32581,
    50265 => -32581,
    50266 => -32580,
    50267 => -32580,
    50268 => -32580,
    50269 => -32579,
    50270 => -32579,
    50271 => -32579,
    50272 => -32578,
    50273 => -32578,
    50274 => -32578,
    50275 => -32577,
    50276 => -32577,
    50277 => -32577,
    50278 => -32576,
    50279 => -32576,
    50280 => -32576,
    50281 => -32575,
    50282 => -32575,
    50283 => -32575,
    50284 => -32574,
    50285 => -32574,
    50286 => -32574,
    50287 => -32573,
    50288 => -32573,
    50289 => -32573,
    50290 => -32572,
    50291 => -32572,
    50292 => -32571,
    50293 => -32571,
    50294 => -32571,
    50295 => -32570,
    50296 => -32570,
    50297 => -32570,
    50298 => -32569,
    50299 => -32569,
    50300 => -32569,
    50301 => -32568,
    50302 => -32568,
    50303 => -32568,
    50304 => -32567,
    50305 => -32567,
    50306 => -32567,
    50307 => -32566,
    50308 => -32566,
    50309 => -32566,
    50310 => -32565,
    50311 => -32565,
    50312 => -32565,
    50313 => -32564,
    50314 => -32564,
    50315 => -32564,
    50316 => -32563,
    50317 => -32563,
    50318 => -32562,
    50319 => -32562,
    50320 => -32562,
    50321 => -32561,
    50322 => -32561,
    50323 => -32561,
    50324 => -32560,
    50325 => -32560,
    50326 => -32560,
    50327 => -32559,
    50328 => -32559,
    50329 => -32559,
    50330 => -32558,
    50331 => -32558,
    50332 => -32558,
    50333 => -32557,
    50334 => -32557,
    50335 => -32556,
    50336 => -32556,
    50337 => -32556,
    50338 => -32555,
    50339 => -32555,
    50340 => -32555,
    50341 => -32554,
    50342 => -32554,
    50343 => -32554,
    50344 => -32553,
    50345 => -32553,
    50346 => -32553,
    50347 => -32552,
    50348 => -32552,
    50349 => -32551,
    50350 => -32551,
    50351 => -32551,
    50352 => -32550,
    50353 => -32550,
    50354 => -32550,
    50355 => -32549,
    50356 => -32549,
    50357 => -32549,
    50358 => -32548,
    50359 => -32548,
    50360 => -32547,
    50361 => -32547,
    50362 => -32547,
    50363 => -32546,
    50364 => -32546,
    50365 => -32546,
    50366 => -32545,
    50367 => -32545,
    50368 => -32545,
    50369 => -32544,
    50370 => -32544,
    50371 => -32543,
    50372 => -32543,
    50373 => -32543,
    50374 => -32542,
    50375 => -32542,
    50376 => -32542,
    50377 => -32541,
    50378 => -32541,
    50379 => -32541,
    50380 => -32540,
    50381 => -32540,
    50382 => -32539,
    50383 => -32539,
    50384 => -32539,
    50385 => -32538,
    50386 => -32538,
    50387 => -32538,
    50388 => -32537,
    50389 => -32537,
    50390 => -32536,
    50391 => -32536,
    50392 => -32536,
    50393 => -32535,
    50394 => -32535,
    50395 => -32535,
    50396 => -32534,
    50397 => -32534,
    50398 => -32533,
    50399 => -32533,
    50400 => -32533,
    50401 => -32532,
    50402 => -32532,
    50403 => -32532,
    50404 => -32531,
    50405 => -32531,
    50406 => -32530,
    50407 => -32530,
    50408 => -32530,
    50409 => -32529,
    50410 => -32529,
    50411 => -32529,
    50412 => -32528,
    50413 => -32528,
    50414 => -32527,
    50415 => -32527,
    50416 => -32527,
    50417 => -32526,
    50418 => -32526,
    50419 => -32526,
    50420 => -32525,
    50421 => -32525,
    50422 => -32524,
    50423 => -32524,
    50424 => -32524,
    50425 => -32523,
    50426 => -32523,
    50427 => -32522,
    50428 => -32522,
    50429 => -32522,
    50430 => -32521,
    50431 => -32521,
    50432 => -32521,
    50433 => -32520,
    50434 => -32520,
    50435 => -32519,
    50436 => -32519,
    50437 => -32519,
    50438 => -32518,
    50439 => -32518,
    50440 => -32517,
    50441 => -32517,
    50442 => -32517,
    50443 => -32516,
    50444 => -32516,
    50445 => -32516,
    50446 => -32515,
    50447 => -32515,
    50448 => -32514,
    50449 => -32514,
    50450 => -32514,
    50451 => -32513,
    50452 => -32513,
    50453 => -32512,
    50454 => -32512,
    50455 => -32512,
    50456 => -32511,
    50457 => -32511,
    50458 => -32510,
    50459 => -32510,
    50460 => -32510,
    50461 => -32509,
    50462 => -32509,
    50463 => -32509,
    50464 => -32508,
    50465 => -32508,
    50466 => -32507,
    50467 => -32507,
    50468 => -32507,
    50469 => -32506,
    50470 => -32506,
    50471 => -32505,
    50472 => -32505,
    50473 => -32505,
    50474 => -32504,
    50475 => -32504,
    50476 => -32503,
    50477 => -32503,
    50478 => -32503,
    50479 => -32502,
    50480 => -32502,
    50481 => -32501,
    50482 => -32501,
    50483 => -32501,
    50484 => -32500,
    50485 => -32500,
    50486 => -32499,
    50487 => -32499,
    50488 => -32499,
    50489 => -32498,
    50490 => -32498,
    50491 => -32497,
    50492 => -32497,
    50493 => -32497,
    50494 => -32496,
    50495 => -32496,
    50496 => -32495,
    50497 => -32495,
    50498 => -32495,
    50499 => -32494,
    50500 => -32494,
    50501 => -32493,
    50502 => -32493,
    50503 => -32493,
    50504 => -32492,
    50505 => -32492,
    50506 => -32491,
    50507 => -32491,
    50508 => -32490,
    50509 => -32490,
    50510 => -32490,
    50511 => -32489,
    50512 => -32489,
    50513 => -32488,
    50514 => -32488,
    50515 => -32488,
    50516 => -32487,
    50517 => -32487,
    50518 => -32486,
    50519 => -32486,
    50520 => -32486,
    50521 => -32485,
    50522 => -32485,
    50523 => -32484,
    50524 => -32484,
    50525 => -32484,
    50526 => -32483,
    50527 => -32483,
    50528 => -32482,
    50529 => -32482,
    50530 => -32481,
    50531 => -32481,
    50532 => -32481,
    50533 => -32480,
    50534 => -32480,
    50535 => -32479,
    50536 => -32479,
    50537 => -32479,
    50538 => -32478,
    50539 => -32478,
    50540 => -32477,
    50541 => -32477,
    50542 => -32476,
    50543 => -32476,
    50544 => -32476,
    50545 => -32475,
    50546 => -32475,
    50547 => -32474,
    50548 => -32474,
    50549 => -32474,
    50550 => -32473,
    50551 => -32473,
    50552 => -32472,
    50553 => -32472,
    50554 => -32471,
    50555 => -32471,
    50556 => -32471,
    50557 => -32470,
    50558 => -32470,
    50559 => -32469,
    50560 => -32469,
    50561 => -32468,
    50562 => -32468,
    50563 => -32468,
    50564 => -32467,
    50565 => -32467,
    50566 => -32466,
    50567 => -32466,
    50568 => -32466,
    50569 => -32465,
    50570 => -32465,
    50571 => -32464,
    50572 => -32464,
    50573 => -32463,
    50574 => -32463,
    50575 => -32463,
    50576 => -32462,
    50577 => -32462,
    50578 => -32461,
    50579 => -32461,
    50580 => -32460,
    50581 => -32460,
    50582 => -32460,
    50583 => -32459,
    50584 => -32459,
    50585 => -32458,
    50586 => -32458,
    50587 => -32457,
    50588 => -32457,
    50589 => -32457,
    50590 => -32456,
    50591 => -32456,
    50592 => -32455,
    50593 => -32455,
    50594 => -32454,
    50595 => -32454,
    50596 => -32453,
    50597 => -32453,
    50598 => -32453,
    50599 => -32452,
    50600 => -32452,
    50601 => -32451,
    50602 => -32451,
    50603 => -32450,
    50604 => -32450,
    50605 => -32450,
    50606 => -32449,
    50607 => -32449,
    50608 => -32448,
    50609 => -32448,
    50610 => -32447,
    50611 => -32447,
    50612 => -32447,
    50613 => -32446,
    50614 => -32446,
    50615 => -32445,
    50616 => -32445,
    50617 => -32444,
    50618 => -32444,
    50619 => -32443,
    50620 => -32443,
    50621 => -32443,
    50622 => -32442,
    50623 => -32442,
    50624 => -32441,
    50625 => -32441,
    50626 => -32440,
    50627 => -32440,
    50628 => -32439,
    50629 => -32439,
    50630 => -32439,
    50631 => -32438,
    50632 => -32438,
    50633 => -32437,
    50634 => -32437,
    50635 => -32436,
    50636 => -32436,
    50637 => -32435,
    50638 => -32435,
    50639 => -32435,
    50640 => -32434,
    50641 => -32434,
    50642 => -32433,
    50643 => -32433,
    50644 => -32432,
    50645 => -32432,
    50646 => -32431,
    50647 => -32431,
    50648 => -32431,
    50649 => -32430,
    50650 => -32430,
    50651 => -32429,
    50652 => -32429,
    50653 => -32428,
    50654 => -32428,
    50655 => -32427,
    50656 => -32427,
    50657 => -32426,
    50658 => -32426,
    50659 => -32426,
    50660 => -32425,
    50661 => -32425,
    50662 => -32424,
    50663 => -32424,
    50664 => -32423,
    50665 => -32423,
    50666 => -32422,
    50667 => -32422,
    50668 => -32422,
    50669 => -32421,
    50670 => -32421,
    50671 => -32420,
    50672 => -32420,
    50673 => -32419,
    50674 => -32419,
    50675 => -32418,
    50676 => -32418,
    50677 => -32417,
    50678 => -32417,
    50679 => -32416,
    50680 => -32416,
    50681 => -32416,
    50682 => -32415,
    50683 => -32415,
    50684 => -32414,
    50685 => -32414,
    50686 => -32413,
    50687 => -32413,
    50688 => -32412,
    50689 => -32412,
    50690 => -32411,
    50691 => -32411,
    50692 => -32411,
    50693 => -32410,
    50694 => -32410,
    50695 => -32409,
    50696 => -32409,
    50697 => -32408,
    50698 => -32408,
    50699 => -32407,
    50700 => -32407,
    50701 => -32406,
    50702 => -32406,
    50703 => -32405,
    50704 => -32405,
    50705 => -32404,
    50706 => -32404,
    50707 => -32404,
    50708 => -32403,
    50709 => -32403,
    50710 => -32402,
    50711 => -32402,
    50712 => -32401,
    50713 => -32401,
    50714 => -32400,
    50715 => -32400,
    50716 => -32399,
    50717 => -32399,
    50718 => -32398,
    50719 => -32398,
    50720 => -32397,
    50721 => -32397,
    50722 => -32397,
    50723 => -32396,
    50724 => -32396,
    50725 => -32395,
    50726 => -32395,
    50727 => -32394,
    50728 => -32394,
    50729 => -32393,
    50730 => -32393,
    50731 => -32392,
    50732 => -32392,
    50733 => -32391,
    50734 => -32391,
    50735 => -32390,
    50736 => -32390,
    50737 => -32389,
    50738 => -32389,
    50739 => -32388,
    50740 => -32388,
    50741 => -32387,
    50742 => -32387,
    50743 => -32387,
    50744 => -32386,
    50745 => -32386,
    50746 => -32385,
    50747 => -32385,
    50748 => -32384,
    50749 => -32384,
    50750 => -32383,
    50751 => -32383,
    50752 => -32382,
    50753 => -32382,
    50754 => -32381,
    50755 => -32381,
    50756 => -32380,
    50757 => -32380,
    50758 => -32379,
    50759 => -32379,
    50760 => -32378,
    50761 => -32378,
    50762 => -32377,
    50763 => -32377,
    50764 => -32376,
    50765 => -32376,
    50766 => -32375,
    50767 => -32375,
    50768 => -32375,
    50769 => -32374,
    50770 => -32374,
    50771 => -32373,
    50772 => -32373,
    50773 => -32372,
    50774 => -32372,
    50775 => -32371,
    50776 => -32371,
    50777 => -32370,
    50778 => -32370,
    50779 => -32369,
    50780 => -32369,
    50781 => -32368,
    50782 => -32368,
    50783 => -32367,
    50784 => -32367,
    50785 => -32366,
    50786 => -32366,
    50787 => -32365,
    50788 => -32365,
    50789 => -32364,
    50790 => -32364,
    50791 => -32363,
    50792 => -32363,
    50793 => -32362,
    50794 => -32362,
    50795 => -32361,
    50796 => -32361,
    50797 => -32360,
    50798 => -32360,
    50799 => -32359,
    50800 => -32359,
    50801 => -32358,
    50802 => -32358,
    50803 => -32357,
    50804 => -32357,
    50805 => -32356,
    50806 => -32356,
    50807 => -32355,
    50808 => -32355,
    50809 => -32354,
    50810 => -32354,
    50811 => -32353,
    50812 => -32353,
    50813 => -32352,
    50814 => -32352,
    50815 => -32351,
    50816 => -32351,
    50817 => -32350,
    50818 => -32350,
    50819 => -32349,
    50820 => -32349,
    50821 => -32348,
    50822 => -32348,
    50823 => -32347,
    50824 => -32347,
    50825 => -32346,
    50826 => -32346,
    50827 => -32345,
    50828 => -32345,
    50829 => -32344,
    50830 => -32344,
    50831 => -32343,
    50832 => -32343,
    50833 => -32342,
    50834 => -32342,
    50835 => -32341,
    50836 => -32341,
    50837 => -32340,
    50838 => -32340,
    50839 => -32339,
    50840 => -32339,
    50841 => -32338,
    50842 => -32338,
    50843 => -32337,
    50844 => -32337,
    50845 => -32336,
    50846 => -32336,
    50847 => -32335,
    50848 => -32335,
    50849 => -32334,
    50850 => -32334,
    50851 => -32333,
    50852 => -32333,
    50853 => -32332,
    50854 => -32332,
    50855 => -32331,
    50856 => -32331,
    50857 => -32330,
    50858 => -32330,
    50859 => -32329,
    50860 => -32329,
    50861 => -32328,
    50862 => -32328,
    50863 => -32327,
    50864 => -32327,
    50865 => -32326,
    50866 => -32326,
    50867 => -32325,
    50868 => -32325,
    50869 => -32324,
    50870 => -32324,
    50871 => -32323,
    50872 => -32322,
    50873 => -32322,
    50874 => -32321,
    50875 => -32321,
    50876 => -32320,
    50877 => -32320,
    50878 => -32319,
    50879 => -32319,
    50880 => -32318,
    50881 => -32318,
    50882 => -32317,
    50883 => -32317,
    50884 => -32316,
    50885 => -32316,
    50886 => -32315,
    50887 => -32315,
    50888 => -32314,
    50889 => -32314,
    50890 => -32313,
    50891 => -32313,
    50892 => -32312,
    50893 => -32312,
    50894 => -32311,
    50895 => -32311,
    50896 => -32310,
    50897 => -32310,
    50898 => -32309,
    50899 => -32308,
    50900 => -32308,
    50901 => -32307,
    50902 => -32307,
    50903 => -32306,
    50904 => -32306,
    50905 => -32305,
    50906 => -32305,
    50907 => -32304,
    50908 => -32304,
    50909 => -32303,
    50910 => -32303,
    50911 => -32302,
    50912 => -32302,
    50913 => -32301,
    50914 => -32301,
    50915 => -32300,
    50916 => -32300,
    50917 => -32299,
    50918 => -32298,
    50919 => -32298,
    50920 => -32297,
    50921 => -32297,
    50922 => -32296,
    50923 => -32296,
    50924 => -32295,
    50925 => -32295,
    50926 => -32294,
    50927 => -32294,
    50928 => -32293,
    50929 => -32293,
    50930 => -32292,
    50931 => -32292,
    50932 => -32291,
    50933 => -32290,
    50934 => -32290,
    50935 => -32289,
    50936 => -32289,
    50937 => -32288,
    50938 => -32288,
    50939 => -32287,
    50940 => -32287,
    50941 => -32286,
    50942 => -32286,
    50943 => -32285,
    50944 => -32285,
    50945 => -32284,
    50946 => -32284,
    50947 => -32283,
    50948 => -32282,
    50949 => -32282,
    50950 => -32281,
    50951 => -32281,
    50952 => -32280,
    50953 => -32280,
    50954 => -32279,
    50955 => -32279,
    50956 => -32278,
    50957 => -32278,
    50958 => -32277,
    50959 => -32277,
    50960 => -32276,
    50961 => -32275,
    50962 => -32275,
    50963 => -32274,
    50964 => -32274,
    50965 => -32273,
    50966 => -32273,
    50967 => -32272,
    50968 => -32272,
    50969 => -32271,
    50970 => -32271,
    50971 => -32270,
    50972 => -32269,
    50973 => -32269,
    50974 => -32268,
    50975 => -32268,
    50976 => -32267,
    50977 => -32267,
    50978 => -32266,
    50979 => -32266,
    50980 => -32265,
    50981 => -32265,
    50982 => -32264,
    50983 => -32263,
    50984 => -32263,
    50985 => -32262,
    50986 => -32262,
    50987 => -32261,
    50988 => -32261,
    50989 => -32260,
    50990 => -32260,
    50991 => -32259,
    50992 => -32258,
    50993 => -32258,
    50994 => -32257,
    50995 => -32257,
    50996 => -32256,
    50997 => -32256,
    50998 => -32255,
    50999 => -32255,
    51000 => -32254,
    51001 => -32253,
    51002 => -32253,
    51003 => -32252,
    51004 => -32252,
    51005 => -32251,
    51006 => -32251,
    51007 => -32250,
    51008 => -32250,
    51009 => -32249,
    51010 => -32248,
    51011 => -32248,
    51012 => -32247,
    51013 => -32247,
    51014 => -32246,
    51015 => -32246,
    51016 => -32245,
    51017 => -32245,
    51018 => -32244,
    51019 => -32243,
    51020 => -32243,
    51021 => -32242,
    51022 => -32242,
    51023 => -32241,
    51024 => -32241,
    51025 => -32240,
    51026 => -32240,
    51027 => -32239,
    51028 => -32238,
    51029 => -32238,
    51030 => -32237,
    51031 => -32237,
    51032 => -32236,
    51033 => -32236,
    51034 => -32235,
    51035 => -32234,
    51036 => -32234,
    51037 => -32233,
    51038 => -32233,
    51039 => -32232,
    51040 => -32232,
    51041 => -32231,
    51042 => -32231,
    51043 => -32230,
    51044 => -32229,
    51045 => -32229,
    51046 => -32228,
    51047 => -32228,
    51048 => -32227,
    51049 => -32227,
    51050 => -32226,
    51051 => -32225,
    51052 => -32225,
    51053 => -32224,
    51054 => -32224,
    51055 => -32223,
    51056 => -32223,
    51057 => -32222,
    51058 => -32221,
    51059 => -32221,
    51060 => -32220,
    51061 => -32220,
    51062 => -32219,
    51063 => -32219,
    51064 => -32218,
    51065 => -32217,
    51066 => -32217,
    51067 => -32216,
    51068 => -32216,
    51069 => -32215,
    51070 => -32215,
    51071 => -32214,
    51072 => -32213,
    51073 => -32213,
    51074 => -32212,
    51075 => -32212,
    51076 => -32211,
    51077 => -32211,
    51078 => -32210,
    51079 => -32209,
    51080 => -32209,
    51081 => -32208,
    51082 => -32208,
    51083 => -32207,
    51084 => -32206,
    51085 => -32206,
    51086 => -32205,
    51087 => -32205,
    51088 => -32204,
    51089 => -32204,
    51090 => -32203,
    51091 => -32202,
    51092 => -32202,
    51093 => -32201,
    51094 => -32201,
    51095 => -32200,
    51096 => -32200,
    51097 => -32199,
    51098 => -32198,
    51099 => -32198,
    51100 => -32197,
    51101 => -32197,
    51102 => -32196,
    51103 => -32195,
    51104 => -32195,
    51105 => -32194,
    51106 => -32194,
    51107 => -32193,
    51108 => -32193,
    51109 => -32192,
    51110 => -32191,
    51111 => -32191,
    51112 => -32190,
    51113 => -32190,
    51114 => -32189,
    51115 => -32188,
    51116 => -32188,
    51117 => -32187,
    51118 => -32187,
    51119 => -32186,
    51120 => -32185,
    51121 => -32185,
    51122 => -32184,
    51123 => -32184,
    51124 => -32183,
    51125 => -32183,
    51126 => -32182,
    51127 => -32181,
    51128 => -32181,
    51129 => -32180,
    51130 => -32180,
    51131 => -32179,
    51132 => -32178,
    51133 => -32178,
    51134 => -32177,
    51135 => -32177,
    51136 => -32176,
    51137 => -32175,
    51138 => -32175,
    51139 => -32174,
    51140 => -32174,
    51141 => -32173,
    51142 => -32172,
    51143 => -32172,
    51144 => -32171,
    51145 => -32171,
    51146 => -32170,
    51147 => -32169,
    51148 => -32169,
    51149 => -32168,
    51150 => -32168,
    51151 => -32167,
    51152 => -32166,
    51153 => -32166,
    51154 => -32165,
    51155 => -32165,
    51156 => -32164,
    51157 => -32163,
    51158 => -32163,
    51159 => -32162,
    51160 => -32162,
    51161 => -32161,
    51162 => -32160,
    51163 => -32160,
    51164 => -32159,
    51165 => -32159,
    51166 => -32158,
    51167 => -32157,
    51168 => -32157,
    51169 => -32156,
    51170 => -32156,
    51171 => -32155,
    51172 => -32154,
    51173 => -32154,
    51174 => -32153,
    51175 => -32153,
    51176 => -32152,
    51177 => -32151,
    51178 => -32151,
    51179 => -32150,
    51180 => -32150,
    51181 => -32149,
    51182 => -32148,
    51183 => -32148,
    51184 => -32147,
    51185 => -32147,
    51186 => -32146,
    51187 => -32145,
    51188 => -32145,
    51189 => -32144,
    51190 => -32144,
    51191 => -32143,
    51192 => -32142,
    51193 => -32142,
    51194 => -32141,
    51195 => -32140,
    51196 => -32140,
    51197 => -32139,
    51198 => -32139,
    51199 => -32138,
    51200 => -32137,
    51201 => -32137,
    51202 => -32136,
    51203 => -32136,
    51204 => -32135,
    51205 => -32134,
    51206 => -32134,
    51207 => -32133,
    51208 => -32132,
    51209 => -32132,
    51210 => -32131,
    51211 => -32131,
    51212 => -32130,
    51213 => -32129,
    51214 => -32129,
    51215 => -32128,
    51216 => -32128,
    51217 => -32127,
    51218 => -32126,
    51219 => -32126,
    51220 => -32125,
    51221 => -32124,
    51222 => -32124,
    51223 => -32123,
    51224 => -32123,
    51225 => -32122,
    51226 => -32121,
    51227 => -32121,
    51228 => -32120,
    51229 => -32119,
    51230 => -32119,
    51231 => -32118,
    51232 => -32118,
    51233 => -32117,
    51234 => -32116,
    51235 => -32116,
    51236 => -32115,
    51237 => -32115,
    51238 => -32114,
    51239 => -32113,
    51240 => -32113,
    51241 => -32112,
    51242 => -32111,
    51243 => -32111,
    51244 => -32110,
    51245 => -32110,
    51246 => -32109,
    51247 => -32108,
    51248 => -32108,
    51249 => -32107,
    51250 => -32106,
    51251 => -32106,
    51252 => -32105,
    51253 => -32104,
    51254 => -32104,
    51255 => -32103,
    51256 => -32103,
    51257 => -32102,
    51258 => -32101,
    51259 => -32101,
    51260 => -32100,
    51261 => -32099,
    51262 => -32099,
    51263 => -32098,
    51264 => -32098,
    51265 => -32097,
    51266 => -32096,
    51267 => -32096,
    51268 => -32095,
    51269 => -32094,
    51270 => -32094,
    51271 => -32093,
    51272 => -32092,
    51273 => -32092,
    51274 => -32091,
    51275 => -32091,
    51276 => -32090,
    51277 => -32089,
    51278 => -32089,
    51279 => -32088,
    51280 => -32087,
    51281 => -32087,
    51282 => -32086,
    51283 => -32086,
    51284 => -32085,
    51285 => -32084,
    51286 => -32084,
    51287 => -32083,
    51288 => -32082,
    51289 => -32082,
    51290 => -32081,
    51291 => -32080,
    51292 => -32080,
    51293 => -32079,
    51294 => -32078,
    51295 => -32078,
    51296 => -32077,
    51297 => -32077,
    51298 => -32076,
    51299 => -32075,
    51300 => -32075,
    51301 => -32074,
    51302 => -32073,
    51303 => -32073,
    51304 => -32072,
    51305 => -32071,
    51306 => -32071,
    51307 => -32070,
    51308 => -32069,
    51309 => -32069,
    51310 => -32068,
    51311 => -32068,
    51312 => -32067,
    51313 => -32066,
    51314 => -32066,
    51315 => -32065,
    51316 => -32064,
    51317 => -32064,
    51318 => -32063,
    51319 => -32062,
    51320 => -32062,
    51321 => -32061,
    51322 => -32060,
    51323 => -32060,
    51324 => -32059,
    51325 => -32058,
    51326 => -32058,
    51327 => -32057,
    51328 => -32057,
    51329 => -32056,
    51330 => -32055,
    51331 => -32055,
    51332 => -32054,
    51333 => -32053,
    51334 => -32053,
    51335 => -32052,
    51336 => -32051,
    51337 => -32051,
    51338 => -32050,
    51339 => -32049,
    51340 => -32049,
    51341 => -32048,
    51342 => -32047,
    51343 => -32047,
    51344 => -32046,
    51345 => -32045,
    51346 => -32045,
    51347 => -32044,
    51348 => -32043,
    51349 => -32043,
    51350 => -32042,
    51351 => -32041,
    51352 => -32041,
    51353 => -32040,
    51354 => -32040,
    51355 => -32039,
    51356 => -32038,
    51357 => -32038,
    51358 => -32037,
    51359 => -32036,
    51360 => -32036,
    51361 => -32035,
    51362 => -32034,
    51363 => -32034,
    51364 => -32033,
    51365 => -32032,
    51366 => -32032,
    51367 => -32031,
    51368 => -32030,
    51369 => -32030,
    51370 => -32029,
    51371 => -32028,
    51372 => -32028,
    51373 => -32027,
    51374 => -32026,
    51375 => -32026,
    51376 => -32025,
    51377 => -32024,
    51378 => -32024,
    51379 => -32023,
    51380 => -32022,
    51381 => -32022,
    51382 => -32021,
    51383 => -32020,
    51384 => -32020,
    51385 => -32019,
    51386 => -32018,
    51387 => -32018,
    51388 => -32017,
    51389 => -32016,
    51390 => -32016,
    51391 => -32015,
    51392 => -32014,
    51393 => -32014,
    51394 => -32013,
    51395 => -32012,
    51396 => -32012,
    51397 => -32011,
    51398 => -32010,
    51399 => -32010,
    51400 => -32009,
    51401 => -32008,
    51402 => -32008,
    51403 => -32007,
    51404 => -32006,
    51405 => -32006,
    51406 => -32005,
    51407 => -32004,
    51408 => -32004,
    51409 => -32003,
    51410 => -32002,
    51411 => -32002,
    51412 => -32001,
    51413 => -32000,
    51414 => -31999,
    51415 => -31999,
    51416 => -31998,
    51417 => -31997,
    51418 => -31997,
    51419 => -31996,
    51420 => -31995,
    51421 => -31995,
    51422 => -31994,
    51423 => -31993,
    51424 => -31993,
    51425 => -31992,
    51426 => -31991,
    51427 => -31991,
    51428 => -31990,
    51429 => -31989,
    51430 => -31989,
    51431 => -31988,
    51432 => -31987,
    51433 => -31987,
    51434 => -31986,
    51435 => -31985,
    51436 => -31985,
    51437 => -31984,
    51438 => -31983,
    51439 => -31982,
    51440 => -31982,
    51441 => -31981,
    51442 => -31980,
    51443 => -31980,
    51444 => -31979,
    51445 => -31978,
    51446 => -31978,
    51447 => -31977,
    51448 => -31976,
    51449 => -31976,
    51450 => -31975,
    51451 => -31974,
    51452 => -31974,
    51453 => -31973,
    51454 => -31972,
    51455 => -31972,
    51456 => -31971,
    51457 => -31970,
    51458 => -31969,
    51459 => -31969,
    51460 => -31968,
    51461 => -31967,
    51462 => -31967,
    51463 => -31966,
    51464 => -31965,
    51465 => -31965,
    51466 => -31964,
    51467 => -31963,
    51468 => -31963,
    51469 => -31962,
    51470 => -31961,
    51471 => -31960,
    51472 => -31960,
    51473 => -31959,
    51474 => -31958,
    51475 => -31958,
    51476 => -31957,
    51477 => -31956,
    51478 => -31956,
    51479 => -31955,
    51480 => -31954,
    51481 => -31954,
    51482 => -31953,
    51483 => -31952,
    51484 => -31951,
    51485 => -31951,
    51486 => -31950,
    51487 => -31949,
    51488 => -31949,
    51489 => -31948,
    51490 => -31947,
    51491 => -31947,
    51492 => -31946,
    51493 => -31945,
    51494 => -31944,
    51495 => -31944,
    51496 => -31943,
    51497 => -31942,
    51498 => -31942,
    51499 => -31941,
    51500 => -31940,
    51501 => -31940,
    51502 => -31939,
    51503 => -31938,
    51504 => -31937,
    51505 => -31937,
    51506 => -31936,
    51507 => -31935,
    51508 => -31935,
    51509 => -31934,
    51510 => -31933,
    51511 => -31933,
    51512 => -31932,
    51513 => -31931,
    51514 => -31930,
    51515 => -31930,
    51516 => -31929,
    51517 => -31928,
    51518 => -31928,
    51519 => -31927,
    51520 => -31926,
    51521 => -31925,
    51522 => -31925,
    51523 => -31924,
    51524 => -31923,
    51525 => -31923,
    51526 => -31922,
    51527 => -31921,
    51528 => -31921,
    51529 => -31920,
    51530 => -31919,
    51531 => -31918,
    51532 => -31918,
    51533 => -31917,
    51534 => -31916,
    51535 => -31916,
    51536 => -31915,
    51537 => -31914,
    51538 => -31913,
    51539 => -31913,
    51540 => -31912,
    51541 => -31911,
    51542 => -31911,
    51543 => -31910,
    51544 => -31909,
    51545 => -31908,
    51546 => -31908,
    51547 => -31907,
    51548 => -31906,
    51549 => -31906,
    51550 => -31905,
    51551 => -31904,
    51552 => -31903,
    51553 => -31903,
    51554 => -31902,
    51555 => -31901,
    51556 => -31901,
    51557 => -31900,
    51558 => -31899,
    51559 => -31898,
    51560 => -31898,
    51561 => -31897,
    51562 => -31896,
    51563 => -31896,
    51564 => -31895,
    51565 => -31894,
    51566 => -31893,
    51567 => -31893,
    51568 => -31892,
    51569 => -31891,
    51570 => -31890,
    51571 => -31890,
    51572 => -31889,
    51573 => -31888,
    51574 => -31888,
    51575 => -31887,
    51576 => -31886,
    51577 => -31885,
    51578 => -31885,
    51579 => -31884,
    51580 => -31883,
    51581 => -31882,
    51582 => -31882,
    51583 => -31881,
    51584 => -31880,
    51585 => -31880,
    51586 => -31879,
    51587 => -31878,
    51588 => -31877,
    51589 => -31877,
    51590 => -31876,
    51591 => -31875,
    51592 => -31875,
    51593 => -31874,
    51594 => -31873,
    51595 => -31872,
    51596 => -31872,
    51597 => -31871,
    51598 => -31870,
    51599 => -31869,
    51600 => -31869,
    51601 => -31868,
    51602 => -31867,
    51603 => -31866,
    51604 => -31866,
    51605 => -31865,
    51606 => -31864,
    51607 => -31864,
    51608 => -31863,
    51609 => -31862,
    51610 => -31861,
    51611 => -31861,
    51612 => -31860,
    51613 => -31859,
    51614 => -31858,
    51615 => -31858,
    51616 => -31857,
    51617 => -31856,
    51618 => -31855,
    51619 => -31855,
    51620 => -31854,
    51621 => -31853,
    51622 => -31853,
    51623 => -31852,
    51624 => -31851,
    51625 => -31850,
    51626 => -31850,
    51627 => -31849,
    51628 => -31848,
    51629 => -31847,
    51630 => -31847,
    51631 => -31846,
    51632 => -31845,
    51633 => -31844,
    51634 => -31844,
    51635 => -31843,
    51636 => -31842,
    51637 => -31841,
    51638 => -31841,
    51639 => -31840,
    51640 => -31839,
    51641 => -31838,
    51642 => -31838,
    51643 => -31837,
    51644 => -31836,
    51645 => -31836,
    51646 => -31835,
    51647 => -31834,
    51648 => -31833,
    51649 => -31833,
    51650 => -31832,
    51651 => -31831,
    51652 => -31830,
    51653 => -31830,
    51654 => -31829,
    51655 => -31828,
    51656 => -31827,
    51657 => -31827,
    51658 => -31826,
    51659 => -31825,
    51660 => -31824,
    51661 => -31824,
    51662 => -31823,
    51663 => -31822,
    51664 => -31821,
    51665 => -31821,
    51666 => -31820,
    51667 => -31819,
    51668 => -31818,
    51669 => -31818,
    51670 => -31817,
    51671 => -31816,
    51672 => -31815,
    51673 => -31815,
    51674 => -31814,
    51675 => -31813,
    51676 => -31812,
    51677 => -31812,
    51678 => -31811,
    51679 => -31810,
    51680 => -31809,
    51681 => -31809,
    51682 => -31808,
    51683 => -31807,
    51684 => -31806,
    51685 => -31806,
    51686 => -31805,
    51687 => -31804,
    51688 => -31803,
    51689 => -31802,
    51690 => -31802,
    51691 => -31801,
    51692 => -31800,
    51693 => -31799,
    51694 => -31799,
    51695 => -31798,
    51696 => -31797,
    51697 => -31796,
    51698 => -31796,
    51699 => -31795,
    51700 => -31794,
    51701 => -31793,
    51702 => -31793,
    51703 => -31792,
    51704 => -31791,
    51705 => -31790,
    51706 => -31790,
    51707 => -31789,
    51708 => -31788,
    51709 => -31787,
    51710 => -31787,
    51711 => -31786,
    51712 => -31785,
    51713 => -31784,
    51714 => -31783,
    51715 => -31783,
    51716 => -31782,
    51717 => -31781,
    51718 => -31780,
    51719 => -31780,
    51720 => -31779,
    51721 => -31778,
    51722 => -31777,
    51723 => -31777,
    51724 => -31776,
    51725 => -31775,
    51726 => -31774,
    51727 => -31774,
    51728 => -31773,
    51729 => -31772,
    51730 => -31771,
    51731 => -31770,
    51732 => -31770,
    51733 => -31769,
    51734 => -31768,
    51735 => -31767,
    51736 => -31767,
    51737 => -31766,
    51738 => -31765,
    51739 => -31764,
    51740 => -31764,
    51741 => -31763,
    51742 => -31762,
    51743 => -31761,
    51744 => -31760,
    51745 => -31760,
    51746 => -31759,
    51747 => -31758,
    51748 => -31757,
    51749 => -31757,
    51750 => -31756,
    51751 => -31755,
    51752 => -31754,
    51753 => -31753,
    51754 => -31753,
    51755 => -31752,
    51756 => -31751,
    51757 => -31750,
    51758 => -31750,
    51759 => -31749,
    51760 => -31748,
    51761 => -31747,
    51762 => -31746,
    51763 => -31746,
    51764 => -31745,
    51765 => -31744,
    51766 => -31743,
    51767 => -31743,
    51768 => -31742,
    51769 => -31741,
    51770 => -31740,
    51771 => -31739,
    51772 => -31739,
    51773 => -31738,
    51774 => -31737,
    51775 => -31736,
    51776 => -31736,
    51777 => -31735,
    51778 => -31734,
    51779 => -31733,
    51780 => -31732,
    51781 => -31732,
    51782 => -31731,
    51783 => -31730,
    51784 => -31729,
    51785 => -31729,
    51786 => -31728,
    51787 => -31727,
    51788 => -31726,
    51789 => -31725,
    51790 => -31725,
    51791 => -31724,
    51792 => -31723,
    51793 => -31722,
    51794 => -31721,
    51795 => -31721,
    51796 => -31720,
    51797 => -31719,
    51798 => -31718,
    51799 => -31718,
    51800 => -31717,
    51801 => -31716,
    51802 => -31715,
    51803 => -31714,
    51804 => -31714,
    51805 => -31713,
    51806 => -31712,
    51807 => -31711,
    51808 => -31710,
    51809 => -31710,
    51810 => -31709,
    51811 => -31708,
    51812 => -31707,
    51813 => -31706,
    51814 => -31706,
    51815 => -31705,
    51816 => -31704,
    51817 => -31703,
    51818 => -31702,
    51819 => -31702,
    51820 => -31701,
    51821 => -31700,
    51822 => -31699,
    51823 => -31698,
    51824 => -31698,
    51825 => -31697,
    51826 => -31696,
    51827 => -31695,
    51828 => -31695,
    51829 => -31694,
    51830 => -31693,
    51831 => -31692,
    51832 => -31691,
    51833 => -31691,
    51834 => -31690,
    51835 => -31689,
    51836 => -31688,
    51837 => -31687,
    51838 => -31687,
    51839 => -31686,
    51840 => -31685,
    51841 => -31684,
    51842 => -31683,
    51843 => -31683,
    51844 => -31682,
    51845 => -31681,
    51846 => -31680,
    51847 => -31679,
    51848 => -31679,
    51849 => -31678,
    51850 => -31677,
    51851 => -31676,
    51852 => -31675,
    51853 => -31674,
    51854 => -31674,
    51855 => -31673,
    51856 => -31672,
    51857 => -31671,
    51858 => -31670,
    51859 => -31670,
    51860 => -31669,
    51861 => -31668,
    51862 => -31667,
    51863 => -31666,
    51864 => -31666,
    51865 => -31665,
    51866 => -31664,
    51867 => -31663,
    51868 => -31662,
    51869 => -31662,
    51870 => -31661,
    51871 => -31660,
    51872 => -31659,
    51873 => -31658,
    51874 => -31658,
    51875 => -31657,
    51876 => -31656,
    51877 => -31655,
    51878 => -31654,
    51879 => -31653,
    51880 => -31653,
    51881 => -31652,
    51882 => -31651,
    51883 => -31650,
    51884 => -31649,
    51885 => -31649,
    51886 => -31648,
    51887 => -31647,
    51888 => -31646,
    51889 => -31645,
    51890 => -31645,
    51891 => -31644,
    51892 => -31643,
    51893 => -31642,
    51894 => -31641,
    51895 => -31640,
    51896 => -31640,
    51897 => -31639,
    51898 => -31638,
    51899 => -31637,
    51900 => -31636,
    51901 => -31636,
    51902 => -31635,
    51903 => -31634,
    51904 => -31633,
    51905 => -31632,
    51906 => -31631,
    51907 => -31631,
    51908 => -31630,
    51909 => -31629,
    51910 => -31628,
    51911 => -31627,
    51912 => -31627,
    51913 => -31626,
    51914 => -31625,
    51915 => -31624,
    51916 => -31623,
    51917 => -31622,
    51918 => -31622,
    51919 => -31621,
    51920 => -31620,
    51921 => -31619,
    51922 => -31618,
    51923 => -31617,
    51924 => -31617,
    51925 => -31616,
    51926 => -31615,
    51927 => -31614,
    51928 => -31613,
    51929 => -31613,
    51930 => -31612,
    51931 => -31611,
    51932 => -31610,
    51933 => -31609,
    51934 => -31608,
    51935 => -31608,
    51936 => -31607,
    51937 => -31606,
    51938 => -31605,
    51939 => -31604,
    51940 => -31603,
    51941 => -31603,
    51942 => -31602,
    51943 => -31601,
    51944 => -31600,
    51945 => -31599,
    51946 => -31598,
    51947 => -31598,
    51948 => -31597,
    51949 => -31596,
    51950 => -31595,
    51951 => -31594,
    51952 => -31593,
    51953 => -31593,
    51954 => -31592,
    51955 => -31591,
    51956 => -31590,
    51957 => -31589,
    51958 => -31588,
    51959 => -31588,
    51960 => -31587,
    51961 => -31586,
    51962 => -31585,
    51963 => -31584,
    51964 => -31583,
    51965 => -31583,
    51966 => -31582,
    51967 => -31581,
    51968 => -31580,
    51969 => -31579,
    51970 => -31578,
    51971 => -31578,
    51972 => -31577,
    51973 => -31576,
    51974 => -31575,
    51975 => -31574,
    51976 => -31573,
    51977 => -31572,
    51978 => -31572,
    51979 => -31571,
    51980 => -31570,
    51981 => -31569,
    51982 => -31568,
    51983 => -31567,
    51984 => -31567,
    51985 => -31566,
    51986 => -31565,
    51987 => -31564,
    51988 => -31563,
    51989 => -31562,
    51990 => -31562,
    51991 => -31561,
    51992 => -31560,
    51993 => -31559,
    51994 => -31558,
    51995 => -31557,
    51996 => -31556,
    51997 => -31556,
    51998 => -31555,
    51999 => -31554,
    52000 => -31553,
    52001 => -31552,
    52002 => -31551,
    52003 => -31551,
    52004 => -31550,
    52005 => -31549,
    52006 => -31548,
    52007 => -31547,
    52008 => -31546,
    52009 => -31545,
    52010 => -31545,
    52011 => -31544,
    52012 => -31543,
    52013 => -31542,
    52014 => -31541,
    52015 => -31540,
    52016 => -31539,
    52017 => -31539,
    52018 => -31538,
    52019 => -31537,
    52020 => -31536,
    52021 => -31535,
    52022 => -31534,
    52023 => -31534,
    52024 => -31533,
    52025 => -31532,
    52026 => -31531,
    52027 => -31530,
    52028 => -31529,
    52029 => -31528,
    52030 => -31528,
    52031 => -31527,
    52032 => -31526,
    52033 => -31525,
    52034 => -31524,
    52035 => -31523,
    52036 => -31522,
    52037 => -31522,
    52038 => -31521,
    52039 => -31520,
    52040 => -31519,
    52041 => -31518,
    52042 => -31517,
    52043 => -31516,
    52044 => -31516,
    52045 => -31515,
    52046 => -31514,
    52047 => -31513,
    52048 => -31512,
    52049 => -31511,
    52050 => -31510,
    52051 => -31510,
    52052 => -31509,
    52053 => -31508,
    52054 => -31507,
    52055 => -31506,
    52056 => -31505,
    52057 => -31504,
    52058 => -31503,
    52059 => -31503,
    52060 => -31502,
    52061 => -31501,
    52062 => -31500,
    52063 => -31499,
    52064 => -31498,
    52065 => -31497,
    52066 => -31497,
    52067 => -31496,
    52068 => -31495,
    52069 => -31494,
    52070 => -31493,
    52071 => -31492,
    52072 => -31491,
    52073 => -31490,
    52074 => -31490,
    52075 => -31489,
    52076 => -31488,
    52077 => -31487,
    52078 => -31486,
    52079 => -31485,
    52080 => -31484,
    52081 => -31484,
    52082 => -31483,
    52083 => -31482,
    52084 => -31481,
    52085 => -31480,
    52086 => -31479,
    52087 => -31478,
    52088 => -31477,
    52089 => -31477,
    52090 => -31476,
    52091 => -31475,
    52092 => -31474,
    52093 => -31473,
    52094 => -31472,
    52095 => -31471,
    52096 => -31470,
    52097 => -31470,
    52098 => -31469,
    52099 => -31468,
    52100 => -31467,
    52101 => -31466,
    52102 => -31465,
    52103 => -31464,
    52104 => -31463,
    52105 => -31463,
    52106 => -31462,
    52107 => -31461,
    52108 => -31460,
    52109 => -31459,
    52110 => -31458,
    52111 => -31457,
    52112 => -31456,
    52113 => -31456,
    52114 => -31455,
    52115 => -31454,
    52116 => -31453,
    52117 => -31452,
    52118 => -31451,
    52119 => -31450,
    52120 => -31449,
    52121 => -31448,
    52122 => -31448,
    52123 => -31447,
    52124 => -31446,
    52125 => -31445,
    52126 => -31444,
    52127 => -31443,
    52128 => -31442,
    52129 => -31441,
    52130 => -31441,
    52131 => -31440,
    52132 => -31439,
    52133 => -31438,
    52134 => -31437,
    52135 => -31436,
    52136 => -31435,
    52137 => -31434,
    52138 => -31433,
    52139 => -31433,
    52140 => -31432,
    52141 => -31431,
    52142 => -31430,
    52143 => -31429,
    52144 => -31428,
    52145 => -31427,
    52146 => -31426,
    52147 => -31425,
    52148 => -31425,
    52149 => -31424,
    52150 => -31423,
    52151 => -31422,
    52152 => -31421,
    52153 => -31420,
    52154 => -31419,
    52155 => -31418,
    52156 => -31417,
    52157 => -31417,
    52158 => -31416,
    52159 => -31415,
    52160 => -31414,
    52161 => -31413,
    52162 => -31412,
    52163 => -31411,
    52164 => -31410,
    52165 => -31409,
    52166 => -31408,
    52167 => -31408,
    52168 => -31407,
    52169 => -31406,
    52170 => -31405,
    52171 => -31404,
    52172 => -31403,
    52173 => -31402,
    52174 => -31401,
    52175 => -31400,
    52176 => -31400,
    52177 => -31399,
    52178 => -31398,
    52179 => -31397,
    52180 => -31396,
    52181 => -31395,
    52182 => -31394,
    52183 => -31393,
    52184 => -31392,
    52185 => -31391,
    52186 => -31391,
    52187 => -31390,
    52188 => -31389,
    52189 => -31388,
    52190 => -31387,
    52191 => -31386,
    52192 => -31385,
    52193 => -31384,
    52194 => -31383,
    52195 => -31382,
    52196 => -31381,
    52197 => -31381,
    52198 => -31380,
    52199 => -31379,
    52200 => -31378,
    52201 => -31377,
    52202 => -31376,
    52203 => -31375,
    52204 => -31374,
    52205 => -31373,
    52206 => -31372,
    52207 => -31372,
    52208 => -31371,
    52209 => -31370,
    52210 => -31369,
    52211 => -31368,
    52212 => -31367,
    52213 => -31366,
    52214 => -31365,
    52215 => -31364,
    52216 => -31363,
    52217 => -31362,
    52218 => -31362,
    52219 => -31361,
    52220 => -31360,
    52221 => -31359,
    52222 => -31358,
    52223 => -31357,
    52224 => -31356,
    52225 => -31355,
    52226 => -31354,
    52227 => -31353,
    52228 => -31352,
    52229 => -31352,
    52230 => -31351,
    52231 => -31350,
    52232 => -31349,
    52233 => -31348,
    52234 => -31347,
    52235 => -31346,
    52236 => -31345,
    52237 => -31344,
    52238 => -31343,
    52239 => -31342,
    52240 => -31341,
    52241 => -31341,
    52242 => -31340,
    52243 => -31339,
    52244 => -31338,
    52245 => -31337,
    52246 => -31336,
    52247 => -31335,
    52248 => -31334,
    52249 => -31333,
    52250 => -31332,
    52251 => -31331,
    52252 => -31330,
    52253 => -31329,
    52254 => -31329,
    52255 => -31328,
    52256 => -31327,
    52257 => -31326,
    52258 => -31325,
    52259 => -31324,
    52260 => -31323,
    52261 => -31322,
    52262 => -31321,
    52263 => -31320,
    52264 => -31319,
    52265 => -31318,
    52266 => -31318,
    52267 => -31317,
    52268 => -31316,
    52269 => -31315,
    52270 => -31314,
    52271 => -31313,
    52272 => -31312,
    52273 => -31311,
    52274 => -31310,
    52275 => -31309,
    52276 => -31308,
    52277 => -31307,
    52278 => -31306,
    52279 => -31305,
    52280 => -31305,
    52281 => -31304,
    52282 => -31303,
    52283 => -31302,
    52284 => -31301,
    52285 => -31300,
    52286 => -31299,
    52287 => -31298,
    52288 => -31297,
    52289 => -31296,
    52290 => -31295,
    52291 => -31294,
    52292 => -31293,
    52293 => -31292,
    52294 => -31292,
    52295 => -31291,
    52296 => -31290,
    52297 => -31289,
    52298 => -31288,
    52299 => -31287,
    52300 => -31286,
    52301 => -31285,
    52302 => -31284,
    52303 => -31283,
    52304 => -31282,
    52305 => -31281,
    52306 => -31280,
    52307 => -31279,
    52308 => -31278,
    52309 => -31278,
    52310 => -31277,
    52311 => -31276,
    52312 => -31275,
    52313 => -31274,
    52314 => -31273,
    52315 => -31272,
    52316 => -31271,
    52317 => -31270,
    52318 => -31269,
    52319 => -31268,
    52320 => -31267,
    52321 => -31266,
    52322 => -31265,
    52323 => -31264,
    52324 => -31263,
    52325 => -31262,
    52326 => -31262,
    52327 => -31261,
    52328 => -31260,
    52329 => -31259,
    52330 => -31258,
    52331 => -31257,
    52332 => -31256,
    52333 => -31255,
    52334 => -31254,
    52335 => -31253,
    52336 => -31252,
    52337 => -31251,
    52338 => -31250,
    52339 => -31249,
    52340 => -31248,
    52341 => -31247,
    52342 => -31246,
    52343 => -31246,
    52344 => -31245,
    52345 => -31244,
    52346 => -31243,
    52347 => -31242,
    52348 => -31241,
    52349 => -31240,
    52350 => -31239,
    52351 => -31238,
    52352 => -31237,
    52353 => -31236,
    52354 => -31235,
    52355 => -31234,
    52356 => -31233,
    52357 => -31232,
    52358 => -31231,
    52359 => -31230,
    52360 => -31229,
    52361 => -31228,
    52362 => -31227,
    52363 => -31227,
    52364 => -31226,
    52365 => -31225,
    52366 => -31224,
    52367 => -31223,
    52368 => -31222,
    52369 => -31221,
    52370 => -31220,
    52371 => -31219,
    52372 => -31218,
    52373 => -31217,
    52374 => -31216,
    52375 => -31215,
    52376 => -31214,
    52377 => -31213,
    52378 => -31212,
    52379 => -31211,
    52380 => -31210,
    52381 => -31209,
    52382 => -31208,
    52383 => -31207,
    52384 => -31206,
    52385 => -31206,
    52386 => -31205,
    52387 => -31204,
    52388 => -31203,
    52389 => -31202,
    52390 => -31201,
    52391 => -31200,
    52392 => -31199,
    52393 => -31198,
    52394 => -31197,
    52395 => -31196,
    52396 => -31195,
    52397 => -31194,
    52398 => -31193,
    52399 => -31192,
    52400 => -31191,
    52401 => -31190,
    52402 => -31189,
    52403 => -31188,
    52404 => -31187,
    52405 => -31186,
    52406 => -31185,
    52407 => -31184,
    52408 => -31183,
    52409 => -31182,
    52410 => -31181,
    52411 => -31181,
    52412 => -31180,
    52413 => -31179,
    52414 => -31178,
    52415 => -31177,
    52416 => -31176,
    52417 => -31175,
    52418 => -31174,
    52419 => -31173,
    52420 => -31172,
    52421 => -31171,
    52422 => -31170,
    52423 => -31169,
    52424 => -31168,
    52425 => -31167,
    52426 => -31166,
    52427 => -31165,
    52428 => -31164,
    52429 => -31163,
    52430 => -31162,
    52431 => -31161,
    52432 => -31160,
    52433 => -31159,
    52434 => -31158,
    52435 => -31157,
    52436 => -31156,
    52437 => -31155,
    52438 => -31154,
    52439 => -31153,
    52440 => -31152,
    52441 => -31151,
    52442 => -31150,
    52443 => -31149,
    52444 => -31148,
    52445 => -31148,
    52446 => -31147,
    52447 => -31146,
    52448 => -31145,
    52449 => -31144,
    52450 => -31143,
    52451 => -31142,
    52452 => -31141,
    52453 => -31140,
    52454 => -31139,
    52455 => -31138,
    52456 => -31137,
    52457 => -31136,
    52458 => -31135,
    52459 => -31134,
    52460 => -31133,
    52461 => -31132,
    52462 => -31131,
    52463 => -31130,
    52464 => -31129,
    52465 => -31128,
    52466 => -31127,
    52467 => -31126,
    52468 => -31125,
    52469 => -31124,
    52470 => -31123,
    52471 => -31122,
    52472 => -31121,
    52473 => -31120,
    52474 => -31119,
    52475 => -31118,
    52476 => -31117,
    52477 => -31116,
    52478 => -31115,
    52479 => -31114,
    52480 => -31113,
    52481 => -31112,
    52482 => -31111,
    52483 => -31110,
    52484 => -31109,
    52485 => -31108,
    52486 => -31107,
    52487 => -31106,
    52488 => -31105,
    52489 => -31104,
    52490 => -31103,
    52491 => -31102,
    52492 => -31101,
    52493 => -31100,
    52494 => -31099,
    52495 => -31098,
    52496 => -31097,
    52497 => -31096,
    52498 => -31095,
    52499 => -31094,
    52500 => -31093,
    52501 => -31092,
    52502 => -31091,
    52503 => -31090,
    52504 => -31089,
    52505 => -31088,
    52506 => -31087,
    52507 => -31086,
    52508 => -31085,
    52509 => -31084,
    52510 => -31083,
    52511 => -31083,
    52512 => -31082,
    52513 => -31081,
    52514 => -31080,
    52515 => -31079,
    52516 => -31078,
    52517 => -31077,
    52518 => -31076,
    52519 => -31075,
    52520 => -31074,
    52521 => -31073,
    52522 => -31072,
    52523 => -31071,
    52524 => -31070,
    52525 => -31069,
    52526 => -31068,
    52527 => -31067,
    52528 => -31066,
    52529 => -31065,
    52530 => -31064,
    52531 => -31063,
    52532 => -31062,
    52533 => -31061,
    52534 => -31060,
    52535 => -31059,
    52536 => -31058,
    52537 => -31057,
    52538 => -31056,
    52539 => -31055,
    52540 => -31054,
    52541 => -31053,
    52542 => -31052,
    52543 => -31051,
    52544 => -31050,
    52545 => -31049,
    52546 => -31048,
    52547 => -31047,
    52548 => -31046,
    52549 => -31045,
    52550 => -31044,
    52551 => -31043,
    52552 => -31041,
    52553 => -31040,
    52554 => -31039,
    52555 => -31038,
    52556 => -31037,
    52557 => -31036,
    52558 => -31035,
    52559 => -31034,
    52560 => -31033,
    52561 => -31032,
    52562 => -31031,
    52563 => -31030,
    52564 => -31029,
    52565 => -31028,
    52566 => -31027,
    52567 => -31026,
    52568 => -31025,
    52569 => -31024,
    52570 => -31023,
    52571 => -31022,
    52572 => -31021,
    52573 => -31020,
    52574 => -31019,
    52575 => -31018,
    52576 => -31017,
    52577 => -31016,
    52578 => -31015,
    52579 => -31014,
    52580 => -31013,
    52581 => -31012,
    52582 => -31011,
    52583 => -31010,
    52584 => -31009,
    52585 => -31008,
    52586 => -31007,
    52587 => -31006,
    52588 => -31005,
    52589 => -31004,
    52590 => -31003,
    52591 => -31002,
    52592 => -31001,
    52593 => -31000,
    52594 => -30999,
    52595 => -30998,
    52596 => -30997,
    52597 => -30996,
    52598 => -30995,
    52599 => -30994,
    52600 => -30993,
    52601 => -30992,
    52602 => -30991,
    52603 => -30990,
    52604 => -30989,
    52605 => -30988,
    52606 => -30987,
    52607 => -30986,
    52608 => -30985,
    52609 => -30984,
    52610 => -30983,
    52611 => -30982,
    52612 => -30981,
    52613 => -30980,
    52614 => -30979,
    52615 => -30978,
    52616 => -30977,
    52617 => -30976,
    52618 => -30974,
    52619 => -30973,
    52620 => -30972,
    52621 => -30971,
    52622 => -30970,
    52623 => -30969,
    52624 => -30968,
    52625 => -30967,
    52626 => -30966,
    52627 => -30965,
    52628 => -30964,
    52629 => -30963,
    52630 => -30962,
    52631 => -30961,
    52632 => -30960,
    52633 => -30959,
    52634 => -30958,
    52635 => -30957,
    52636 => -30956,
    52637 => -30955,
    52638 => -30954,
    52639 => -30953,
    52640 => -30952,
    52641 => -30951,
    52642 => -30950,
    52643 => -30949,
    52644 => -30948,
    52645 => -30947,
    52646 => -30946,
    52647 => -30945,
    52648 => -30944,
    52649 => -30943,
    52650 => -30942,
    52651 => -30941,
    52652 => -30939,
    52653 => -30938,
    52654 => -30937,
    52655 => -30936,
    52656 => -30935,
    52657 => -30934,
    52658 => -30933,
    52659 => -30932,
    52660 => -30931,
    52661 => -30930,
    52662 => -30929,
    52663 => -30928,
    52664 => -30927,
    52665 => -30926,
    52666 => -30925,
    52667 => -30924,
    52668 => -30923,
    52669 => -30922,
    52670 => -30921,
    52671 => -30920,
    52672 => -30919,
    52673 => -30918,
    52674 => -30917,
    52675 => -30916,
    52676 => -30915,
    52677 => -30914,
    52678 => -30912,
    52679 => -30911,
    52680 => -30910,
    52681 => -30909,
    52682 => -30908,
    52683 => -30907,
    52684 => -30906,
    52685 => -30905,
    52686 => -30904,
    52687 => -30903,
    52688 => -30902,
    52689 => -30901,
    52690 => -30900,
    52691 => -30899,
    52692 => -30898,
    52693 => -30897,
    52694 => -30896,
    52695 => -30895,
    52696 => -30894,
    52697 => -30893,
    52698 => -30892,
    52699 => -30891,
    52700 => -30889,
    52701 => -30888,
    52702 => -30887,
    52703 => -30886,
    52704 => -30885,
    52705 => -30884,
    52706 => -30883,
    52707 => -30882,
    52708 => -30881,
    52709 => -30880,
    52710 => -30879,
    52711 => -30878,
    52712 => -30877,
    52713 => -30876,
    52714 => -30875,
    52715 => -30874,
    52716 => -30873,
    52717 => -30872,
    52718 => -30871,
    52719 => -30870,
    52720 => -30868,
    52721 => -30867,
    52722 => -30866,
    52723 => -30865,
    52724 => -30864,
    52725 => -30863,
    52726 => -30862,
    52727 => -30861,
    52728 => -30860,
    52729 => -30859,
    52730 => -30858,
    52731 => -30857,
    52732 => -30856,
    52733 => -30855,
    52734 => -30854,
    52735 => -30853,
    52736 => -30852,
    52737 => -30851,
    52738 => -30849,
    52739 => -30848,
    52740 => -30847,
    52741 => -30846,
    52742 => -30845,
    52743 => -30844,
    52744 => -30843,
    52745 => -30842,
    52746 => -30841,
    52747 => -30840,
    52748 => -30839,
    52749 => -30838,
    52750 => -30837,
    52751 => -30836,
    52752 => -30835,
    52753 => -30834,
    52754 => -30832,
    52755 => -30831,
    52756 => -30830,
    52757 => -30829,
    52758 => -30828,
    52759 => -30827,
    52760 => -30826,
    52761 => -30825,
    52762 => -30824,
    52763 => -30823,
    52764 => -30822,
    52765 => -30821,
    52766 => -30820,
    52767 => -30819,
    52768 => -30818,
    52769 => -30816,
    52770 => -30815,
    52771 => -30814,
    52772 => -30813,
    52773 => -30812,
    52774 => -30811,
    52775 => -30810,
    52776 => -30809,
    52777 => -30808,
    52778 => -30807,
    52779 => -30806,
    52780 => -30805,
    52781 => -30804,
    52782 => -30803,
    52783 => -30802,
    52784 => -30800,
    52785 => -30799,
    52786 => -30798,
    52787 => -30797,
    52788 => -30796,
    52789 => -30795,
    52790 => -30794,
    52791 => -30793,
    52792 => -30792,
    52793 => -30791,
    52794 => -30790,
    52795 => -30789,
    52796 => -30788,
    52797 => -30786,
    52798 => -30785,
    52799 => -30784,
    52800 => -30783,
    52801 => -30782,
    52802 => -30781,
    52803 => -30780,
    52804 => -30779,
    52805 => -30778,
    52806 => -30777,
    52807 => -30776,
    52808 => -30775,
    52809 => -30774,
    52810 => -30772,
    52811 => -30771,
    52812 => -30770,
    52813 => -30769,
    52814 => -30768,
    52815 => -30767,
    52816 => -30766,
    52817 => -30765,
    52818 => -30764,
    52819 => -30763,
    52820 => -30762,
    52821 => -30761,
    52822 => -30760,
    52823 => -30758,
    52824 => -30757,
    52825 => -30756,
    52826 => -30755,
    52827 => -30754,
    52828 => -30753,
    52829 => -30752,
    52830 => -30751,
    52831 => -30750,
    52832 => -30749,
    52833 => -30748,
    52834 => -30746,
    52835 => -30745,
    52836 => -30744,
    52837 => -30743,
    52838 => -30742,
    52839 => -30741,
    52840 => -30740,
    52841 => -30739,
    52842 => -30738,
    52843 => -30737,
    52844 => -30736,
    52845 => -30735,
    52846 => -30733,
    52847 => -30732,
    52848 => -30731,
    52849 => -30730,
    52850 => -30729,
    52851 => -30728,
    52852 => -30727,
    52853 => -30726,
    52854 => -30725,
    52855 => -30724,
    52856 => -30723,
    52857 => -30721,
    52858 => -30720,
    52859 => -30719,
    52860 => -30718,
    52861 => -30717,
    52862 => -30716,
    52863 => -30715,
    52864 => -30714,
    52865 => -30713,
    52866 => -30712,
    52867 => -30711,
    52868 => -30709,
    52869 => -30708,
    52870 => -30707,
    52871 => -30706,
    52872 => -30705,
    52873 => -30704,
    52874 => -30703,
    52875 => -30702,
    52876 => -30701,
    52877 => -30700,
    52878 => -30698,
    52879 => -30697,
    52880 => -30696,
    52881 => -30695,
    52882 => -30694,
    52883 => -30693,
    52884 => -30692,
    52885 => -30691,
    52886 => -30690,
    52887 => -30689,
    52888 => -30687,
    52889 => -30686,
    52890 => -30685,
    52891 => -30684,
    52892 => -30683,
    52893 => -30682,
    52894 => -30681,
    52895 => -30680,
    52896 => -30679,
    52897 => -30678,
    52898 => -30676,
    52899 => -30675,
    52900 => -30674,
    52901 => -30673,
    52902 => -30672,
    52903 => -30671,
    52904 => -30670,
    52905 => -30669,
    52906 => -30668,
    52907 => -30666,
    52908 => -30665,
    52909 => -30664,
    52910 => -30663,
    52911 => -30662,
    52912 => -30661,
    52913 => -30660,
    52914 => -30659,
    52915 => -30658,
    52916 => -30656,
    52917 => -30655,
    52918 => -30654,
    52919 => -30653,
    52920 => -30652,
    52921 => -30651,
    52922 => -30650,
    52923 => -30649,
    52924 => -30648,
    52925 => -30646,
    52926 => -30645,
    52927 => -30644,
    52928 => -30643,
    52929 => -30642,
    52930 => -30641,
    52931 => -30640,
    52932 => -30639,
    52933 => -30638,
    52934 => -30636,
    52935 => -30635,
    52936 => -30634,
    52937 => -30633,
    52938 => -30632,
    52939 => -30631,
    52940 => -30630,
    52941 => -30629,
    52942 => -30628,
    52943 => -30626,
    52944 => -30625,
    52945 => -30624,
    52946 => -30623,
    52947 => -30622,
    52948 => -30621,
    52949 => -30620,
    52950 => -30619,
    52951 => -30617,
    52952 => -30616,
    52953 => -30615,
    52954 => -30614,
    52955 => -30613,
    52956 => -30612,
    52957 => -30611,
    52958 => -30610,
    52959 => -30609,
    52960 => -30607,
    52961 => -30606,
    52962 => -30605,
    52963 => -30604,
    52964 => -30603,
    52965 => -30602,
    52966 => -30601,
    52967 => -30600,
    52968 => -30598,
    52969 => -30597,
    52970 => -30596,
    52971 => -30595,
    52972 => -30594,
    52973 => -30593,
    52974 => -30592,
    52975 => -30591,
    52976 => -30589,
    52977 => -30588,
    52978 => -30587,
    52979 => -30586,
    52980 => -30585,
    52981 => -30584,
    52982 => -30583,
    52983 => -30582,
    52984 => -30580,
    52985 => -30579,
    52986 => -30578,
    52987 => -30577,
    52988 => -30576,
    52989 => -30575,
    52990 => -30574,
    52991 => -30573,
    52992 => -30571,
    52993 => -30570,
    52994 => -30569,
    52995 => -30568,
    52996 => -30567,
    52997 => -30566,
    52998 => -30565,
    52999 => -30563,
    53000 => -30562,
    53001 => -30561,
    53002 => -30560,
    53003 => -30559,
    53004 => -30558,
    53005 => -30557,
    53006 => -30556,
    53007 => -30554,
    53008 => -30553,
    53009 => -30552,
    53010 => -30551,
    53011 => -30550,
    53012 => -30549,
    53013 => -30548,
    53014 => -30546,
    53015 => -30545,
    53016 => -30544,
    53017 => -30543,
    53018 => -30542,
    53019 => -30541,
    53020 => -30540,
    53021 => -30538,
    53022 => -30537,
    53023 => -30536,
    53024 => -30535,
    53025 => -30534,
    53026 => -30533,
    53027 => -30532,
    53028 => -30530,
    53029 => -30529,
    53030 => -30528,
    53031 => -30527,
    53032 => -30526,
    53033 => -30525,
    53034 => -30524,
    53035 => -30522,
    53036 => -30521,
    53037 => -30520,
    53038 => -30519,
    53039 => -30518,
    53040 => -30517,
    53041 => -30516,
    53042 => -30514,
    53043 => -30513,
    53044 => -30512,
    53045 => -30511,
    53046 => -30510,
    53047 => -30509,
    53048 => -30508,
    53049 => -30506,
    53050 => -30505,
    53051 => -30504,
    53052 => -30503,
    53053 => -30502,
    53054 => -30501,
    53055 => -30500,
    53056 => -30498,
    53057 => -30497,
    53058 => -30496,
    53059 => -30495,
    53060 => -30494,
    53061 => -30493,
    53062 => -30492,
    53063 => -30490,
    53064 => -30489,
    53065 => -30488,
    53066 => -30487,
    53067 => -30486,
    53068 => -30485,
    53069 => -30483,
    53070 => -30482,
    53071 => -30481,
    53072 => -30480,
    53073 => -30479,
    53074 => -30478,
    53075 => -30477,
    53076 => -30475,
    53077 => -30474,
    53078 => -30473,
    53079 => -30472,
    53080 => -30471,
    53081 => -30470,
    53082 => -30468,
    53083 => -30467,
    53084 => -30466,
    53085 => -30465,
    53086 => -30464,
    53087 => -30463,
    53088 => -30462,
    53089 => -30460,
    53090 => -30459,
    53091 => -30458,
    53092 => -30457,
    53093 => -30456,
    53094 => -30455,
    53095 => -30453,
    53096 => -30452,
    53097 => -30451,
    53098 => -30450,
    53099 => -30449,
    53100 => -30448,
    53101 => -30446,
    53102 => -30445,
    53103 => -30444,
    53104 => -30443,
    53105 => -30442,
    53106 => -30441,
    53107 => -30439,
    53108 => -30438,
    53109 => -30437,
    53110 => -30436,
    53111 => -30435,
    53112 => -30434,
    53113 => -30433,
    53114 => -30431,
    53115 => -30430,
    53116 => -30429,
    53117 => -30428,
    53118 => -30427,
    53119 => -30426,
    53120 => -30424,
    53121 => -30423,
    53122 => -30422,
    53123 => -30421,
    53124 => -30420,
    53125 => -30419,
    53126 => -30417,
    53127 => -30416,
    53128 => -30415,
    53129 => -30414,
    53130 => -30413,
    53131 => -30412,
    53132 => -30410,
    53133 => -30409,
    53134 => -30408,
    53135 => -30407,
    53136 => -30406,
    53137 => -30404,
    53138 => -30403,
    53139 => -30402,
    53140 => -30401,
    53141 => -30400,
    53142 => -30399,
    53143 => -30397,
    53144 => -30396,
    53145 => -30395,
    53146 => -30394,
    53147 => -30393,
    53148 => -30392,
    53149 => -30390,
    53150 => -30389,
    53151 => -30388,
    53152 => -30387,
    53153 => -30386,
    53154 => -30385,
    53155 => -30383,
    53156 => -30382,
    53157 => -30381,
    53158 => -30380,
    53159 => -30379,
    53160 => -30377,
    53161 => -30376,
    53162 => -30375,
    53163 => -30374,
    53164 => -30373,
    53165 => -30372,
    53166 => -30370,
    53167 => -30369,
    53168 => -30368,
    53169 => -30367,
    53170 => -30366,
    53171 => -30365,
    53172 => -30363,
    53173 => -30362,
    53174 => -30361,
    53175 => -30360,
    53176 => -30359,
    53177 => -30357,
    53178 => -30356,
    53179 => -30355,
    53180 => -30354,
    53181 => -30353,
    53182 => -30351,
    53183 => -30350,
    53184 => -30349,
    53185 => -30348,
    53186 => -30347,
    53187 => -30346,
    53188 => -30344,
    53189 => -30343,
    53190 => -30342,
    53191 => -30341,
    53192 => -30340,
    53193 => -30338,
    53194 => -30337,
    53195 => -30336,
    53196 => -30335,
    53197 => -30334,
    53198 => -30333,
    53199 => -30331,
    53200 => -30330,
    53201 => -30329,
    53202 => -30328,
    53203 => -30327,
    53204 => -30325,
    53205 => -30324,
    53206 => -30323,
    53207 => -30322,
    53208 => -30321,
    53209 => -30319,
    53210 => -30318,
    53211 => -30317,
    53212 => -30316,
    53213 => -30315,
    53214 => -30313,
    53215 => -30312,
    53216 => -30311,
    53217 => -30310,
    53218 => -30309,
    53219 => -30308,
    53220 => -30306,
    53221 => -30305,
    53222 => -30304,
    53223 => -30303,
    53224 => -30302,
    53225 => -30300,
    53226 => -30299,
    53227 => -30298,
    53228 => -30297,
    53229 => -30296,
    53230 => -30294,
    53231 => -30293,
    53232 => -30292,
    53233 => -30291,
    53234 => -30290,
    53235 => -30288,
    53236 => -30287,
    53237 => -30286,
    53238 => -30285,
    53239 => -30284,
    53240 => -30282,
    53241 => -30281,
    53242 => -30280,
    53243 => -30279,
    53244 => -30278,
    53245 => -30276,
    53246 => -30275,
    53247 => -30274,
    53248 => -30273,
    53249 => -30272,
    53250 => -30270,
    53251 => -30269,
    53252 => -30268,
    53253 => -30267,
    53254 => -30266,
    53255 => -30264,
    53256 => -30263,
    53257 => -30262,
    53258 => -30261,
    53259 => -30260,
    53260 => -30258,
    53261 => -30257,
    53262 => -30256,
    53263 => -30255,
    53264 => -30253,
    53265 => -30252,
    53266 => -30251,
    53267 => -30250,
    53268 => -30249,
    53269 => -30247,
    53270 => -30246,
    53271 => -30245,
    53272 => -30244,
    53273 => -30243,
    53274 => -30241,
    53275 => -30240,
    53276 => -30239,
    53277 => -30238,
    53278 => -30237,
    53279 => -30235,
    53280 => -30234,
    53281 => -30233,
    53282 => -30232,
    53283 => -30231,
    53284 => -30229,
    53285 => -30228,
    53286 => -30227,
    53287 => -30226,
    53288 => -30224,
    53289 => -30223,
    53290 => -30222,
    53291 => -30221,
    53292 => -30220,
    53293 => -30218,
    53294 => -30217,
    53295 => -30216,
    53296 => -30215,
    53297 => -30214,
    53298 => -30212,
    53299 => -30211,
    53300 => -30210,
    53301 => -30209,
    53302 => -30207,
    53303 => -30206,
    53304 => -30205,
    53305 => -30204,
    53306 => -30203,
    53307 => -30201,
    53308 => -30200,
    53309 => -30199,
    53310 => -30198,
    53311 => -30196,
    53312 => -30195,
    53313 => -30194,
    53314 => -30193,
    53315 => -30192,
    53316 => -30190,
    53317 => -30189,
    53318 => -30188,
    53319 => -30187,
    53320 => -30185,
    53321 => -30184,
    53322 => -30183,
    53323 => -30182,
    53324 => -30181,
    53325 => -30179,
    53326 => -30178,
    53327 => -30177,
    53328 => -30176,
    53329 => -30174,
    53330 => -30173,
    53331 => -30172,
    53332 => -30171,
    53333 => -30170,
    53334 => -30168,
    53335 => -30167,
    53336 => -30166,
    53337 => -30165,
    53338 => -30163,
    53339 => -30162,
    53340 => -30161,
    53341 => -30160,
    53342 => -30159,
    53343 => -30157,
    53344 => -30156,
    53345 => -30155,
    53346 => -30154,
    53347 => -30152,
    53348 => -30151,
    53349 => -30150,
    53350 => -30149,
    53351 => -30147,
    53352 => -30146,
    53353 => -30145,
    53354 => -30144,
    53355 => -30143,
    53356 => -30141,
    53357 => -30140,
    53358 => -30139,
    53359 => -30138,
    53360 => -30136,
    53361 => -30135,
    53362 => -30134,
    53363 => -30133,
    53364 => -30131,
    53365 => -30130,
    53366 => -30129,
    53367 => -30128,
    53368 => -30126,
    53369 => -30125,
    53370 => -30124,
    53371 => -30123,
    53372 => -30122,
    53373 => -30120,
    53374 => -30119,
    53375 => -30118,
    53376 => -30117,
    53377 => -30115,
    53378 => -30114,
    53379 => -30113,
    53380 => -30112,
    53381 => -30110,
    53382 => -30109,
    53383 => -30108,
    53384 => -30107,
    53385 => -30105,
    53386 => -30104,
    53387 => -30103,
    53388 => -30102,
    53389 => -30100,
    53390 => -30099,
    53391 => -30098,
    53392 => -30097,
    53393 => -30096,
    53394 => -30094,
    53395 => -30093,
    53396 => -30092,
    53397 => -30091,
    53398 => -30089,
    53399 => -30088,
    53400 => -30087,
    53401 => -30086,
    53402 => -30084,
    53403 => -30083,
    53404 => -30082,
    53405 => -30081,
    53406 => -30079,
    53407 => -30078,
    53408 => -30077,
    53409 => -30076,
    53410 => -30074,
    53411 => -30073,
    53412 => -30072,
    53413 => -30071,
    53414 => -30069,
    53415 => -30068,
    53416 => -30067,
    53417 => -30066,
    53418 => -30064,
    53419 => -30063,
    53420 => -30062,
    53421 => -30061,
    53422 => -30059,
    53423 => -30058,
    53424 => -30057,
    53425 => -30056,
    53426 => -30054,
    53427 => -30053,
    53428 => -30052,
    53429 => -30051,
    53430 => -30049,
    53431 => -30048,
    53432 => -30047,
    53433 => -30046,
    53434 => -30044,
    53435 => -30043,
    53436 => -30042,
    53437 => -30041,
    53438 => -30039,
    53439 => -30038,
    53440 => -30037,
    53441 => -30036,
    53442 => -30034,
    53443 => -30033,
    53444 => -30032,
    53445 => -30031,
    53446 => -30029,
    53447 => -30028,
    53448 => -30027,
    53449 => -30026,
    53450 => -30024,
    53451 => -30023,
    53452 => -30022,
    53453 => -30020,
    53454 => -30019,
    53455 => -30018,
    53456 => -30017,
    53457 => -30015,
    53458 => -30014,
    53459 => -30013,
    53460 => -30012,
    53461 => -30010,
    53462 => -30009,
    53463 => -30008,
    53464 => -30007,
    53465 => -30005,
    53466 => -30004,
    53467 => -30003,
    53468 => -30002,
    53469 => -30000,
    53470 => -29999,
    53471 => -29998,
    53472 => -29997,
    53473 => -29995,
    53474 => -29994,
    53475 => -29993,
    53476 => -29991,
    53477 => -29990,
    53478 => -29989,
    53479 => -29988,
    53480 => -29986,
    53481 => -29985,
    53482 => -29984,
    53483 => -29983,
    53484 => -29981,
    53485 => -29980,
    53486 => -29979,
    53487 => -29978,
    53488 => -29976,
    53489 => -29975,
    53490 => -29974,
    53491 => -29972,
    53492 => -29971,
    53493 => -29970,
    53494 => -29969,
    53495 => -29967,
    53496 => -29966,
    53497 => -29965,
    53498 => -29964,
    53499 => -29962,
    53500 => -29961,
    53501 => -29960,
    53502 => -29958,
    53503 => -29957,
    53504 => -29956,
    53505 => -29955,
    53506 => -29953,
    53507 => -29952,
    53508 => -29951,
    53509 => -29950,
    53510 => -29948,
    53511 => -29947,
    53512 => -29946,
    53513 => -29944,
    53514 => -29943,
    53515 => -29942,
    53516 => -29941,
    53517 => -29939,
    53518 => -29938,
    53519 => -29937,
    53520 => -29936,
    53521 => -29934,
    53522 => -29933,
    53523 => -29932,
    53524 => -29930,
    53525 => -29929,
    53526 => -29928,
    53527 => -29927,
    53528 => -29925,
    53529 => -29924,
    53530 => -29923,
    53531 => -29921,
    53532 => -29920,
    53533 => -29919,
    53534 => -29918,
    53535 => -29916,
    53536 => -29915,
    53537 => -29914,
    53538 => -29912,
    53539 => -29911,
    53540 => -29910,
    53541 => -29909,
    53542 => -29907,
    53543 => -29906,
    53544 => -29905,
    53545 => -29903,
    53546 => -29902,
    53547 => -29901,
    53548 => -29900,
    53549 => -29898,
    53550 => -29897,
    53551 => -29896,
    53552 => -29894,
    53553 => -29893,
    53554 => -29892,
    53555 => -29891,
    53556 => -29889,
    53557 => -29888,
    53558 => -29887,
    53559 => -29885,
    53560 => -29884,
    53561 => -29883,
    53562 => -29882,
    53563 => -29880,
    53564 => -29879,
    53565 => -29878,
    53566 => -29876,
    53567 => -29875,
    53568 => -29874,
    53569 => -29873,
    53570 => -29871,
    53571 => -29870,
    53572 => -29869,
    53573 => -29867,
    53574 => -29866,
    53575 => -29865,
    53576 => -29864,
    53577 => -29862,
    53578 => -29861,
    53579 => -29860,
    53580 => -29858,
    53581 => -29857,
    53582 => -29856,
    53583 => -29854,
    53584 => -29853,
    53585 => -29852,
    53586 => -29851,
    53587 => -29849,
    53588 => -29848,
    53589 => -29847,
    53590 => -29845,
    53591 => -29844,
    53592 => -29843,
    53593 => -29842,
    53594 => -29840,
    53595 => -29839,
    53596 => -29838,
    53597 => -29836,
    53598 => -29835,
    53599 => -29834,
    53600 => -29832,
    53601 => -29831,
    53602 => -29830,
    53603 => -29829,
    53604 => -29827,
    53605 => -29826,
    53606 => -29825,
    53607 => -29823,
    53608 => -29822,
    53609 => -29821,
    53610 => -29819,
    53611 => -29818,
    53612 => -29817,
    53613 => -29816,
    53614 => -29814,
    53615 => -29813,
    53616 => -29812,
    53617 => -29810,
    53618 => -29809,
    53619 => -29808,
    53620 => -29806,
    53621 => -29805,
    53622 => -29804,
    53623 => -29802,
    53624 => -29801,
    53625 => -29800,
    53626 => -29799,
    53627 => -29797,
    53628 => -29796,
    53629 => -29795,
    53630 => -29793,
    53631 => -29792,
    53632 => -29791,
    53633 => -29789,
    53634 => -29788,
    53635 => -29787,
    53636 => -29785,
    53637 => -29784,
    53638 => -29783,
    53639 => -29782,
    53640 => -29780,
    53641 => -29779,
    53642 => -29778,
    53643 => -29776,
    53644 => -29775,
    53645 => -29774,
    53646 => -29772,
    53647 => -29771,
    53648 => -29770,
    53649 => -29768,
    53650 => -29767,
    53651 => -29766,
    53652 => -29764,
    53653 => -29763,
    53654 => -29762,
    53655 => -29761,
    53656 => -29759,
    53657 => -29758,
    53658 => -29757,
    53659 => -29755,
    53660 => -29754,
    53661 => -29753,
    53662 => -29751,
    53663 => -29750,
    53664 => -29749,
    53665 => -29747,
    53666 => -29746,
    53667 => -29745,
    53668 => -29743,
    53669 => -29742,
    53670 => -29741,
    53671 => -29739,
    53672 => -29738,
    53673 => -29737,
    53674 => -29736,
    53675 => -29734,
    53676 => -29733,
    53677 => -29732,
    53678 => -29730,
    53679 => -29729,
    53680 => -29728,
    53681 => -29726,
    53682 => -29725,
    53683 => -29724,
    53684 => -29722,
    53685 => -29721,
    53686 => -29720,
    53687 => -29718,
    53688 => -29717,
    53689 => -29716,
    53690 => -29714,
    53691 => -29713,
    53692 => -29712,
    53693 => -29710,
    53694 => -29709,
    53695 => -29708,
    53696 => -29706,
    53697 => -29705,
    53698 => -29704,
    53699 => -29702,
    53700 => -29701,
    53701 => -29700,
    53702 => -29698,
    53703 => -29697,
    53704 => -29696,
    53705 => -29694,
    53706 => -29693,
    53707 => -29692,
    53708 => -29690,
    53709 => -29689,
    53710 => -29688,
    53711 => -29687,
    53712 => -29685,
    53713 => -29684,
    53714 => -29683,
    53715 => -29681,
    53716 => -29680,
    53717 => -29679,
    53718 => -29677,
    53719 => -29676,
    53720 => -29675,
    53721 => -29673,
    53722 => -29672,
    53723 => -29671,
    53724 => -29669,
    53725 => -29668,
    53726 => -29667,
    53727 => -29665,
    53728 => -29664,
    53729 => -29663,
    53730 => -29661,
    53731 => -29660,
    53732 => -29659,
    53733 => -29657,
    53734 => -29656,
    53735 => -29655,
    53736 => -29653,
    53737 => -29652,
    53738 => -29651,
    53739 => -29649,
    53740 => -29648,
    53741 => -29646,
    53742 => -29645,
    53743 => -29644,
    53744 => -29642,
    53745 => -29641,
    53746 => -29640,
    53747 => -29638,
    53748 => -29637,
    53749 => -29636,
    53750 => -29634,
    53751 => -29633,
    53752 => -29632,
    53753 => -29630,
    53754 => -29629,
    53755 => -29628,
    53756 => -29626,
    53757 => -29625,
    53758 => -29624,
    53759 => -29622,
    53760 => -29621,
    53761 => -29620,
    53762 => -29618,
    53763 => -29617,
    53764 => -29616,
    53765 => -29614,
    53766 => -29613,
    53767 => -29612,
    53768 => -29610,
    53769 => -29609,
    53770 => -29608,
    53771 => -29606,
    53772 => -29605,
    53773 => -29604,
    53774 => -29602,
    53775 => -29601,
    53776 => -29599,
    53777 => -29598,
    53778 => -29597,
    53779 => -29595,
    53780 => -29594,
    53781 => -29593,
    53782 => -29591,
    53783 => -29590,
    53784 => -29589,
    53785 => -29587,
    53786 => -29586,
    53787 => -29585,
    53788 => -29583,
    53789 => -29582,
    53790 => -29581,
    53791 => -29579,
    53792 => -29578,
    53793 => -29577,
    53794 => -29575,
    53795 => -29574,
    53796 => -29572,
    53797 => -29571,
    53798 => -29570,
    53799 => -29568,
    53800 => -29567,
    53801 => -29566,
    53802 => -29564,
    53803 => -29563,
    53804 => -29562,
    53805 => -29560,
    53806 => -29559,
    53807 => -29558,
    53808 => -29556,
    53809 => -29555,
    53810 => -29554,
    53811 => -29552,
    53812 => -29551,
    53813 => -29549,
    53814 => -29548,
    53815 => -29547,
    53816 => -29545,
    53817 => -29544,
    53818 => -29543,
    53819 => -29541,
    53820 => -29540,
    53821 => -29539,
    53822 => -29537,
    53823 => -29536,
    53824 => -29534,
    53825 => -29533,
    53826 => -29532,
    53827 => -29530,
    53828 => -29529,
    53829 => -29528,
    53830 => -29526,
    53831 => -29525,
    53832 => -29524,
    53833 => -29522,
    53834 => -29521,
    53835 => -29520,
    53836 => -29518,
    53837 => -29517,
    53838 => -29515,
    53839 => -29514,
    53840 => -29513,
    53841 => -29511,
    53842 => -29510,
    53843 => -29509,
    53844 => -29507,
    53845 => -29506,
    53846 => -29504,
    53847 => -29503,
    53848 => -29502,
    53849 => -29500,
    53850 => -29499,
    53851 => -29498,
    53852 => -29496,
    53853 => -29495,
    53854 => -29494,
    53855 => -29492,
    53856 => -29491,
    53857 => -29489,
    53858 => -29488,
    53859 => -29487,
    53860 => -29485,
    53861 => -29484,
    53862 => -29483,
    53863 => -29481,
    53864 => -29480,
    53865 => -29478,
    53866 => -29477,
    53867 => -29476,
    53868 => -29474,
    53869 => -29473,
    53870 => -29472,
    53871 => -29470,
    53872 => -29469,
    53873 => -29468,
    53874 => -29466,
    53875 => -29465,
    53876 => -29463,
    53877 => -29462,
    53878 => -29461,
    53879 => -29459,
    53880 => -29458,
    53881 => -29457,
    53882 => -29455,
    53883 => -29454,
    53884 => -29452,
    53885 => -29451,
    53886 => -29450,
    53887 => -29448,
    53888 => -29447,
    53889 => -29445,
    53890 => -29444,
    53891 => -29443,
    53892 => -29441,
    53893 => -29440,
    53894 => -29439,
    53895 => -29437,
    53896 => -29436,
    53897 => -29434,
    53898 => -29433,
    53899 => -29432,
    53900 => -29430,
    53901 => -29429,
    53902 => -29428,
    53903 => -29426,
    53904 => -29425,
    53905 => -29423,
    53906 => -29422,
    53907 => -29421,
    53908 => -29419,
    53909 => -29418,
    53910 => -29416,
    53911 => -29415,
    53912 => -29414,
    53913 => -29412,
    53914 => -29411,
    53915 => -29410,
    53916 => -29408,
    53917 => -29407,
    53918 => -29405,
    53919 => -29404,
    53920 => -29403,
    53921 => -29401,
    53922 => -29400,
    53923 => -29398,
    53924 => -29397,
    53925 => -29396,
    53926 => -29394,
    53927 => -29393,
    53928 => -29392,
    53929 => -29390,
    53930 => -29389,
    53931 => -29387,
    53932 => -29386,
    53933 => -29385,
    53934 => -29383,
    53935 => -29382,
    53936 => -29380,
    53937 => -29379,
    53938 => -29378,
    53939 => -29376,
    53940 => -29375,
    53941 => -29373,
    53942 => -29372,
    53943 => -29371,
    53944 => -29369,
    53945 => -29368,
    53946 => -29366,
    53947 => -29365,
    53948 => -29364,
    53949 => -29362,
    53950 => -29361,
    53951 => -29360,
    53952 => -29358,
    53953 => -29357,
    53954 => -29355,
    53955 => -29354,
    53956 => -29353,
    53957 => -29351,
    53958 => -29350,
    53959 => -29348,
    53960 => -29347,
    53961 => -29346,
    53962 => -29344,
    53963 => -29343,
    53964 => -29341,
    53965 => -29340,
    53966 => -29339,
    53967 => -29337,
    53968 => -29336,
    53969 => -29334,
    53970 => -29333,
    53971 => -29332,
    53972 => -29330,
    53973 => -29329,
    53974 => -29327,
    53975 => -29326,
    53976 => -29325,
    53977 => -29323,
    53978 => -29322,
    53979 => -29320,
    53980 => -29319,
    53981 => -29318,
    53982 => -29316,
    53983 => -29315,
    53984 => -29313,
    53985 => -29312,
    53986 => -29311,
    53987 => -29309,
    53988 => -29308,
    53989 => -29306,
    53990 => -29305,
    53991 => -29304,
    53992 => -29302,
    53993 => -29301,
    53994 => -29299,
    53995 => -29298,
    53996 => -29296,
    53997 => -29295,
    53998 => -29294,
    53999 => -29292,
    54000 => -29291,
    54001 => -29289,
    54002 => -29288,
    54003 => -29287,
    54004 => -29285,
    54005 => -29284,
    54006 => -29282,
    54007 => -29281,
    54008 => -29280,
    54009 => -29278,
    54010 => -29277,
    54011 => -29275,
    54012 => -29274,
    54013 => -29273,
    54014 => -29271,
    54015 => -29270,
    54016 => -29268,
    54017 => -29267,
    54018 => -29265,
    54019 => -29264,
    54020 => -29263,
    54021 => -29261,
    54022 => -29260,
    54023 => -29258,
    54024 => -29257,
    54025 => -29256,
    54026 => -29254,
    54027 => -29253,
    54028 => -29251,
    54029 => -29250,
    54030 => -29248,
    54031 => -29247,
    54032 => -29246,
    54033 => -29244,
    54034 => -29243,
    54035 => -29241,
    54036 => -29240,
    54037 => -29239,
    54038 => -29237,
    54039 => -29236,
    54040 => -29234,
    54041 => -29233,
    54042 => -29231,
    54043 => -29230,
    54044 => -29229,
    54045 => -29227,
    54046 => -29226,
    54047 => -29224,
    54048 => -29223,
    54049 => -29222,
    54050 => -29220,
    54051 => -29219,
    54052 => -29217,
    54053 => -29216,
    54054 => -29214,
    54055 => -29213,
    54056 => -29212,
    54057 => -29210,
    54058 => -29209,
    54059 => -29207,
    54060 => -29206,
    54061 => -29204,
    54062 => -29203,
    54063 => -29202,
    54064 => -29200,
    54065 => -29199,
    54066 => -29197,
    54067 => -29196,
    54068 => -29194,
    54069 => -29193,
    54070 => -29192,
    54071 => -29190,
    54072 => -29189,
    54073 => -29187,
    54074 => -29186,
    54075 => -29184,
    54076 => -29183,
    54077 => -29182,
    54078 => -29180,
    54079 => -29179,
    54080 => -29177,
    54081 => -29176,
    54082 => -29174,
    54083 => -29173,
    54084 => -29172,
    54085 => -29170,
    54086 => -29169,
    54087 => -29167,
    54088 => -29166,
    54089 => -29164,
    54090 => -29163,
    54091 => -29162,
    54092 => -29160,
    54093 => -29159,
    54094 => -29157,
    54095 => -29156,
    54096 => -29154,
    54097 => -29153,
    54098 => -29152,
    54099 => -29150,
    54100 => -29149,
    54101 => -29147,
    54102 => -29146,
    54103 => -29144,
    54104 => -29143,
    54105 => -29142,
    54106 => -29140,
    54107 => -29139,
    54108 => -29137,
    54109 => -29136,
    54110 => -29134,
    54111 => -29133,
    54112 => -29131,
    54113 => -29130,
    54114 => -29129,
    54115 => -29127,
    54116 => -29126,
    54117 => -29124,
    54118 => -29123,
    54119 => -29121,
    54120 => -29120,
    54121 => -29118,
    54122 => -29117,
    54123 => -29116,
    54124 => -29114,
    54125 => -29113,
    54126 => -29111,
    54127 => -29110,
    54128 => -29108,
    54129 => -29107,
    54130 => -29106,
    54131 => -29104,
    54132 => -29103,
    54133 => -29101,
    54134 => -29100,
    54135 => -29098,
    54136 => -29097,
    54137 => -29095,
    54138 => -29094,
    54139 => -29093,
    54140 => -29091,
    54141 => -29090,
    54142 => -29088,
    54143 => -29087,
    54144 => -29085,
    54145 => -29084,
    54146 => -29082,
    54147 => -29081,
    54148 => -29079,
    54149 => -29078,
    54150 => -29077,
    54151 => -29075,
    54152 => -29074,
    54153 => -29072,
    54154 => -29071,
    54155 => -29069,
    54156 => -29068,
    54157 => -29066,
    54158 => -29065,
    54159 => -29064,
    54160 => -29062,
    54161 => -29061,
    54162 => -29059,
    54163 => -29058,
    54164 => -29056,
    54165 => -29055,
    54166 => -29053,
    54167 => -29052,
    54168 => -29050,
    54169 => -29049,
    54170 => -29048,
    54171 => -29046,
    54172 => -29045,
    54173 => -29043,
    54174 => -29042,
    54175 => -29040,
    54176 => -29039,
    54177 => -29037,
    54178 => -29036,
    54179 => -29034,
    54180 => -29033,
    54181 => -29032,
    54182 => -29030,
    54183 => -29029,
    54184 => -29027,
    54185 => -29026,
    54186 => -29024,
    54187 => -29023,
    54188 => -29021,
    54189 => -29020,
    54190 => -29018,
    54191 => -29017,
    54192 => -29016,
    54193 => -29014,
    54194 => -29013,
    54195 => -29011,
    54196 => -29010,
    54197 => -29008,
    54198 => -29007,
    54199 => -29005,
    54200 => -29004,
    54201 => -29002,
    54202 => -29001,
    54203 => -28999,
    54204 => -28998,
    54205 => -28997,
    54206 => -28995,
    54207 => -28994,
    54208 => -28992,
    54209 => -28991,
    54210 => -28989,
    54211 => -28988,
    54212 => -28986,
    54213 => -28985,
    54214 => -28983,
    54215 => -28982,
    54216 => -28980,
    54217 => -28979,
    54218 => -28977,
    54219 => -28976,
    54220 => -28975,
    54221 => -28973,
    54222 => -28972,
    54223 => -28970,
    54224 => -28969,
    54225 => -28967,
    54226 => -28966,
    54227 => -28964,
    54228 => -28963,
    54229 => -28961,
    54230 => -28960,
    54231 => -28958,
    54232 => -28957,
    54233 => -28955,
    54234 => -28954,
    54235 => -28953,
    54236 => -28951,
    54237 => -28950,
    54238 => -28948,
    54239 => -28947,
    54240 => -28945,
    54241 => -28944,
    54242 => -28942,
    54243 => -28941,
    54244 => -28939,
    54245 => -28938,
    54246 => -28936,
    54247 => -28935,
    54248 => -28933,
    54249 => -28932,
    54250 => -28930,
    54251 => -28929,
    54252 => -28927,
    54253 => -28926,
    54254 => -28925,
    54255 => -28923,
    54256 => -28922,
    54257 => -28920,
    54258 => -28919,
    54259 => -28917,
    54260 => -28916,
    54261 => -28914,
    54262 => -28913,
    54263 => -28911,
    54264 => -28910,
    54265 => -28908,
    54266 => -28907,
    54267 => -28905,
    54268 => -28904,
    54269 => -28902,
    54270 => -28901,
    54271 => -28899,
    54272 => -28898,
    54273 => -28896,
    54274 => -28895,
    54275 => -28893,
    54276 => -28892,
    54277 => -28891,
    54278 => -28889,
    54279 => -28888,
    54280 => -28886,
    54281 => -28885,
    54282 => -28883,
    54283 => -28882,
    54284 => -28880,
    54285 => -28879,
    54286 => -28877,
    54287 => -28876,
    54288 => -28874,
    54289 => -28873,
    54290 => -28871,
    54291 => -28870,
    54292 => -28868,
    54293 => -28867,
    54294 => -28865,
    54295 => -28864,
    54296 => -28862,
    54297 => -28861,
    54298 => -28859,
    54299 => -28858,
    54300 => -28856,
    54301 => -28855,
    54302 => -28853,
    54303 => -28852,
    54304 => -28850,
    54305 => -28849,
    54306 => -28847,
    54307 => -28846,
    54308 => -28844,
    54309 => -28843,
    54310 => -28841,
    54311 => -28840,
    54312 => -28838,
    54313 => -28837,
    54314 => -28835,
    54315 => -28834,
    54316 => -28832,
    54317 => -28831,
    54318 => -28830,
    54319 => -28828,
    54320 => -28827,
    54321 => -28825,
    54322 => -28824,
    54323 => -28822,
    54324 => -28821,
    54325 => -28819,
    54326 => -28818,
    54327 => -28816,
    54328 => -28815,
    54329 => -28813,
    54330 => -28812,
    54331 => -28810,
    54332 => -28809,
    54333 => -28807,
    54334 => -28806,
    54335 => -28804,
    54336 => -28803,
    54337 => -28801,
    54338 => -28800,
    54339 => -28798,
    54340 => -28797,
    54341 => -28795,
    54342 => -28794,
    54343 => -28792,
    54344 => -28791,
    54345 => -28789,
    54346 => -28788,
    54347 => -28786,
    54348 => -28785,
    54349 => -28783,
    54350 => -28782,
    54351 => -28780,
    54352 => -28779,
    54353 => -28777,
    54354 => -28776,
    54355 => -28774,
    54356 => -28773,
    54357 => -28771,
    54358 => -28770,
    54359 => -28768,
    54360 => -28767,
    54361 => -28765,
    54362 => -28764,
    54363 => -28762,
    54364 => -28761,
    54365 => -28759,
    54366 => -28758,
    54367 => -28756,
    54368 => -28755,
    54369 => -28753,
    54370 => -28752,
    54371 => -28750,
    54372 => -28748,
    54373 => -28747,
    54374 => -28745,
    54375 => -28744,
    54376 => -28742,
    54377 => -28741,
    54378 => -28739,
    54379 => -28738,
    54380 => -28736,
    54381 => -28735,
    54382 => -28733,
    54383 => -28732,
    54384 => -28730,
    54385 => -28729,
    54386 => -28727,
    54387 => -28726,
    54388 => -28724,
    54389 => -28723,
    54390 => -28721,
    54391 => -28720,
    54392 => -28718,
    54393 => -28717,
    54394 => -28715,
    54395 => -28714,
    54396 => -28712,
    54397 => -28711,
    54398 => -28709,
    54399 => -28708,
    54400 => -28706,
    54401 => -28705,
    54402 => -28703,
    54403 => -28702,
    54404 => -28700,
    54405 => -28699,
    54406 => -28697,
    54407 => -28696,
    54408 => -28694,
    54409 => -28693,
    54410 => -28691,
    54411 => -28690,
    54412 => -28688,
    54413 => -28686,
    54414 => -28685,
    54415 => -28683,
    54416 => -28682,
    54417 => -28680,
    54418 => -28679,
    54419 => -28677,
    54420 => -28676,
    54421 => -28674,
    54422 => -28673,
    54423 => -28671,
    54424 => -28670,
    54425 => -28668,
    54426 => -28667,
    54427 => -28665,
    54428 => -28664,
    54429 => -28662,
    54430 => -28661,
    54431 => -28659,
    54432 => -28658,
    54433 => -28656,
    54434 => -28655,
    54435 => -28653,
    54436 => -28651,
    54437 => -28650,
    54438 => -28648,
    54439 => -28647,
    54440 => -28645,
    54441 => -28644,
    54442 => -28642,
    54443 => -28641,
    54444 => -28639,
    54445 => -28638,
    54446 => -28636,
    54447 => -28635,
    54448 => -28633,
    54449 => -28632,
    54450 => -28630,
    54451 => -28629,
    54452 => -28627,
    54453 => -28626,
    54454 => -28624,
    54455 => -28622,
    54456 => -28621,
    54457 => -28619,
    54458 => -28618,
    54459 => -28616,
    54460 => -28615,
    54461 => -28613,
    54462 => -28612,
    54463 => -28610,
    54464 => -28609,
    54465 => -28607,
    54466 => -28606,
    54467 => -28604,
    54468 => -28603,
    54469 => -28601,
    54470 => -28600,
    54471 => -28598,
    54472 => -28596,
    54473 => -28595,
    54474 => -28593,
    54475 => -28592,
    54476 => -28590,
    54477 => -28589,
    54478 => -28587,
    54479 => -28586,
    54480 => -28584,
    54481 => -28583,
    54482 => -28581,
    54483 => -28580,
    54484 => -28578,
    54485 => -28576,
    54486 => -28575,
    54487 => -28573,
    54488 => -28572,
    54489 => -28570,
    54490 => -28569,
    54491 => -28567,
    54492 => -28566,
    54493 => -28564,
    54494 => -28563,
    54495 => -28561,
    54496 => -28560,
    54497 => -28558,
    54498 => -28556,
    54499 => -28555,
    54500 => -28553,
    54501 => -28552,
    54502 => -28550,
    54503 => -28549,
    54504 => -28547,
    54505 => -28546,
    54506 => -28544,
    54507 => -28543,
    54508 => -28541,
    54509 => -28540,
    54510 => -28538,
    54511 => -28536,
    54512 => -28535,
    54513 => -28533,
    54514 => -28532,
    54515 => -28530,
    54516 => -28529,
    54517 => -28527,
    54518 => -28526,
    54519 => -28524,
    54520 => -28523,
    54521 => -28521,
    54522 => -28519,
    54523 => -28518,
    54524 => -28516,
    54525 => -28515,
    54526 => -28513,
    54527 => -28512,
    54528 => -28510,
    54529 => -28509,
    54530 => -28507,
    54531 => -28505,
    54532 => -28504,
    54533 => -28502,
    54534 => -28501,
    54535 => -28499,
    54536 => -28498,
    54537 => -28496,
    54538 => -28495,
    54539 => -28493,
    54540 => -28492,
    54541 => -28490,
    54542 => -28488,
    54543 => -28487,
    54544 => -28485,
    54545 => -28484,
    54546 => -28482,
    54547 => -28481,
    54548 => -28479,
    54549 => -28478,
    54550 => -28476,
    54551 => -28474,
    54552 => -28473,
    54553 => -28471,
    54554 => -28470,
    54555 => -28468,
    54556 => -28467,
    54557 => -28465,
    54558 => -28464,
    54559 => -28462,
    54560 => -28460,
    54561 => -28459,
    54562 => -28457,
    54563 => -28456,
    54564 => -28454,
    54565 => -28453,
    54566 => -28451,
    54567 => -28450,
    54568 => -28448,
    54569 => -28446,
    54570 => -28445,
    54571 => -28443,
    54572 => -28442,
    54573 => -28440,
    54574 => -28439,
    54575 => -28437,
    54576 => -28436,
    54577 => -28434,
    54578 => -28432,
    54579 => -28431,
    54580 => -28429,
    54581 => -28428,
    54582 => -28426,
    54583 => -28425,
    54584 => -28423,
    54585 => -28421,
    54586 => -28420,
    54587 => -28418,
    54588 => -28417,
    54589 => -28415,
    54590 => -28414,
    54591 => -28412,
    54592 => -28411,
    54593 => -28409,
    54594 => -28407,
    54595 => -28406,
    54596 => -28404,
    54597 => -28403,
    54598 => -28401,
    54599 => -28400,
    54600 => -28398,
    54601 => -28396,
    54602 => -28395,
    54603 => -28393,
    54604 => -28392,
    54605 => -28390,
    54606 => -28389,
    54607 => -28387,
    54608 => -28385,
    54609 => -28384,
    54610 => -28382,
    54611 => -28381,
    54612 => -28379,
    54613 => -28378,
    54614 => -28376,
    54615 => -28374,
    54616 => -28373,
    54617 => -28371,
    54618 => -28370,
    54619 => -28368,
    54620 => -28367,
    54621 => -28365,
    54622 => -28363,
    54623 => -28362,
    54624 => -28360,
    54625 => -28359,
    54626 => -28357,
    54627 => -28356,
    54628 => -28354,
    54629 => -28352,
    54630 => -28351,
    54631 => -28349,
    54632 => -28348,
    54633 => -28346,
    54634 => -28345,
    54635 => -28343,
    54636 => -28341,
    54637 => -28340,
    54638 => -28338,
    54639 => -28337,
    54640 => -28335,
    54641 => -28333,
    54642 => -28332,
    54643 => -28330,
    54644 => -28329,
    54645 => -28327,
    54646 => -28326,
    54647 => -28324,
    54648 => -28322,
    54649 => -28321,
    54650 => -28319,
    54651 => -28318,
    54652 => -28316,
    54653 => -28315,
    54654 => -28313,
    54655 => -28311,
    54656 => -28310,
    54657 => -28308,
    54658 => -28307,
    54659 => -28305,
    54660 => -28303,
    54661 => -28302,
    54662 => -28300,
    54663 => -28299,
    54664 => -28297,
    54665 => -28296,
    54666 => -28294,
    54667 => -28292,
    54668 => -28291,
    54669 => -28289,
    54670 => -28288,
    54671 => -28286,
    54672 => -28284,
    54673 => -28283,
    54674 => -28281,
    54675 => -28280,
    54676 => -28278,
    54677 => -28277,
    54678 => -28275,
    54679 => -28273,
    54680 => -28272,
    54681 => -28270,
    54682 => -28269,
    54683 => -28267,
    54684 => -28265,
    54685 => -28264,
    54686 => -28262,
    54687 => -28261,
    54688 => -28259,
    54689 => -28257,
    54690 => -28256,
    54691 => -28254,
    54692 => -28253,
    54693 => -28251,
    54694 => -28249,
    54695 => -28248,
    54696 => -28246,
    54697 => -28245,
    54698 => -28243,
    54699 => -28242,
    54700 => -28240,
    54701 => -28238,
    54702 => -28237,
    54703 => -28235,
    54704 => -28234,
    54705 => -28232,
    54706 => -28230,
    54707 => -28229,
    54708 => -28227,
    54709 => -28226,
    54710 => -28224,
    54711 => -28222,
    54712 => -28221,
    54713 => -28219,
    54714 => -28218,
    54715 => -28216,
    54716 => -28214,
    54717 => -28213,
    54718 => -28211,
    54719 => -28210,
    54720 => -28208,
    54721 => -28206,
    54722 => -28205,
    54723 => -28203,
    54724 => -28202,
    54725 => -28200,
    54726 => -28198,
    54727 => -28197,
    54728 => -28195,
    54729 => -28194,
    54730 => -28192,
    54731 => -28190,
    54732 => -28189,
    54733 => -28187,
    54734 => -28186,
    54735 => -28184,
    54736 => -28182,
    54737 => -28181,
    54738 => -28179,
    54739 => -28178,
    54740 => -28176,
    54741 => -28174,
    54742 => -28173,
    54743 => -28171,
    54744 => -28170,
    54745 => -28168,
    54746 => -28166,
    54747 => -28165,
    54748 => -28163,
    54749 => -28162,
    54750 => -28160,
    54751 => -28158,
    54752 => -28157,
    54753 => -28155,
    54754 => -28154,
    54755 => -28152,
    54756 => -28150,
    54757 => -28149,
    54758 => -28147,
    54759 => -28145,
    54760 => -28144,
    54761 => -28142,
    54762 => -28141,
    54763 => -28139,
    54764 => -28137,
    54765 => -28136,
    54766 => -28134,
    54767 => -28133,
    54768 => -28131,
    54769 => -28129,
    54770 => -28128,
    54771 => -28126,
    54772 => -28125,
    54773 => -28123,
    54774 => -28121,
    54775 => -28120,
    54776 => -28118,
    54777 => -28116,
    54778 => -28115,
    54779 => -28113,
    54780 => -28112,
    54781 => -28110,
    54782 => -28108,
    54783 => -28107,
    54784 => -28105,
    54785 => -28104,
    54786 => -28102,
    54787 => -28100,
    54788 => -28099,
    54789 => -28097,
    54790 => -28095,
    54791 => -28094,
    54792 => -28092,
    54793 => -28091,
    54794 => -28089,
    54795 => -28087,
    54796 => -28086,
    54797 => -28084,
    54798 => -28083,
    54799 => -28081,
    54800 => -28079,
    54801 => -28078,
    54802 => -28076,
    54803 => -28074,
    54804 => -28073,
    54805 => -28071,
    54806 => -28070,
    54807 => -28068,
    54808 => -28066,
    54809 => -28065,
    54810 => -28063,
    54811 => -28061,
    54812 => -28060,
    54813 => -28058,
    54814 => -28057,
    54815 => -28055,
    54816 => -28053,
    54817 => -28052,
    54818 => -28050,
    54819 => -28049,
    54820 => -28047,
    54821 => -28045,
    54822 => -28044,
    54823 => -28042,
    54824 => -28040,
    54825 => -28039,
    54826 => -28037,
    54827 => -28036,
    54828 => -28034,
    54829 => -28032,
    54830 => -28031,
    54831 => -28029,
    54832 => -28027,
    54833 => -28026,
    54834 => -28024,
    54835 => -28022,
    54836 => -28021,
    54837 => -28019,
    54838 => -28018,
    54839 => -28016,
    54840 => -28014,
    54841 => -28013,
    54842 => -28011,
    54843 => -28009,
    54844 => -28008,
    54845 => -28006,
    54846 => -28005,
    54847 => -28003,
    54848 => -28001,
    54849 => -28000,
    54850 => -27998,
    54851 => -27996,
    54852 => -27995,
    54853 => -27993,
    54854 => -27992,
    54855 => -27990,
    54856 => -27988,
    54857 => -27987,
    54858 => -27985,
    54859 => -27983,
    54860 => -27982,
    54861 => -27980,
    54862 => -27978,
    54863 => -27977,
    54864 => -27975,
    54865 => -27974,
    54866 => -27972,
    54867 => -27970,
    54868 => -27969,
    54869 => -27967,
    54870 => -27965,
    54871 => -27964,
    54872 => -27962,
    54873 => -27960,
    54874 => -27959,
    54875 => -27957,
    54876 => -27956,
    54877 => -27954,
    54878 => -27952,
    54879 => -27951,
    54880 => -27949,
    54881 => -27947,
    54882 => -27946,
    54883 => -27944,
    54884 => -27942,
    54885 => -27941,
    54886 => -27939,
    54887 => -27937,
    54888 => -27936,
    54889 => -27934,
    54890 => -27933,
    54891 => -27931,
    54892 => -27929,
    54893 => -27928,
    54894 => -27926,
    54895 => -27924,
    54896 => -27923,
    54897 => -27921,
    54898 => -27919,
    54899 => -27918,
    54900 => -27916,
    54901 => -27914,
    54902 => -27913,
    54903 => -27911,
    54904 => -27910,
    54905 => -27908,
    54906 => -27906,
    54907 => -27905,
    54908 => -27903,
    54909 => -27901,
    54910 => -27900,
    54911 => -27898,
    54912 => -27896,
    54913 => -27895,
    54914 => -27893,
    54915 => -27891,
    54916 => -27890,
    54917 => -27888,
    54918 => -27886,
    54919 => -27885,
    54920 => -27883,
    54921 => -27882,
    54922 => -27880,
    54923 => -27878,
    54924 => -27877,
    54925 => -27875,
    54926 => -27873,
    54927 => -27872,
    54928 => -27870,
    54929 => -27868,
    54930 => -27867,
    54931 => -27865,
    54932 => -27863,
    54933 => -27862,
    54934 => -27860,
    54935 => -27858,
    54936 => -27857,
    54937 => -27855,
    54938 => -27853,
    54939 => -27852,
    54940 => -27850,
    54941 => -27848,
    54942 => -27847,
    54943 => -27845,
    54944 => -27843,
    54945 => -27842,
    54946 => -27840,
    54947 => -27839,
    54948 => -27837,
    54949 => -27835,
    54950 => -27834,
    54951 => -27832,
    54952 => -27830,
    54953 => -27829,
    54954 => -27827,
    54955 => -27825,
    54956 => -27824,
    54957 => -27822,
    54958 => -27820,
    54959 => -27819,
    54960 => -27817,
    54961 => -27815,
    54962 => -27814,
    54963 => -27812,
    54964 => -27810,
    54965 => -27809,
    54966 => -27807,
    54967 => -27805,
    54968 => -27804,
    54969 => -27802,
    54970 => -27800,
    54971 => -27799,
    54972 => -27797,
    54973 => -27795,
    54974 => -27794,
    54975 => -27792,
    54976 => -27790,
    54977 => -27789,
    54978 => -27787,
    54979 => -27785,
    54980 => -27784,
    54981 => -27782,
    54982 => -27780,
    54983 => -27779,
    54984 => -27777,
    54985 => -27775,
    54986 => -27774,
    54987 => -27772,
    54988 => -27770,
    54989 => -27769,
    54990 => -27767,
    54991 => -27765,
    54992 => -27764,
    54993 => -27762,
    54994 => -27760,
    54995 => -27759,
    54996 => -27757,
    54997 => -27755,
    54998 => -27754,
    54999 => -27752,
    55000 => -27750,
    55001 => -27749,
    55002 => -27747,
    55003 => -27745,
    55004 => -27744,
    55005 => -27742,
    55006 => -27740,
    55007 => -27739,
    55008 => -27737,
    55009 => -27735,
    55010 => -27734,
    55011 => -27732,
    55012 => -27730,
    55013 => -27729,
    55014 => -27727,
    55015 => -27725,
    55016 => -27724,
    55017 => -27722,
    55018 => -27720,
    55019 => -27719,
    55020 => -27717,
    55021 => -27715,
    55022 => -27714,
    55023 => -27712,
    55024 => -27710,
    55025 => -27708,
    55026 => -27707,
    55027 => -27705,
    55028 => -27703,
    55029 => -27702,
    55030 => -27700,
    55031 => -27698,
    55032 => -27697,
    55033 => -27695,
    55034 => -27693,
    55035 => -27692,
    55036 => -27690,
    55037 => -27688,
    55038 => -27687,
    55039 => -27685,
    55040 => -27683,
    55041 => -27682,
    55042 => -27680,
    55043 => -27678,
    55044 => -27677,
    55045 => -27675,
    55046 => -27673,
    55047 => -27672,
    55048 => -27670,
    55049 => -27668,
    55050 => -27666,
    55051 => -27665,
    55052 => -27663,
    55053 => -27661,
    55054 => -27660,
    55055 => -27658,
    55056 => -27656,
    55057 => -27655,
    55058 => -27653,
    55059 => -27651,
    55060 => -27650,
    55061 => -27648,
    55062 => -27646,
    55063 => -27645,
    55064 => -27643,
    55065 => -27641,
    55066 => -27640,
    55067 => -27638,
    55068 => -27636,
    55069 => -27634,
    55070 => -27633,
    55071 => -27631,
    55072 => -27629,
    55073 => -27628,
    55074 => -27626,
    55075 => -27624,
    55076 => -27623,
    55077 => -27621,
    55078 => -27619,
    55079 => -27618,
    55080 => -27616,
    55081 => -27614,
    55082 => -27613,
    55083 => -27611,
    55084 => -27609,
    55085 => -27607,
    55086 => -27606,
    55087 => -27604,
    55088 => -27602,
    55089 => -27601,
    55090 => -27599,
    55091 => -27597,
    55092 => -27596,
    55093 => -27594,
    55094 => -27592,
    55095 => -27590,
    55096 => -27589,
    55097 => -27587,
    55098 => -27585,
    55099 => -27584,
    55100 => -27582,
    55101 => -27580,
    55102 => -27579,
    55103 => -27577,
    55104 => -27575,
    55105 => -27574,
    55106 => -27572,
    55107 => -27570,
    55108 => -27568,
    55109 => -27567,
    55110 => -27565,
    55111 => -27563,
    55112 => -27562,
    55113 => -27560,
    55114 => -27558,
    55115 => -27557,
    55116 => -27555,
    55117 => -27553,
    55118 => -27551,
    55119 => -27550,
    55120 => -27548,
    55121 => -27546,
    55122 => -27545,
    55123 => -27543,
    55124 => -27541,
    55125 => -27540,
    55126 => -27538,
    55127 => -27536,
    55128 => -27534,
    55129 => -27533,
    55130 => -27531,
    55131 => -27529,
    55132 => -27528,
    55133 => -27526,
    55134 => -27524,
    55135 => -27523,
    55136 => -27521,
    55137 => -27519,
    55138 => -27517,
    55139 => -27516,
    55140 => -27514,
    55141 => -27512,
    55142 => -27511,
    55143 => -27509,
    55144 => -27507,
    55145 => -27505,
    55146 => -27504,
    55147 => -27502,
    55148 => -27500,
    55149 => -27499,
    55150 => -27497,
    55151 => -27495,
    55152 => -27493,
    55153 => -27492,
    55154 => -27490,
    55155 => -27488,
    55156 => -27487,
    55157 => -27485,
    55158 => -27483,
    55159 => -27482,
    55160 => -27480,
    55161 => -27478,
    55162 => -27476,
    55163 => -27475,
    55164 => -27473,
    55165 => -27471,
    55166 => -27470,
    55167 => -27468,
    55168 => -27466,
    55169 => -27464,
    55170 => -27463,
    55171 => -27461,
    55172 => -27459,
    55173 => -27458,
    55174 => -27456,
    55175 => -27454,
    55176 => -27452,
    55177 => -27451,
    55178 => -27449,
    55179 => -27447,
    55180 => -27446,
    55181 => -27444,
    55182 => -27442,
    55183 => -27440,
    55184 => -27439,
    55185 => -27437,
    55186 => -27435,
    55187 => -27434,
    55188 => -27432,
    55189 => -27430,
    55190 => -27428,
    55191 => -27427,
    55192 => -27425,
    55193 => -27423,
    55194 => -27421,
    55195 => -27420,
    55196 => -27418,
    55197 => -27416,
    55198 => -27415,
    55199 => -27413,
    55200 => -27411,
    55201 => -27409,
    55202 => -27408,
    55203 => -27406,
    55204 => -27404,
    55205 => -27403,
    55206 => -27401,
    55207 => -27399,
    55208 => -27397,
    55209 => -27396,
    55210 => -27394,
    55211 => -27392,
    55212 => -27390,
    55213 => -27389,
    55214 => -27387,
    55215 => -27385,
    55216 => -27384,
    55217 => -27382,
    55218 => -27380,
    55219 => -27378,
    55220 => -27377,
    55221 => -27375,
    55222 => -27373,
    55223 => -27372,
    55224 => -27370,
    55225 => -27368,
    55226 => -27366,
    55227 => -27365,
    55228 => -27363,
    55229 => -27361,
    55230 => -27359,
    55231 => -27358,
    55232 => -27356,
    55233 => -27354,
    55234 => -27352,
    55235 => -27351,
    55236 => -27349,
    55237 => -27347,
    55238 => -27346,
    55239 => -27344,
    55240 => -27342,
    55241 => -27340,
    55242 => -27339,
    55243 => -27337,
    55244 => -27335,
    55245 => -27333,
    55246 => -27332,
    55247 => -27330,
    55248 => -27328,
    55249 => -27327,
    55250 => -27325,
    55251 => -27323,
    55252 => -27321,
    55253 => -27320,
    55254 => -27318,
    55255 => -27316,
    55256 => -27314,
    55257 => -27313,
    55258 => -27311,
    55259 => -27309,
    55260 => -27307,
    55261 => -27306,
    55262 => -27304,
    55263 => -27302,
    55264 => -27300,
    55265 => -27299,
    55266 => -27297,
    55267 => -27295,
    55268 => -27294,
    55269 => -27292,
    55270 => -27290,
    55271 => -27288,
    55272 => -27287,
    55273 => -27285,
    55274 => -27283,
    55275 => -27281,
    55276 => -27280,
    55277 => -27278,
    55278 => -27276,
    55279 => -27274,
    55280 => -27273,
    55281 => -27271,
    55282 => -27269,
    55283 => -27267,
    55284 => -27266,
    55285 => -27264,
    55286 => -27262,
    55287 => -27260,
    55288 => -27259,
    55289 => -27257,
    55290 => -27255,
    55291 => -27253,
    55292 => -27252,
    55293 => -27250,
    55294 => -27248,
    55295 => -27247,
    55296 => -27245,
    55297 => -27243,
    55298 => -27241,
    55299 => -27240,
    55300 => -27238,
    55301 => -27236,
    55302 => -27234,
    55303 => -27233,
    55304 => -27231,
    55305 => -27229,
    55306 => -27227,
    55307 => -27226,
    55308 => -27224,
    55309 => -27222,
    55310 => -27220,
    55311 => -27219,
    55312 => -27217,
    55313 => -27215,
    55314 => -27213,
    55315 => -27212,
    55316 => -27210,
    55317 => -27208,
    55318 => -27206,
    55319 => -27205,
    55320 => -27203,
    55321 => -27201,
    55322 => -27199,
    55323 => -27198,
    55324 => -27196,
    55325 => -27194,
    55326 => -27192,
    55327 => -27191,
    55328 => -27189,
    55329 => -27187,
    55330 => -27185,
    55331 => -27184,
    55332 => -27182,
    55333 => -27180,
    55334 => -27178,
    55335 => -27177,
    55336 => -27175,
    55337 => -27173,
    55338 => -27171,
    55339 => -27169,
    55340 => -27168,
    55341 => -27166,
    55342 => -27164,
    55343 => -27162,
    55344 => -27161,
    55345 => -27159,
    55346 => -27157,
    55347 => -27155,
    55348 => -27154,
    55349 => -27152,
    55350 => -27150,
    55351 => -27148,
    55352 => -27147,
    55353 => -27145,
    55354 => -27143,
    55355 => -27141,
    55356 => -27140,
    55357 => -27138,
    55358 => -27136,
    55359 => -27134,
    55360 => -27133,
    55361 => -27131,
    55362 => -27129,
    55363 => -27127,
    55364 => -27126,
    55365 => -27124,
    55366 => -27122,
    55367 => -27120,
    55368 => -27118,
    55369 => -27117,
    55370 => -27115,
    55371 => -27113,
    55372 => -27111,
    55373 => -27110,
    55374 => -27108,
    55375 => -27106,
    55376 => -27104,
    55377 => -27103,
    55378 => -27101,
    55379 => -27099,
    55380 => -27097,
    55381 => -27096,
    55382 => -27094,
    55383 => -27092,
    55384 => -27090,
    55385 => -27088,
    55386 => -27087,
    55387 => -27085,
    55388 => -27083,
    55389 => -27081,
    55390 => -27080,
    55391 => -27078,
    55392 => -27076,
    55393 => -27074,
    55394 => -27073,
    55395 => -27071,
    55396 => -27069,
    55397 => -27067,
    55398 => -27065,
    55399 => -27064,
    55400 => -27062,
    55401 => -27060,
    55402 => -27058,
    55403 => -27057,
    55404 => -27055,
    55405 => -27053,
    55406 => -27051,
    55407 => -27049,
    55408 => -27048,
    55409 => -27046,
    55410 => -27044,
    55411 => -27042,
    55412 => -27041,
    55413 => -27039,
    55414 => -27037,
    55415 => -27035,
    55416 => -27034,
    55417 => -27032,
    55418 => -27030,
    55419 => -27028,
    55420 => -27026,
    55421 => -27025,
    55422 => -27023,
    55423 => -27021,
    55424 => -27019,
    55425 => -27018,
    55426 => -27016,
    55427 => -27014,
    55428 => -27012,
    55429 => -27010,
    55430 => -27009,
    55431 => -27007,
    55432 => -27005,
    55433 => -27003,
    55434 => -27002,
    55435 => -27000,
    55436 => -26998,
    55437 => -26996,
    55438 => -26994,
    55439 => -26993,
    55440 => -26991,
    55441 => -26989,
    55442 => -26987,
    55443 => -26986,
    55444 => -26984,
    55445 => -26982,
    55446 => -26980,
    55447 => -26978,
    55448 => -26977,
    55449 => -26975,
    55450 => -26973,
    55451 => -26971,
    55452 => -26969,
    55453 => -26968,
    55454 => -26966,
    55455 => -26964,
    55456 => -26962,
    55457 => -26961,
    55458 => -26959,
    55459 => -26957,
    55460 => -26955,
    55461 => -26953,
    55462 => -26952,
    55463 => -26950,
    55464 => -26948,
    55465 => -26946,
    55466 => -26944,
    55467 => -26943,
    55468 => -26941,
    55469 => -26939,
    55470 => -26937,
    55471 => -26936,
    55472 => -26934,
    55473 => -26932,
    55474 => -26930,
    55475 => -26928,
    55476 => -26927,
    55477 => -26925,
    55478 => -26923,
    55479 => -26921,
    55480 => -26919,
    55481 => -26918,
    55482 => -26916,
    55483 => -26914,
    55484 => -26912,
    55485 => -26910,
    55486 => -26909,
    55487 => -26907,
    55488 => -26905,
    55489 => -26903,
    55490 => -26901,
    55491 => -26900,
    55492 => -26898,
    55493 => -26896,
    55494 => -26894,
    55495 => -26893,
    55496 => -26891,
    55497 => -26889,
    55498 => -26887,
    55499 => -26885,
    55500 => -26884,
    55501 => -26882,
    55502 => -26880,
    55503 => -26878,
    55504 => -26876,
    55505 => -26875,
    55506 => -26873,
    55507 => -26871,
    55508 => -26869,
    55509 => -26867,
    55510 => -26866,
    55511 => -26864,
    55512 => -26862,
    55513 => -26860,
    55514 => -26858,
    55515 => -26857,
    55516 => -26855,
    55517 => -26853,
    55518 => -26851,
    55519 => -26849,
    55520 => -26848,
    55521 => -26846,
    55522 => -26844,
    55523 => -26842,
    55524 => -26840,
    55525 => -26839,
    55526 => -26837,
    55527 => -26835,
    55528 => -26833,
    55529 => -26831,
    55530 => -26830,
    55531 => -26828,
    55532 => -26826,
    55533 => -26824,
    55534 => -26822,
    55535 => -26821,
    55536 => -26819,
    55537 => -26817,
    55538 => -26815,
    55539 => -26813,
    55540 => -26811,
    55541 => -26810,
    55542 => -26808,
    55543 => -26806,
    55544 => -26804,
    55545 => -26802,
    55546 => -26801,
    55547 => -26799,
    55548 => -26797,
    55549 => -26795,
    55550 => -26793,
    55551 => -26792,
    55552 => -26790,
    55553 => -26788,
    55554 => -26786,
    55555 => -26784,
    55556 => -26783,
    55557 => -26781,
    55558 => -26779,
    55559 => -26777,
    55560 => -26775,
    55561 => -26774,
    55562 => -26772,
    55563 => -26770,
    55564 => -26768,
    55565 => -26766,
    55566 => -26764,
    55567 => -26763,
    55568 => -26761,
    55569 => -26759,
    55570 => -26757,
    55571 => -26755,
    55572 => -26754,
    55573 => -26752,
    55574 => -26750,
    55575 => -26748,
    55576 => -26746,
    55577 => -26745,
    55578 => -26743,
    55579 => -26741,
    55580 => -26739,
    55581 => -26737,
    55582 => -26735,
    55583 => -26734,
    55584 => -26732,
    55585 => -26730,
    55586 => -26728,
    55587 => -26726,
    55588 => -26725,
    55589 => -26723,
    55590 => -26721,
    55591 => -26719,
    55592 => -26717,
    55593 => -26715,
    55594 => -26714,
    55595 => -26712,
    55596 => -26710,
    55597 => -26708,
    55598 => -26706,
    55599 => -26705,
    55600 => -26703,
    55601 => -26701,
    55602 => -26699,
    55603 => -26697,
    55604 => -26695,
    55605 => -26694,
    55606 => -26692,
    55607 => -26690,
    55608 => -26688,
    55609 => -26686,
    55610 => -26684,
    55611 => -26683,
    55612 => -26681,
    55613 => -26679,
    55614 => -26677,
    55615 => -26675,
    55616 => -26674,
    55617 => -26672,
    55618 => -26670,
    55619 => -26668,
    55620 => -26666,
    55621 => -26664,
    55622 => -26663,
    55623 => -26661,
    55624 => -26659,
    55625 => -26657,
    55626 => -26655,
    55627 => -26653,
    55628 => -26652,
    55629 => -26650,
    55630 => -26648,
    55631 => -26646,
    55632 => -26644,
    55633 => -26642,
    55634 => -26641,
    55635 => -26639,
    55636 => -26637,
    55637 => -26635,
    55638 => -26633,
    55639 => -26631,
    55640 => -26630,
    55641 => -26628,
    55642 => -26626,
    55643 => -26624,
    55644 => -26622,
    55645 => -26621,
    55646 => -26619,
    55647 => -26617,
    55648 => -26615,
    55649 => -26613,
    55650 => -26611,
    55651 => -26610,
    55652 => -26608,
    55653 => -26606,
    55654 => -26604,
    55655 => -26602,
    55656 => -26600,
    55657 => -26599,
    55658 => -26597,
    55659 => -26595,
    55660 => -26593,
    55661 => -26591,
    55662 => -26589,
    55663 => -26588,
    55664 => -26586,
    55665 => -26584,
    55666 => -26582,
    55667 => -26580,
    55668 => -26578,
    55669 => -26576,
    55670 => -26575,
    55671 => -26573,
    55672 => -26571,
    55673 => -26569,
    55674 => -26567,
    55675 => -26565,
    55676 => -26564,
    55677 => -26562,
    55678 => -26560,
    55679 => -26558,
    55680 => -26556,
    55681 => -26554,
    55682 => -26553,
    55683 => -26551,
    55684 => -26549,
    55685 => -26547,
    55686 => -26545,
    55687 => -26543,
    55688 => -26542,
    55689 => -26540,
    55690 => -26538,
    55691 => -26536,
    55692 => -26534,
    55693 => -26532,
    55694 => -26530,
    55695 => -26529,
    55696 => -26527,
    55697 => -26525,
    55698 => -26523,
    55699 => -26521,
    55700 => -26519,
    55701 => -26518,
    55702 => -26516,
    55703 => -26514,
    55704 => -26512,
    55705 => -26510,
    55706 => -26508,
    55707 => -26506,
    55708 => -26505,
    55709 => -26503,
    55710 => -26501,
    55711 => -26499,
    55712 => -26497,
    55713 => -26495,
    55714 => -26494,
    55715 => -26492,
    55716 => -26490,
    55717 => -26488,
    55718 => -26486,
    55719 => -26484,
    55720 => -26482,
    55721 => -26481,
    55722 => -26479,
    55723 => -26477,
    55724 => -26475,
    55725 => -26473,
    55726 => -26471,
    55727 => -26469,
    55728 => -26468,
    55729 => -26466,
    55730 => -26464,
    55731 => -26462,
    55732 => -26460,
    55733 => -26458,
    55734 => -26457,
    55735 => -26455,
    55736 => -26453,
    55737 => -26451,
    55738 => -26449,
    55739 => -26447,
    55740 => -26445,
    55741 => -26444,
    55742 => -26442,
    55743 => -26440,
    55744 => -26438,
    55745 => -26436,
    55746 => -26434,
    55747 => -26432,
    55748 => -26431,
    55749 => -26429,
    55750 => -26427,
    55751 => -26425,
    55752 => -26423,
    55753 => -26421,
    55754 => -26419,
    55755 => -26418,
    55756 => -26416,
    55757 => -26414,
    55758 => -26412,
    55759 => -26410,
    55760 => -26408,
    55761 => -26406,
    55762 => -26405,
    55763 => -26403,
    55764 => -26401,
    55765 => -26399,
    55766 => -26397,
    55767 => -26395,
    55768 => -26393,
    55769 => -26392,
    55770 => -26390,
    55771 => -26388,
    55772 => -26386,
    55773 => -26384,
    55774 => -26382,
    55775 => -26380,
    55776 => -26378,
    55777 => -26377,
    55778 => -26375,
    55779 => -26373,
    55780 => -26371,
    55781 => -26369,
    55782 => -26367,
    55783 => -26365,
    55784 => -26364,
    55785 => -26362,
    55786 => -26360,
    55787 => -26358,
    55788 => -26356,
    55789 => -26354,
    55790 => -26352,
    55791 => -26350,
    55792 => -26349,
    55793 => -26347,
    55794 => -26345,
    55795 => -26343,
    55796 => -26341,
    55797 => -26339,
    55798 => -26337,
    55799 => -26336,
    55800 => -26334,
    55801 => -26332,
    55802 => -26330,
    55803 => -26328,
    55804 => -26326,
    55805 => -26324,
    55806 => -26322,
    55807 => -26321,
    55808 => -26319,
    55809 => -26317,
    55810 => -26315,
    55811 => -26313,
    55812 => -26311,
    55813 => -26309,
    55814 => -26307,
    55815 => -26306,
    55816 => -26304,
    55817 => -26302,
    55818 => -26300,
    55819 => -26298,
    55820 => -26296,
    55821 => -26294,
    55822 => -26292,
    55823 => -26291,
    55824 => -26289,
    55825 => -26287,
    55826 => -26285,
    55827 => -26283,
    55828 => -26281,
    55829 => -26279,
    55830 => -26277,
    55831 => -26276,
    55832 => -26274,
    55833 => -26272,
    55834 => -26270,
    55835 => -26268,
    55836 => -26266,
    55837 => -26264,
    55838 => -26262,
    55839 => -26261,
    55840 => -26259,
    55841 => -26257,
    55842 => -26255,
    55843 => -26253,
    55844 => -26251,
    55845 => -26249,
    55846 => -26247,
    55847 => -26246,
    55848 => -26244,
    55849 => -26242,
    55850 => -26240,
    55851 => -26238,
    55852 => -26236,
    55853 => -26234,
    55854 => -26232,
    55855 => -26230,
    55856 => -26229,
    55857 => -26227,
    55858 => -26225,
    55859 => -26223,
    55860 => -26221,
    55861 => -26219,
    55862 => -26217,
    55863 => -26215,
    55864 => -26214,
    55865 => -26212,
    55866 => -26210,
    55867 => -26208,
    55868 => -26206,
    55869 => -26204,
    55870 => -26202,
    55871 => -26200,
    55872 => -26198,
    55873 => -26197,
    55874 => -26195,
    55875 => -26193,
    55876 => -26191,
    55877 => -26189,
    55878 => -26187,
    55879 => -26185,
    55880 => -26183,
    55881 => -26181,
    55882 => -26180,
    55883 => -26178,
    55884 => -26176,
    55885 => -26174,
    55886 => -26172,
    55887 => -26170,
    55888 => -26168,
    55889 => -26166,
    55890 => -26164,
    55891 => -26163,
    55892 => -26161,
    55893 => -26159,
    55894 => -26157,
    55895 => -26155,
    55896 => -26153,
    55897 => -26151,
    55898 => -26149,
    55899 => -26147,
    55900 => -26146,
    55901 => -26144,
    55902 => -26142,
    55903 => -26140,
    55904 => -26138,
    55905 => -26136,
    55906 => -26134,
    55907 => -26132,
    55908 => -26130,
    55909 => -26128,
    55910 => -26127,
    55911 => -26125,
    55912 => -26123,
    55913 => -26121,
    55914 => -26119,
    55915 => -26117,
    55916 => -26115,
    55917 => -26113,
    55918 => -26111,
    55919 => -26109,
    55920 => -26108,
    55921 => -26106,
    55922 => -26104,
    55923 => -26102,
    55924 => -26100,
    55925 => -26098,
    55926 => -26096,
    55927 => -26094,
    55928 => -26092,
    55929 => -26090,
    55930 => -26089,
    55931 => -26087,
    55932 => -26085,
    55933 => -26083,
    55934 => -26081,
    55935 => -26079,
    55936 => -26077,
    55937 => -26075,
    55938 => -26073,
    55939 => -26071,
    55940 => -26070,
    55941 => -26068,
    55942 => -26066,
    55943 => -26064,
    55944 => -26062,
    55945 => -26060,
    55946 => -26058,
    55947 => -26056,
    55948 => -26054,
    55949 => -26052,
    55950 => -26051,
    55951 => -26049,
    55952 => -26047,
    55953 => -26045,
    55954 => -26043,
    55955 => -26041,
    55956 => -26039,
    55957 => -26037,
    55958 => -26035,
    55959 => -26033,
    55960 => -26031,
    55961 => -26030,
    55962 => -26028,
    55963 => -26026,
    55964 => -26024,
    55965 => -26022,
    55966 => -26020,
    55967 => -26018,
    55968 => -26016,
    55969 => -26014,
    55970 => -26012,
    55971 => -26010,
    55972 => -26009,
    55973 => -26007,
    55974 => -26005,
    55975 => -26003,
    55976 => -26001,
    55977 => -25999,
    55978 => -25997,
    55979 => -25995,
    55980 => -25993,
    55981 => -25991,
    55982 => -25989,
    55983 => -25988,
    55984 => -25986,
    55985 => -25984,
    55986 => -25982,
    55987 => -25980,
    55988 => -25978,
    55989 => -25976,
    55990 => -25974,
    55991 => -25972,
    55992 => -25970,
    55993 => -25968,
    55994 => -25966,
    55995 => -25965,
    55996 => -25963,
    55997 => -25961,
    55998 => -25959,
    55999 => -25957,
    56000 => -25955,
    56001 => -25953,
    56002 => -25951,
    56003 => -25949,
    56004 => -25947,
    56005 => -25945,
    56006 => -25943,
    56007 => -25942,
    56008 => -25940,
    56009 => -25938,
    56010 => -25936,
    56011 => -25934,
    56012 => -25932,
    56013 => -25930,
    56014 => -25928,
    56015 => -25926,
    56016 => -25924,
    56017 => -25922,
    56018 => -25920,
    56019 => -25918,
    56020 => -25917,
    56021 => -25915,
    56022 => -25913,
    56023 => -25911,
    56024 => -25909,
    56025 => -25907,
    56026 => -25905,
    56027 => -25903,
    56028 => -25901,
    56029 => -25899,
    56030 => -25897,
    56031 => -25895,
    56032 => -25893,
    56033 => -25892,
    56034 => -25890,
    56035 => -25888,
    56036 => -25886,
    56037 => -25884,
    56038 => -25882,
    56039 => -25880,
    56040 => -25878,
    56041 => -25876,
    56042 => -25874,
    56043 => -25872,
    56044 => -25870,
    56045 => -25868,
    56046 => -25866,
    56047 => -25865,
    56048 => -25863,
    56049 => -25861,
    56050 => -25859,
    56051 => -25857,
    56052 => -25855,
    56053 => -25853,
    56054 => -25851,
    56055 => -25849,
    56056 => -25847,
    56057 => -25845,
    56058 => -25843,
    56059 => -25841,
    56060 => -25839,
    56061 => -25838,
    56062 => -25836,
    56063 => -25834,
    56064 => -25832,
    56065 => -25830,
    56066 => -25828,
    56067 => -25826,
    56068 => -25824,
    56069 => -25822,
    56070 => -25820,
    56071 => -25818,
    56072 => -25816,
    56073 => -25814,
    56074 => -25812,
    56075 => -25810,
    56076 => -25809,
    56077 => -25807,
    56078 => -25805,
    56079 => -25803,
    56080 => -25801,
    56081 => -25799,
    56082 => -25797,
    56083 => -25795,
    56084 => -25793,
    56085 => -25791,
    56086 => -25789,
    56087 => -25787,
    56088 => -25785,
    56089 => -25783,
    56090 => -25781,
    56091 => -25779,
    56092 => -25778,
    56093 => -25776,
    56094 => -25774,
    56095 => -25772,
    56096 => -25770,
    56097 => -25768,
    56098 => -25766,
    56099 => -25764,
    56100 => -25762,
    56101 => -25760,
    56102 => -25758,
    56103 => -25756,
    56104 => -25754,
    56105 => -25752,
    56106 => -25750,
    56107 => -25748,
    56108 => -25746,
    56109 => -25745,
    56110 => -25743,
    56111 => -25741,
    56112 => -25739,
    56113 => -25737,
    56114 => -25735,
    56115 => -25733,
    56116 => -25731,
    56117 => -25729,
    56118 => -25727,
    56119 => -25725,
    56120 => -25723,
    56121 => -25721,
    56122 => -25719,
    56123 => -25717,
    56124 => -25715,
    56125 => -25713,
    56126 => -25711,
    56127 => -25710,
    56128 => -25708,
    56129 => -25706,
    56130 => -25704,
    56131 => -25702,
    56132 => -25700,
    56133 => -25698,
    56134 => -25696,
    56135 => -25694,
    56136 => -25692,
    56137 => -25690,
    56138 => -25688,
    56139 => -25686,
    56140 => -25684,
    56141 => -25682,
    56142 => -25680,
    56143 => -25678,
    56144 => -25676,
    56145 => -25674,
    56146 => -25672,
    56147 => -25671,
    56148 => -25669,
    56149 => -25667,
    56150 => -25665,
    56151 => -25663,
    56152 => -25661,
    56153 => -25659,
    56154 => -25657,
    56155 => -25655,
    56156 => -25653,
    56157 => -25651,
    56158 => -25649,
    56159 => -25647,
    56160 => -25645,
    56161 => -25643,
    56162 => -25641,
    56163 => -25639,
    56164 => -25637,
    56165 => -25635,
    56166 => -25633,
    56167 => -25631,
    56168 => -25629,
    56169 => -25628,
    56170 => -25626,
    56171 => -25624,
    56172 => -25622,
    56173 => -25620,
    56174 => -25618,
    56175 => -25616,
    56176 => -25614,
    56177 => -25612,
    56178 => -25610,
    56179 => -25608,
    56180 => -25606,
    56181 => -25604,
    56182 => -25602,
    56183 => -25600,
    56184 => -25598,
    56185 => -25596,
    56186 => -25594,
    56187 => -25592,
    56188 => -25590,
    56189 => -25588,
    56190 => -25586,
    56191 => -25584,
    56192 => -25582,
    56193 => -25580,
    56194 => -25578,
    56195 => -25577,
    56196 => -25575,
    56197 => -25573,
    56198 => -25571,
    56199 => -25569,
    56200 => -25567,
    56201 => -25565,
    56202 => -25563,
    56203 => -25561,
    56204 => -25559,
    56205 => -25557,
    56206 => -25555,
    56207 => -25553,
    56208 => -25551,
    56209 => -25549,
    56210 => -25547,
    56211 => -25545,
    56212 => -25543,
    56213 => -25541,
    56214 => -25539,
    56215 => -25537,
    56216 => -25535,
    56217 => -25533,
    56218 => -25531,
    56219 => -25529,
    56220 => -25527,
    56221 => -25525,
    56222 => -25523,
    56223 => -25521,
    56224 => -25519,
    56225 => -25518,
    56226 => -25516,
    56227 => -25514,
    56228 => -25512,
    56229 => -25510,
    56230 => -25508,
    56231 => -25506,
    56232 => -25504,
    56233 => -25502,
    56234 => -25500,
    56235 => -25498,
    56236 => -25496,
    56237 => -25494,
    56238 => -25492,
    56239 => -25490,
    56240 => -25488,
    56241 => -25486,
    56242 => -25484,
    56243 => -25482,
    56244 => -25480,
    56245 => -25478,
    56246 => -25476,
    56247 => -25474,
    56248 => -25472,
    56249 => -25470,
    56250 => -25468,
    56251 => -25466,
    56252 => -25464,
    56253 => -25462,
    56254 => -25460,
    56255 => -25458,
    56256 => -25456,
    56257 => -25454,
    56258 => -25452,
    56259 => -25450,
    56260 => -25448,
    56261 => -25446,
    56262 => -25444,
    56263 => -25442,
    56264 => -25440,
    56265 => -25438,
    56266 => -25437,
    56267 => -25435,
    56268 => -25433,
    56269 => -25431,
    56270 => -25429,
    56271 => -25427,
    56272 => -25425,
    56273 => -25423,
    56274 => -25421,
    56275 => -25419,
    56276 => -25417,
    56277 => -25415,
    56278 => -25413,
    56279 => -25411,
    56280 => -25409,
    56281 => -25407,
    56282 => -25405,
    56283 => -25403,
    56284 => -25401,
    56285 => -25399,
    56286 => -25397,
    56287 => -25395,
    56288 => -25393,
    56289 => -25391,
    56290 => -25389,
    56291 => -25387,
    56292 => -25385,
    56293 => -25383,
    56294 => -25381,
    56295 => -25379,
    56296 => -25377,
    56297 => -25375,
    56298 => -25373,
    56299 => -25371,
    56300 => -25369,
    56301 => -25367,
    56302 => -25365,
    56303 => -25363,
    56304 => -25361,
    56305 => -25359,
    56306 => -25357,
    56307 => -25355,
    56308 => -25353,
    56309 => -25351,
    56310 => -25349,
    56311 => -25347,
    56312 => -25345,
    56313 => -25343,
    56314 => -25341,
    56315 => -25339,
    56316 => -25337,
    56317 => -25335,
    56318 => -25333,
    56319 => -25331,
    56320 => -25329,
    56321 => -25327,
    56322 => -25325,
    56323 => -25323,
    56324 => -25321,
    56325 => -25319,
    56326 => -25317,
    56327 => -25315,
    56328 => -25313,
    56329 => -25311,
    56330 => -25309,
    56331 => -25307,
    56332 => -25305,
    56333 => -25303,
    56334 => -25301,
    56335 => -25299,
    56336 => -25297,
    56337 => -25295,
    56338 => -25293,
    56339 => -25291,
    56340 => -25289,
    56341 => -25287,
    56342 => -25285,
    56343 => -25283,
    56344 => -25281,
    56345 => -25279,
    56346 => -25277,
    56347 => -25275,
    56348 => -25273,
    56349 => -25271,
    56350 => -25269,
    56351 => -25267,
    56352 => -25265,
    56353 => -25263,
    56354 => -25261,
    56355 => -25259,
    56356 => -25257,
    56357 => -25255,
    56358 => -25253,
    56359 => -25251,
    56360 => -25249,
    56361 => -25247,
    56362 => -25245,
    56363 => -25243,
    56364 => -25241,
    56365 => -25239,
    56366 => -25237,
    56367 => -25235,
    56368 => -25233,
    56369 => -25231,
    56370 => -25229,
    56371 => -25227,
    56372 => -25225,
    56373 => -25223,
    56374 => -25221,
    56375 => -25219,
    56376 => -25217,
    56377 => -25215,
    56378 => -25213,
    56379 => -25211,
    56380 => -25209,
    56381 => -25207,
    56382 => -25205,
    56383 => -25203,
    56384 => -25201,
    56385 => -25199,
    56386 => -25197,
    56387 => -25195,
    56388 => -25193,
    56389 => -25191,
    56390 => -25189,
    56391 => -25187,
    56392 => -25185,
    56393 => -25183,
    56394 => -25181,
    56395 => -25179,
    56396 => -25177,
    56397 => -25175,
    56398 => -25173,
    56399 => -25171,
    56400 => -25169,
    56401 => -25167,
    56402 => -25165,
    56403 => -25163,
    56404 => -25161,
    56405 => -25159,
    56406 => -25157,
    56407 => -25155,
    56408 => -25153,
    56409 => -25151,
    56410 => -25149,
    56411 => -25147,
    56412 => -25145,
    56413 => -25143,
    56414 => -25141,
    56415 => -25139,
    56416 => -25137,
    56417 => -25135,
    56418 => -25133,
    56419 => -25131,
    56420 => -25129,
    56421 => -25127,
    56422 => -25125,
    56423 => -25123,
    56424 => -25121,
    56425 => -25119,
    56426 => -25117,
    56427 => -25115,
    56428 => -25113,
    56429 => -25111,
    56430 => -25109,
    56431 => -25107,
    56432 => -25105,
    56433 => -25103,
    56434 => -25101,
    56435 => -25099,
    56436 => -25096,
    56437 => -25094,
    56438 => -25092,
    56439 => -25090,
    56440 => -25088,
    56441 => -25086,
    56442 => -25084,
    56443 => -25082,
    56444 => -25080,
    56445 => -25078,
    56446 => -25076,
    56447 => -25074,
    56448 => -25072,
    56449 => -25070,
    56450 => -25068,
    56451 => -25066,
    56452 => -25064,
    56453 => -25062,
    56454 => -25060,
    56455 => -25058,
    56456 => -25056,
    56457 => -25054,
    56458 => -25052,
    56459 => -25050,
    56460 => -25048,
    56461 => -25046,
    56462 => -25044,
    56463 => -25042,
    56464 => -25040,
    56465 => -25038,
    56466 => -25036,
    56467 => -25034,
    56468 => -25032,
    56469 => -25030,
    56470 => -25028,
    56471 => -25026,
    56472 => -25024,
    56473 => -25022,
    56474 => -25020,
    56475 => -25018,
    56476 => -25016,
    56477 => -25013,
    56478 => -25011,
    56479 => -25009,
    56480 => -25007,
    56481 => -25005,
    56482 => -25003,
    56483 => -25001,
    56484 => -24999,
    56485 => -24997,
    56486 => -24995,
    56487 => -24993,
    56488 => -24991,
    56489 => -24989,
    56490 => -24987,
    56491 => -24985,
    56492 => -24983,
    56493 => -24981,
    56494 => -24979,
    56495 => -24977,
    56496 => -24975,
    56497 => -24973,
    56498 => -24971,
    56499 => -24969,
    56500 => -24967,
    56501 => -24965,
    56502 => -24963,
    56503 => -24961,
    56504 => -24959,
    56505 => -24957,
    56506 => -24955,
    56507 => -24953,
    56508 => -24950,
    56509 => -24948,
    56510 => -24946,
    56511 => -24944,
    56512 => -24942,
    56513 => -24940,
    56514 => -24938,
    56515 => -24936,
    56516 => -24934,
    56517 => -24932,
    56518 => -24930,
    56519 => -24928,
    56520 => -24926,
    56521 => -24924,
    56522 => -24922,
    56523 => -24920,
    56524 => -24918,
    56525 => -24916,
    56526 => -24914,
    56527 => -24912,
    56528 => -24910,
    56529 => -24908,
    56530 => -24906,
    56531 => -24904,
    56532 => -24902,
    56533 => -24899,
    56534 => -24897,
    56535 => -24895,
    56536 => -24893,
    56537 => -24891,
    56538 => -24889,
    56539 => -24887,
    56540 => -24885,
    56541 => -24883,
    56542 => -24881,
    56543 => -24879,
    56544 => -24877,
    56545 => -24875,
    56546 => -24873,
    56547 => -24871,
    56548 => -24869,
    56549 => -24867,
    56550 => -24865,
    56551 => -24863,
    56552 => -24861,
    56553 => -24859,
    56554 => -24857,
    56555 => -24855,
    56556 => -24852,
    56557 => -24850,
    56558 => -24848,
    56559 => -24846,
    56560 => -24844,
    56561 => -24842,
    56562 => -24840,
    56563 => -24838,
    56564 => -24836,
    56565 => -24834,
    56566 => -24832,
    56567 => -24830,
    56568 => -24828,
    56569 => -24826,
    56570 => -24824,
    56571 => -24822,
    56572 => -24820,
    56573 => -24818,
    56574 => -24816,
    56575 => -24814,
    56576 => -24811,
    56577 => -24809,
    56578 => -24807,
    56579 => -24805,
    56580 => -24803,
    56581 => -24801,
    56582 => -24799,
    56583 => -24797,
    56584 => -24795,
    56585 => -24793,
    56586 => -24791,
    56587 => -24789,
    56588 => -24787,
    56589 => -24785,
    56590 => -24783,
    56591 => -24781,
    56592 => -24779,
    56593 => -24777,
    56594 => -24774,
    56595 => -24772,
    56596 => -24770,
    56597 => -24768,
    56598 => -24766,
    56599 => -24764,
    56600 => -24762,
    56601 => -24760,
    56602 => -24758,
    56603 => -24756,
    56604 => -24754,
    56605 => -24752,
    56606 => -24750,
    56607 => -24748,
    56608 => -24746,
    56609 => -24744,
    56610 => -24742,
    56611 => -24740,
    56612 => -24737,
    56613 => -24735,
    56614 => -24733,
    56615 => -24731,
    56616 => -24729,
    56617 => -24727,
    56618 => -24725,
    56619 => -24723,
    56620 => -24721,
    56621 => -24719,
    56622 => -24717,
    56623 => -24715,
    56624 => -24713,
    56625 => -24711,
    56626 => -24709,
    56627 => -24707,
    56628 => -24704,
    56629 => -24702,
    56630 => -24700,
    56631 => -24698,
    56632 => -24696,
    56633 => -24694,
    56634 => -24692,
    56635 => -24690,
    56636 => -24688,
    56637 => -24686,
    56638 => -24684,
    56639 => -24682,
    56640 => -24680,
    56641 => -24678,
    56642 => -24676,
    56643 => -24673,
    56644 => -24671,
    56645 => -24669,
    56646 => -24667,
    56647 => -24665,
    56648 => -24663,
    56649 => -24661,
    56650 => -24659,
    56651 => -24657,
    56652 => -24655,
    56653 => -24653,
    56654 => -24651,
    56655 => -24649,
    56656 => -24647,
    56657 => -24645,
    56658 => -24642,
    56659 => -24640,
    56660 => -24638,
    56661 => -24636,
    56662 => -24634,
    56663 => -24632,
    56664 => -24630,
    56665 => -24628,
    56666 => -24626,
    56667 => -24624,
    56668 => -24622,
    56669 => -24620,
    56670 => -24618,
    56671 => -24616,
    56672 => -24613,
    56673 => -24611,
    56674 => -24609,
    56675 => -24607,
    56676 => -24605,
    56677 => -24603,
    56678 => -24601,
    56679 => -24599,
    56680 => -24597,
    56681 => -24595,
    56682 => -24593,
    56683 => -24591,
    56684 => -24589,
    56685 => -24586,
    56686 => -24584,
    56687 => -24582,
    56688 => -24580,
    56689 => -24578,
    56690 => -24576,
    56691 => -24574,
    56692 => -24572,
    56693 => -24570,
    56694 => -24568,
    56695 => -24566,
    56696 => -24564,
    56697 => -24562,
    56698 => -24559,
    56699 => -24557,
    56700 => -24555,
    56701 => -24553,
    56702 => -24551,
    56703 => -24549,
    56704 => -24547,
    56705 => -24545,
    56706 => -24543,
    56707 => -24541,
    56708 => -24539,
    56709 => -24537,
    56710 => -24534,
    56711 => -24532,
    56712 => -24530,
    56713 => -24528,
    56714 => -24526,
    56715 => -24524,
    56716 => -24522,
    56717 => -24520,
    56718 => -24518,
    56719 => -24516,
    56720 => -24514,
    56721 => -24512,
    56722 => -24509,
    56723 => -24507,
    56724 => -24505,
    56725 => -24503,
    56726 => -24501,
    56727 => -24499,
    56728 => -24497,
    56729 => -24495,
    56730 => -24493,
    56731 => -24491,
    56732 => -24489,
    56733 => -24487,
    56734 => -24484,
    56735 => -24482,
    56736 => -24480,
    56737 => -24478,
    56738 => -24476,
    56739 => -24474,
    56740 => -24472,
    56741 => -24470,
    56742 => -24468,
    56743 => -24466,
    56744 => -24464,
    56745 => -24461,
    56746 => -24459,
    56747 => -24457,
    56748 => -24455,
    56749 => -24453,
    56750 => -24451,
    56751 => -24449,
    56752 => -24447,
    56753 => -24445,
    56754 => -24443,
    56755 => -24441,
    56756 => -24438,
    56757 => -24436,
    56758 => -24434,
    56759 => -24432,
    56760 => -24430,
    56761 => -24428,
    56762 => -24426,
    56763 => -24424,
    56764 => -24422,
    56765 => -24420,
    56766 => -24417,
    56767 => -24415,
    56768 => -24413,
    56769 => -24411,
    56770 => -24409,
    56771 => -24407,
    56772 => -24405,
    56773 => -24403,
    56774 => -24401,
    56775 => -24399,
    56776 => -24397,
    56777 => -24394,
    56778 => -24392,
    56779 => -24390,
    56780 => -24388,
    56781 => -24386,
    56782 => -24384,
    56783 => -24382,
    56784 => -24380,
    56785 => -24378,
    56786 => -24376,
    56787 => -24373,
    56788 => -24371,
    56789 => -24369,
    56790 => -24367,
    56791 => -24365,
    56792 => -24363,
    56793 => -24361,
    56794 => -24359,
    56795 => -24357,
    56796 => -24355,
    56797 => -24352,
    56798 => -24350,
    56799 => -24348,
    56800 => -24346,
    56801 => -24344,
    56802 => -24342,
    56803 => -24340,
    56804 => -24338,
    56805 => -24336,
    56806 => -24334,
    56807 => -24331,
    56808 => -24329,
    56809 => -24327,
    56810 => -24325,
    56811 => -24323,
    56812 => -24321,
    56813 => -24319,
    56814 => -24317,
    56815 => -24315,
    56816 => -24312,
    56817 => -24310,
    56818 => -24308,
    56819 => -24306,
    56820 => -24304,
    56821 => -24302,
    56822 => -24300,
    56823 => -24298,
    56824 => -24296,
    56825 => -24294,
    56826 => -24291,
    56827 => -24289,
    56828 => -24287,
    56829 => -24285,
    56830 => -24283,
    56831 => -24281,
    56832 => -24279,
    56833 => -24277,
    56834 => -24275,
    56835 => -24272,
    56836 => -24270,
    56837 => -24268,
    56838 => -24266,
    56839 => -24264,
    56840 => -24262,
    56841 => -24260,
    56842 => -24258,
    56843 => -24256,
    56844 => -24253,
    56845 => -24251,
    56846 => -24249,
    56847 => -24247,
    56848 => -24245,
    56849 => -24243,
    56850 => -24241,
    56851 => -24239,
    56852 => -24237,
    56853 => -24234,
    56854 => -24232,
    56855 => -24230,
    56856 => -24228,
    56857 => -24226,
    56858 => -24224,
    56859 => -24222,
    56860 => -24220,
    56861 => -24217,
    56862 => -24215,
    56863 => -24213,
    56864 => -24211,
    56865 => -24209,
    56866 => -24207,
    56867 => -24205,
    56868 => -24203,
    56869 => -24201,
    56870 => -24198,
    56871 => -24196,
    56872 => -24194,
    56873 => -24192,
    56874 => -24190,
    56875 => -24188,
    56876 => -24186,
    56877 => -24184,
    56878 => -24181,
    56879 => -24179,
    56880 => -24177,
    56881 => -24175,
    56882 => -24173,
    56883 => -24171,
    56884 => -24169,
    56885 => -24167,
    56886 => -24164,
    56887 => -24162,
    56888 => -24160,
    56889 => -24158,
    56890 => -24156,
    56891 => -24154,
    56892 => -24152,
    56893 => -24150,
    56894 => -24148,
    56895 => -24145,
    56896 => -24143,
    56897 => -24141,
    56898 => -24139,
    56899 => -24137,
    56900 => -24135,
    56901 => -24133,
    56902 => -24131,
    56903 => -24128,
    56904 => -24126,
    56905 => -24124,
    56906 => -24122,
    56907 => -24120,
    56908 => -24118,
    56909 => -24116,
    56910 => -24114,
    56911 => -24111,
    56912 => -24109,
    56913 => -24107,
    56914 => -24105,
    56915 => -24103,
    56916 => -24101,
    56917 => -24099,
    56918 => -24096,
    56919 => -24094,
    56920 => -24092,
    56921 => -24090,
    56922 => -24088,
    56923 => -24086,
    56924 => -24084,
    56925 => -24082,
    56926 => -24079,
    56927 => -24077,
    56928 => -24075,
    56929 => -24073,
    56930 => -24071,
    56931 => -24069,
    56932 => -24067,
    56933 => -24065,
    56934 => -24062,
    56935 => -24060,
    56936 => -24058,
    56937 => -24056,
    56938 => -24054,
    56939 => -24052,
    56940 => -24050,
    56941 => -24047,
    56942 => -24045,
    56943 => -24043,
    56944 => -24041,
    56945 => -24039,
    56946 => -24037,
    56947 => -24035,
    56948 => -24033,
    56949 => -24030,
    56950 => -24028,
    56951 => -24026,
    56952 => -24024,
    56953 => -24022,
    56954 => -24020,
    56955 => -24018,
    56956 => -24015,
    56957 => -24013,
    56958 => -24011,
    56959 => -24009,
    56960 => -24007,
    56961 => -24005,
    56962 => -24003,
    56963 => -24000,
    56964 => -23998,
    56965 => -23996,
    56966 => -23994,
    56967 => -23992,
    56968 => -23990,
    56969 => -23988,
    56970 => -23985,
    56971 => -23983,
    56972 => -23981,
    56973 => -23979,
    56974 => -23977,
    56975 => -23975,
    56976 => -23973,
    56977 => -23971,
    56978 => -23968,
    56979 => -23966,
    56980 => -23964,
    56981 => -23962,
    56982 => -23960,
    56983 => -23958,
    56984 => -23956,
    56985 => -23953,
    56986 => -23951,
    56987 => -23949,
    56988 => -23947,
    56989 => -23945,
    56990 => -23943,
    56991 => -23940,
    56992 => -23938,
    56993 => -23936,
    56994 => -23934,
    56995 => -23932,
    56996 => -23930,
    56997 => -23928,
    56998 => -23925,
    56999 => -23923,
    57000 => -23921,
    57001 => -23919,
    57002 => -23917,
    57003 => -23915,
    57004 => -23913,
    57005 => -23910,
    57006 => -23908,
    57007 => -23906,
    57008 => -23904,
    57009 => -23902,
    57010 => -23900,
    57011 => -23898,
    57012 => -23895,
    57013 => -23893,
    57014 => -23891,
    57015 => -23889,
    57016 => -23887,
    57017 => -23885,
    57018 => -23883,
    57019 => -23880,
    57020 => -23878,
    57021 => -23876,
    57022 => -23874,
    57023 => -23872,
    57024 => -23870,
    57025 => -23867,
    57026 => -23865,
    57027 => -23863,
    57028 => -23861,
    57029 => -23859,
    57030 => -23857,
    57031 => -23855,
    57032 => -23852,
    57033 => -23850,
    57034 => -23848,
    57035 => -23846,
    57036 => -23844,
    57037 => -23842,
    57038 => -23839,
    57039 => -23837,
    57040 => -23835,
    57041 => -23833,
    57042 => -23831,
    57043 => -23829,
    57044 => -23827,
    57045 => -23824,
    57046 => -23822,
    57047 => -23820,
    57048 => -23818,
    57049 => -23816,
    57050 => -23814,
    57051 => -23811,
    57052 => -23809,
    57053 => -23807,
    57054 => -23805,
    57055 => -23803,
    57056 => -23801,
    57057 => -23798,
    57058 => -23796,
    57059 => -23794,
    57060 => -23792,
    57061 => -23790,
    57062 => -23788,
    57063 => -23785,
    57064 => -23783,
    57065 => -23781,
    57066 => -23779,
    57067 => -23777,
    57068 => -23775,
    57069 => -23773,
    57070 => -23770,
    57071 => -23768,
    57072 => -23766,
    57073 => -23764,
    57074 => -23762,
    57075 => -23760,
    57076 => -23757,
    57077 => -23755,
    57078 => -23753,
    57079 => -23751,
    57080 => -23749,
    57081 => -23747,
    57082 => -23744,
    57083 => -23742,
    57084 => -23740,
    57085 => -23738,
    57086 => -23736,
    57087 => -23734,
    57088 => -23731,
    57089 => -23729,
    57090 => -23727,
    57091 => -23725,
    57092 => -23723,
    57093 => -23721,
    57094 => -23718,
    57095 => -23716,
    57096 => -23714,
    57097 => -23712,
    57098 => -23710,
    57099 => -23708,
    57100 => -23705,
    57101 => -23703,
    57102 => -23701,
    57103 => -23699,
    57104 => -23697,
    57105 => -23695,
    57106 => -23692,
    57107 => -23690,
    57108 => -23688,
    57109 => -23686,
    57110 => -23684,
    57111 => -23682,
    57112 => -23679,
    57113 => -23677,
    57114 => -23675,
    57115 => -23673,
    57116 => -23671,
    57117 => -23668,
    57118 => -23666,
    57119 => -23664,
    57120 => -23662,
    57121 => -23660,
    57122 => -23658,
    57123 => -23655,
    57124 => -23653,
    57125 => -23651,
    57126 => -23649,
    57127 => -23647,
    57128 => -23645,
    57129 => -23642,
    57130 => -23640,
    57131 => -23638,
    57132 => -23636,
    57133 => -23634,
    57134 => -23632,
    57135 => -23629,
    57136 => -23627,
    57137 => -23625,
    57138 => -23623,
    57139 => -23621,
    57140 => -23618,
    57141 => -23616,
    57142 => -23614,
    57143 => -23612,
    57144 => -23610,
    57145 => -23608,
    57146 => -23605,
    57147 => -23603,
    57148 => -23601,
    57149 => -23599,
    57150 => -23597,
    57151 => -23595,
    57152 => -23592,
    57153 => -23590,
    57154 => -23588,
    57155 => -23586,
    57156 => -23584,
    57157 => -23581,
    57158 => -23579,
    57159 => -23577,
    57160 => -23575,
    57161 => -23573,
    57162 => -23571,
    57163 => -23568,
    57164 => -23566,
    57165 => -23564,
    57166 => -23562,
    57167 => -23560,
    57168 => -23557,
    57169 => -23555,
    57170 => -23553,
    57171 => -23551,
    57172 => -23549,
    57173 => -23546,
    57174 => -23544,
    57175 => -23542,
    57176 => -23540,
    57177 => -23538,
    57178 => -23536,
    57179 => -23533,
    57180 => -23531,
    57181 => -23529,
    57182 => -23527,
    57183 => -23525,
    57184 => -23522,
    57185 => -23520,
    57186 => -23518,
    57187 => -23516,
    57188 => -23514,
    57189 => -23512,
    57190 => -23509,
    57191 => -23507,
    57192 => -23505,
    57193 => -23503,
    57194 => -23501,
    57195 => -23498,
    57196 => -23496,
    57197 => -23494,
    57198 => -23492,
    57199 => -23490,
    57200 => -23487,
    57201 => -23485,
    57202 => -23483,
    57203 => -23481,
    57204 => -23479,
    57205 => -23476,
    57206 => -23474,
    57207 => -23472,
    57208 => -23470,
    57209 => -23468,
    57210 => -23466,
    57211 => -23463,
    57212 => -23461,
    57213 => -23459,
    57214 => -23457,
    57215 => -23455,
    57216 => -23452,
    57217 => -23450,
    57218 => -23448,
    57219 => -23446,
    57220 => -23444,
    57221 => -23441,
    57222 => -23439,
    57223 => -23437,
    57224 => -23435,
    57225 => -23433,
    57226 => -23430,
    57227 => -23428,
    57228 => -23426,
    57229 => -23424,
    57230 => -23422,
    57231 => -23419,
    57232 => -23417,
    57233 => -23415,
    57234 => -23413,
    57235 => -23411,
    57236 => -23408,
    57237 => -23406,
    57238 => -23404,
    57239 => -23402,
    57240 => -23400,
    57241 => -23397,
    57242 => -23395,
    57243 => -23393,
    57244 => -23391,
    57245 => -23389,
    57246 => -23386,
    57247 => -23384,
    57248 => -23382,
    57249 => -23380,
    57250 => -23378,
    57251 => -23375,
    57252 => -23373,
    57253 => -23371,
    57254 => -23369,
    57255 => -23367,
    57256 => -23364,
    57257 => -23362,
    57258 => -23360,
    57259 => -23358,
    57260 => -23356,
    57261 => -23353,
    57262 => -23351,
    57263 => -23349,
    57264 => -23347,
    57265 => -23345,
    57266 => -23342,
    57267 => -23340,
    57268 => -23338,
    57269 => -23336,
    57270 => -23334,
    57271 => -23331,
    57272 => -23329,
    57273 => -23327,
    57274 => -23325,
    57275 => -23323,
    57276 => -23320,
    57277 => -23318,
    57278 => -23316,
    57279 => -23314,
    57280 => -23311,
    57281 => -23309,
    57282 => -23307,
    57283 => -23305,
    57284 => -23303,
    57285 => -23300,
    57286 => -23298,
    57287 => -23296,
    57288 => -23294,
    57289 => -23292,
    57290 => -23289,
    57291 => -23287,
    57292 => -23285,
    57293 => -23283,
    57294 => -23281,
    57295 => -23278,
    57296 => -23276,
    57297 => -23274,
    57298 => -23272,
    57299 => -23270,
    57300 => -23267,
    57301 => -23265,
    57302 => -23263,
    57303 => -23261,
    57304 => -23258,
    57305 => -23256,
    57306 => -23254,
    57307 => -23252,
    57308 => -23250,
    57309 => -23247,
    57310 => -23245,
    57311 => -23243,
    57312 => -23241,
    57313 => -23239,
    57314 => -23236,
    57315 => -23234,
    57316 => -23232,
    57317 => -23230,
    57318 => -23227,
    57319 => -23225,
    57320 => -23223,
    57321 => -23221,
    57322 => -23219,
    57323 => -23216,
    57324 => -23214,
    57325 => -23212,
    57326 => -23210,
    57327 => -23208,
    57328 => -23205,
    57329 => -23203,
    57330 => -23201,
    57331 => -23199,
    57332 => -23196,
    57333 => -23194,
    57334 => -23192,
    57335 => -23190,
    57336 => -23188,
    57337 => -23185,
    57338 => -23183,
    57339 => -23181,
    57340 => -23179,
    57341 => -23176,
    57342 => -23174,
    57343 => -23172,
    57344 => -23170,
    57345 => -23168,
    57346 => -23165,
    57347 => -23163,
    57348 => -23161,
    57349 => -23159,
    57350 => -23156,
    57351 => -23154,
    57352 => -23152,
    57353 => -23150,
    57354 => -23148,
    57355 => -23145,
    57356 => -23143,
    57357 => -23141,
    57358 => -23139,
    57359 => -23136,
    57360 => -23134,
    57361 => -23132,
    57362 => -23130,
    57363 => -23128,
    57364 => -23125,
    57365 => -23123,
    57366 => -23121,
    57367 => -23119,
    57368 => -23116,
    57369 => -23114,
    57370 => -23112,
    57371 => -23110,
    57372 => -23107,
    57373 => -23105,
    57374 => -23103,
    57375 => -23101,
    57376 => -23099,
    57377 => -23096,
    57378 => -23094,
    57379 => -23092,
    57380 => -23090,
    57381 => -23087,
    57382 => -23085,
    57383 => -23083,
    57384 => -23081,
    57385 => -23079,
    57386 => -23076,
    57387 => -23074,
    57388 => -23072,
    57389 => -23070,
    57390 => -23067,
    57391 => -23065,
    57392 => -23063,
    57393 => -23061,
    57394 => -23058,
    57395 => -23056,
    57396 => -23054,
    57397 => -23052,
    57398 => -23050,
    57399 => -23047,
    57400 => -23045,
    57401 => -23043,
    57402 => -23041,
    57403 => -23038,
    57404 => -23036,
    57405 => -23034,
    57406 => -23032,
    57407 => -23029,
    57408 => -23027,
    57409 => -23025,
    57410 => -23023,
    57411 => -23020,
    57412 => -23018,
    57413 => -23016,
    57414 => -23014,
    57415 => -23012,
    57416 => -23009,
    57417 => -23007,
    57418 => -23005,
    57419 => -23003,
    57420 => -23000,
    57421 => -22998,
    57422 => -22996,
    57423 => -22994,
    57424 => -22991,
    57425 => -22989,
    57426 => -22987,
    57427 => -22985,
    57428 => -22982,
    57429 => -22980,
    57430 => -22978,
    57431 => -22976,
    57432 => -22973,
    57433 => -22971,
    57434 => -22969,
    57435 => -22967,
    57436 => -22965,
    57437 => -22962,
    57438 => -22960,
    57439 => -22958,
    57440 => -22956,
    57441 => -22953,
    57442 => -22951,
    57443 => -22949,
    57444 => -22947,
    57445 => -22944,
    57446 => -22942,
    57447 => -22940,
    57448 => -22938,
    57449 => -22935,
    57450 => -22933,
    57451 => -22931,
    57452 => -22929,
    57453 => -22926,
    57454 => -22924,
    57455 => -22922,
    57456 => -22920,
    57457 => -22917,
    57458 => -22915,
    57459 => -22913,
    57460 => -22911,
    57461 => -22908,
    57462 => -22906,
    57463 => -22904,
    57464 => -22902,
    57465 => -22899,
    57466 => -22897,
    57467 => -22895,
    57468 => -22893,
    57469 => -22890,
    57470 => -22888,
    57471 => -22886,
    57472 => -22884,
    57473 => -22881,
    57474 => -22879,
    57475 => -22877,
    57476 => -22875,
    57477 => -22872,
    57478 => -22870,
    57479 => -22868,
    57480 => -22866,
    57481 => -22863,
    57482 => -22861,
    57483 => -22859,
    57484 => -22857,
    57485 => -22854,
    57486 => -22852,
    57487 => -22850,
    57488 => -22848,
    57489 => -22845,
    57490 => -22843,
    57491 => -22841,
    57492 => -22839,
    57493 => -22836,
    57494 => -22834,
    57495 => -22832,
    57496 => -22830,
    57497 => -22827,
    57498 => -22825,
    57499 => -22823,
    57500 => -22821,
    57501 => -22818,
    57502 => -22816,
    57503 => -22814,
    57504 => -22812,
    57505 => -22809,
    57506 => -22807,
    57507 => -22805,
    57508 => -22803,
    57509 => -22800,
    57510 => -22798,
    57511 => -22796,
    57512 => -22794,
    57513 => -22791,
    57514 => -22789,
    57515 => -22787,
    57516 => -22785,
    57517 => -22782,
    57518 => -22780,
    57519 => -22778,
    57520 => -22776,
    57521 => -22773,
    57522 => -22771,
    57523 => -22769,
    57524 => -22766,
    57525 => -22764,
    57526 => -22762,
    57527 => -22760,
    57528 => -22757,
    57529 => -22755,
    57530 => -22753,
    57531 => -22751,
    57532 => -22748,
    57533 => -22746,
    57534 => -22744,
    57535 => -22742,
    57536 => -22739,
    57537 => -22737,
    57538 => -22735,
    57539 => -22733,
    57540 => -22730,
    57541 => -22728,
    57542 => -22726,
    57543 => -22724,
    57544 => -22721,
    57545 => -22719,
    57546 => -22717,
    57547 => -22714,
    57548 => -22712,
    57549 => -22710,
    57550 => -22708,
    57551 => -22705,
    57552 => -22703,
    57553 => -22701,
    57554 => -22699,
    57555 => -22696,
    57556 => -22694,
    57557 => -22692,
    57558 => -22690,
    57559 => -22687,
    57560 => -22685,
    57561 => -22683,
    57562 => -22680,
    57563 => -22678,
    57564 => -22676,
    57565 => -22674,
    57566 => -22671,
    57567 => -22669,
    57568 => -22667,
    57569 => -22665,
    57570 => -22662,
    57571 => -22660,
    57572 => -22658,
    57573 => -22656,
    57574 => -22653,
    57575 => -22651,
    57576 => -22649,
    57577 => -22646,
    57578 => -22644,
    57579 => -22642,
    57580 => -22640,
    57581 => -22637,
    57582 => -22635,
    57583 => -22633,
    57584 => -22631,
    57585 => -22628,
    57586 => -22626,
    57587 => -22624,
    57588 => -22621,
    57589 => -22619,
    57590 => -22617,
    57591 => -22615,
    57592 => -22612,
    57593 => -22610,
    57594 => -22608,
    57595 => -22606,
    57596 => -22603,
    57597 => -22601,
    57598 => -22599,
    57599 => -22596,
    57600 => -22594,
    57601 => -22592,
    57602 => -22590,
    57603 => -22587,
    57604 => -22585,
    57605 => -22583,
    57606 => -22581,
    57607 => -22578,
    57608 => -22576,
    57609 => -22574,
    57610 => -22571,
    57611 => -22569,
    57612 => -22567,
    57613 => -22565,
    57614 => -22562,
    57615 => -22560,
    57616 => -22558,
    57617 => -22555,
    57618 => -22553,
    57619 => -22551,
    57620 => -22549,
    57621 => -22546,
    57622 => -22544,
    57623 => -22542,
    57624 => -22540,
    57625 => -22537,
    57626 => -22535,
    57627 => -22533,
    57628 => -22530,
    57629 => -22528,
    57630 => -22526,
    57631 => -22524,
    57632 => -22521,
    57633 => -22519,
    57634 => -22517,
    57635 => -22514,
    57636 => -22512,
    57637 => -22510,
    57638 => -22508,
    57639 => -22505,
    57640 => -22503,
    57641 => -22501,
    57642 => -22498,
    57643 => -22496,
    57644 => -22494,
    57645 => -22492,
    57646 => -22489,
    57647 => -22487,
    57648 => -22485,
    57649 => -22482,
    57650 => -22480,
    57651 => -22478,
    57652 => -22476,
    57653 => -22473,
    57654 => -22471,
    57655 => -22469,
    57656 => -22466,
    57657 => -22464,
    57658 => -22462,
    57659 => -22460,
    57660 => -22457,
    57661 => -22455,
    57662 => -22453,
    57663 => -22450,
    57664 => -22448,
    57665 => -22446,
    57666 => -22444,
    57667 => -22441,
    57668 => -22439,
    57669 => -22437,
    57670 => -22434,
    57671 => -22432,
    57672 => -22430,
    57673 => -22428,
    57674 => -22425,
    57675 => -22423,
    57676 => -22421,
    57677 => -22418,
    57678 => -22416,
    57679 => -22414,
    57680 => -22411,
    57681 => -22409,
    57682 => -22407,
    57683 => -22405,
    57684 => -22402,
    57685 => -22400,
    57686 => -22398,
    57687 => -22395,
    57688 => -22393,
    57689 => -22391,
    57690 => -22389,
    57691 => -22386,
    57692 => -22384,
    57693 => -22382,
    57694 => -22379,
    57695 => -22377,
    57696 => -22375,
    57697 => -22373,
    57698 => -22370,
    57699 => -22368,
    57700 => -22366,
    57701 => -22363,
    57702 => -22361,
    57703 => -22359,
    57704 => -22356,
    57705 => -22354,
    57706 => -22352,
    57707 => -22350,
    57708 => -22347,
    57709 => -22345,
    57710 => -22343,
    57711 => -22340,
    57712 => -22338,
    57713 => -22336,
    57714 => -22333,
    57715 => -22331,
    57716 => -22329,
    57717 => -22327,
    57718 => -22324,
    57719 => -22322,
    57720 => -22320,
    57721 => -22317,
    57722 => -22315,
    57723 => -22313,
    57724 => -22310,
    57725 => -22308,
    57726 => -22306,
    57727 => -22304,
    57728 => -22301,
    57729 => -22299,
    57730 => -22297,
    57731 => -22294,
    57732 => -22292,
    57733 => -22290,
    57734 => -22287,
    57735 => -22285,
    57736 => -22283,
    57737 => -22281,
    57738 => -22278,
    57739 => -22276,
    57740 => -22274,
    57741 => -22271,
    57742 => -22269,
    57743 => -22267,
    57744 => -22264,
    57745 => -22262,
    57746 => -22260,
    57747 => -22257,
    57748 => -22255,
    57749 => -22253,
    57750 => -22251,
    57751 => -22248,
    57752 => -22246,
    57753 => -22244,
    57754 => -22241,
    57755 => -22239,
    57756 => -22237,
    57757 => -22234,
    57758 => -22232,
    57759 => -22230,
    57760 => -22227,
    57761 => -22225,
    57762 => -22223,
    57763 => -22221,
    57764 => -22218,
    57765 => -22216,
    57766 => -22214,
    57767 => -22211,
    57768 => -22209,
    57769 => -22207,
    57770 => -22204,
    57771 => -22202,
    57772 => -22200,
    57773 => -22197,
    57774 => -22195,
    57775 => -22193,
    57776 => -22191,
    57777 => -22188,
    57778 => -22186,
    57779 => -22184,
    57780 => -22181,
    57781 => -22179,
    57782 => -22177,
    57783 => -22174,
    57784 => -22172,
    57785 => -22170,
    57786 => -22167,
    57787 => -22165,
    57788 => -22163,
    57789 => -22160,
    57790 => -22158,
    57791 => -22156,
    57792 => -22154,
    57793 => -22151,
    57794 => -22149,
    57795 => -22147,
    57796 => -22144,
    57797 => -22142,
    57798 => -22140,
    57799 => -22137,
    57800 => -22135,
    57801 => -22133,
    57802 => -22130,
    57803 => -22128,
    57804 => -22126,
    57805 => -22123,
    57806 => -22121,
    57807 => -22119,
    57808 => -22116,
    57809 => -22114,
    57810 => -22112,
    57811 => -22110,
    57812 => -22107,
    57813 => -22105,
    57814 => -22103,
    57815 => -22100,
    57816 => -22098,
    57817 => -22096,
    57818 => -22093,
    57819 => -22091,
    57820 => -22089,
    57821 => -22086,
    57822 => -22084,
    57823 => -22082,
    57824 => -22079,
    57825 => -22077,
    57826 => -22075,
    57827 => -22072,
    57828 => -22070,
    57829 => -22068,
    57830 => -22065,
    57831 => -22063,
    57832 => -22061,
    57833 => -22058,
    57834 => -22056,
    57835 => -22054,
    57836 => -22051,
    57837 => -22049,
    57838 => -22047,
    57839 => -22045,
    57840 => -22042,
    57841 => -22040,
    57842 => -22038,
    57843 => -22035,
    57844 => -22033,
    57845 => -22031,
    57846 => -22028,
    57847 => -22026,
    57848 => -22024,
    57849 => -22021,
    57850 => -22019,
    57851 => -22017,
    57852 => -22014,
    57853 => -22012,
    57854 => -22010,
    57855 => -22007,
    57856 => -22005,
    57857 => -22003,
    57858 => -22000,
    57859 => -21998,
    57860 => -21996,
    57861 => -21993,
    57862 => -21991,
    57863 => -21989,
    57864 => -21986,
    57865 => -21984,
    57866 => -21982,
    57867 => -21979,
    57868 => -21977,
    57869 => -21975,
    57870 => -21972,
    57871 => -21970,
    57872 => -21968,
    57873 => -21965,
    57874 => -21963,
    57875 => -21961,
    57876 => -21958,
    57877 => -21956,
    57878 => -21954,
    57879 => -21951,
    57880 => -21949,
    57881 => -21947,
    57882 => -21944,
    57883 => -21942,
    57884 => -21940,
    57885 => -21937,
    57886 => -21935,
    57887 => -21933,
    57888 => -21930,
    57889 => -21928,
    57890 => -21926,
    57891 => -21923,
    57892 => -21921,
    57893 => -21919,
    57894 => -21916,
    57895 => -21914,
    57896 => -21912,
    57897 => -21909,
    57898 => -21907,
    57899 => -21905,
    57900 => -21902,
    57901 => -21900,
    57902 => -21898,
    57903 => -21895,
    57904 => -21893,
    57905 => -21891,
    57906 => -21888,
    57907 => -21886,
    57908 => -21884,
    57909 => -21881,
    57910 => -21879,
    57911 => -21877,
    57912 => -21874,
    57913 => -21872,
    57914 => -21870,
    57915 => -21867,
    57916 => -21865,
    57917 => -21863,
    57918 => -21860,
    57919 => -21858,
    57920 => -21856,
    57921 => -21853,
    57922 => -21851,
    57923 => -21849,
    57924 => -21846,
    57925 => -21844,
    57926 => -21842,
    57927 => -21839,
    57928 => -21837,
    57929 => -21835,
    57930 => -21832,
    57931 => -21830,
    57932 => -21827,
    57933 => -21825,
    57934 => -21823,
    57935 => -21820,
    57936 => -21818,
    57937 => -21816,
    57938 => -21813,
    57939 => -21811,
    57940 => -21809,
    57941 => -21806,
    57942 => -21804,
    57943 => -21802,
    57944 => -21799,
    57945 => -21797,
    57946 => -21795,
    57947 => -21792,
    57948 => -21790,
    57949 => -21788,
    57950 => -21785,
    57951 => -21783,
    57952 => -21781,
    57953 => -21778,
    57954 => -21776,
    57955 => -21774,
    57956 => -21771,
    57957 => -21769,
    57958 => -21766,
    57959 => -21764,
    57960 => -21762,
    57961 => -21759,
    57962 => -21757,
    57963 => -21755,
    57964 => -21752,
    57965 => -21750,
    57966 => -21748,
    57967 => -21745,
    57968 => -21743,
    57969 => -21741,
    57970 => -21738,
    57971 => -21736,
    57972 => -21734,
    57973 => -21731,
    57974 => -21729,
    57975 => -21727,
    57976 => -21724,
    57977 => -21722,
    57978 => -21719,
    57979 => -21717,
    57980 => -21715,
    57981 => -21712,
    57982 => -21710,
    57983 => -21708,
    57984 => -21705,
    57985 => -21703,
    57986 => -21701,
    57987 => -21698,
    57988 => -21696,
    57989 => -21694,
    57990 => -21691,
    57991 => -21689,
    57992 => -21687,
    57993 => -21684,
    57994 => -21682,
    57995 => -21679,
    57996 => -21677,
    57997 => -21675,
    57998 => -21672,
    57999 => -21670,
    58000 => -21668,
    58001 => -21665,
    58002 => -21663,
    58003 => -21661,
    58004 => -21658,
    58005 => -21656,
    58006 => -21654,
    58007 => -21651,
    58008 => -21649,
    58009 => -21646,
    58010 => -21644,
    58011 => -21642,
    58012 => -21639,
    58013 => -21637,
    58014 => -21635,
    58015 => -21632,
    58016 => -21630,
    58017 => -21628,
    58018 => -21625,
    58019 => -21623,
    58020 => -21621,
    58021 => -21618,
    58022 => -21616,
    58023 => -21613,
    58024 => -21611,
    58025 => -21609,
    58026 => -21606,
    58027 => -21604,
    58028 => -21602,
    58029 => -21599,
    58030 => -21597,
    58031 => -21595,
    58032 => -21592,
    58033 => -21590,
    58034 => -21587,
    58035 => -21585,
    58036 => -21583,
    58037 => -21580,
    58038 => -21578,
    58039 => -21576,
    58040 => -21573,
    58041 => -21571,
    58042 => -21569,
    58043 => -21566,
    58044 => -21564,
    58045 => -21561,
    58046 => -21559,
    58047 => -21557,
    58048 => -21554,
    58049 => -21552,
    58050 => -21550,
    58051 => -21547,
    58052 => -21545,
    58053 => -21543,
    58054 => -21540,
    58055 => -21538,
    58056 => -21535,
    58057 => -21533,
    58058 => -21531,
    58059 => -21528,
    58060 => -21526,
    58061 => -21524,
    58062 => -21521,
    58063 => -21519,
    58064 => -21516,
    58065 => -21514,
    58066 => -21512,
    58067 => -21509,
    58068 => -21507,
    58069 => -21505,
    58070 => -21502,
    58071 => -21500,
    58072 => -21498,
    58073 => -21495,
    58074 => -21493,
    58075 => -21490,
    58076 => -21488,
    58077 => -21486,
    58078 => -21483,
    58079 => -21481,
    58080 => -21479,
    58081 => -21476,
    58082 => -21474,
    58083 => -21471,
    58084 => -21469,
    58085 => -21467,
    58086 => -21464,
    58087 => -21462,
    58088 => -21460,
    58089 => -21457,
    58090 => -21455,
    58091 => -21452,
    58092 => -21450,
    58093 => -21448,
    58094 => -21445,
    58095 => -21443,
    58096 => -21441,
    58097 => -21438,
    58098 => -21436,
    58099 => -21433,
    58100 => -21431,
    58101 => -21429,
    58102 => -21426,
    58103 => -21424,
    58104 => -21422,
    58105 => -21419,
    58106 => -21417,
    58107 => -21414,
    58108 => -21412,
    58109 => -21410,
    58110 => -21407,
    58111 => -21405,
    58112 => -21403,
    58113 => -21400,
    58114 => -21398,
    58115 => -21395,
    58116 => -21393,
    58117 => -21391,
    58118 => -21388,
    58119 => -21386,
    58120 => -21383,
    58121 => -21381,
    58122 => -21379,
    58123 => -21376,
    58124 => -21374,
    58125 => -21372,
    58126 => -21369,
    58127 => -21367,
    58128 => -21364,
    58129 => -21362,
    58130 => -21360,
    58131 => -21357,
    58132 => -21355,
    58133 => -21353,
    58134 => -21350,
    58135 => -21348,
    58136 => -21345,
    58137 => -21343,
    58138 => -21341,
    58139 => -21338,
    58140 => -21336,
    58141 => -21333,
    58142 => -21331,
    58143 => -21329,
    58144 => -21326,
    58145 => -21324,
    58146 => -21322,
    58147 => -21319,
    58148 => -21317,
    58149 => -21314,
    58150 => -21312,
    58151 => -21310,
    58152 => -21307,
    58153 => -21305,
    58154 => -21302,
    58155 => -21300,
    58156 => -21298,
    58157 => -21295,
    58158 => -21293,
    58159 => -21290,
    58160 => -21288,
    58161 => -21286,
    58162 => -21283,
    58163 => -21281,
    58164 => -21279,
    58165 => -21276,
    58166 => -21274,
    58167 => -21271,
    58168 => -21269,
    58169 => -21267,
    58170 => -21264,
    58171 => -21262,
    58172 => -21259,
    58173 => -21257,
    58174 => -21255,
    58175 => -21252,
    58176 => -21250,
    58177 => -21247,
    58178 => -21245,
    58179 => -21243,
    58180 => -21240,
    58181 => -21238,
    58182 => -21236,
    58183 => -21233,
    58184 => -21231,
    58185 => -21228,
    58186 => -21226,
    58187 => -21224,
    58188 => -21221,
    58189 => -21219,
    58190 => -21216,
    58191 => -21214,
    58192 => -21212,
    58193 => -21209,
    58194 => -21207,
    58195 => -21204,
    58196 => -21202,
    58197 => -21200,
    58198 => -21197,
    58199 => -21195,
    58200 => -21192,
    58201 => -21190,
    58202 => -21188,
    58203 => -21185,
    58204 => -21183,
    58205 => -21180,
    58206 => -21178,
    58207 => -21176,
    58208 => -21173,
    58209 => -21171,
    58210 => -21168,
    58211 => -21166,
    58212 => -21164,
    58213 => -21161,
    58214 => -21159,
    58215 => -21156,
    58216 => -21154,
    58217 => -21152,
    58218 => -21149,
    58219 => -21147,
    58220 => -21144,
    58221 => -21142,
    58222 => -21140,
    58223 => -21137,
    58224 => -21135,
    58225 => -21132,
    58226 => -21130,
    58227 => -21128,
    58228 => -21125,
    58229 => -21123,
    58230 => -21120,
    58231 => -21118,
    58232 => -21116,
    58233 => -21113,
    58234 => -21111,
    58235 => -21108,
    58236 => -21106,
    58237 => -21104,
    58238 => -21101,
    58239 => -21099,
    58240 => -21096,
    58241 => -21094,
    58242 => -21092,
    58243 => -21089,
    58244 => -21087,
    58245 => -21084,
    58246 => -21082,
    58247 => -21080,
    58248 => -21077,
    58249 => -21075,
    58250 => -21072,
    58251 => -21070,
    58252 => -21068,
    58253 => -21065,
    58254 => -21063,
    58255 => -21060,
    58256 => -21058,
    58257 => -21056,
    58258 => -21053,
    58259 => -21051,
    58260 => -21048,
    58261 => -21046,
    58262 => -21043,
    58263 => -21041,
    58264 => -21039,
    58265 => -21036,
    58266 => -21034,
    58267 => -21031,
    58268 => -21029,
    58269 => -21027,
    58270 => -21024,
    58271 => -21022,
    58272 => -21019,
    58273 => -21017,
    58274 => -21015,
    58275 => -21012,
    58276 => -21010,
    58277 => -21007,
    58278 => -21005,
    58279 => -21003,
    58280 => -21000,
    58281 => -20998,
    58282 => -20995,
    58283 => -20993,
    58284 => -20990,
    58285 => -20988,
    58286 => -20986,
    58287 => -20983,
    58288 => -20981,
    58289 => -20978,
    58290 => -20976,
    58291 => -20974,
    58292 => -20971,
    58293 => -20969,
    58294 => -20966,
    58295 => -20964,
    58296 => -20962,
    58297 => -20959,
    58298 => -20957,
    58299 => -20954,
    58300 => -20952,
    58301 => -20949,
    58302 => -20947,
    58303 => -20945,
    58304 => -20942,
    58305 => -20940,
    58306 => -20937,
    58307 => -20935,
    58308 => -20933,
    58309 => -20930,
    58310 => -20928,
    58311 => -20925,
    58312 => -20923,
    58313 => -20920,
    58314 => -20918,
    58315 => -20916,
    58316 => -20913,
    58317 => -20911,
    58318 => -20908,
    58319 => -20906,
    58320 => -20904,
    58321 => -20901,
    58322 => -20899,
    58323 => -20896,
    58324 => -20894,
    58325 => -20891,
    58326 => -20889,
    58327 => -20887,
    58328 => -20884,
    58329 => -20882,
    58330 => -20879,
    58331 => -20877,
    58332 => -20874,
    58333 => -20872,
    58334 => -20870,
    58335 => -20867,
    58336 => -20865,
    58337 => -20862,
    58338 => -20860,
    58339 => -20858,
    58340 => -20855,
    58341 => -20853,
    58342 => -20850,
    58343 => -20848,
    58344 => -20845,
    58345 => -20843,
    58346 => -20841,
    58347 => -20838,
    58348 => -20836,
    58349 => -20833,
    58350 => -20831,
    58351 => -20828,
    58352 => -20826,
    58353 => -20824,
    58354 => -20821,
    58355 => -20819,
    58356 => -20816,
    58357 => -20814,
    58358 => -20811,
    58359 => -20809,
    58360 => -20807,
    58361 => -20804,
    58362 => -20802,
    58363 => -20799,
    58364 => -20797,
    58365 => -20794,
    58366 => -20792,
    58367 => -20790,
    58368 => -20787,
    58369 => -20785,
    58370 => -20782,
    58371 => -20780,
    58372 => -20777,
    58373 => -20775,
    58374 => -20773,
    58375 => -20770,
    58376 => -20768,
    58377 => -20765,
    58378 => -20763,
    58379 => -20760,
    58380 => -20758,
    58381 => -20756,
    58382 => -20753,
    58383 => -20751,
    58384 => -20748,
    58385 => -20746,
    58386 => -20743,
    58387 => -20741,
    58388 => -20739,
    58389 => -20736,
    58390 => -20734,
    58391 => -20731,
    58392 => -20729,
    58393 => -20726,
    58394 => -20724,
    58395 => -20722,
    58396 => -20719,
    58397 => -20717,
    58398 => -20714,
    58399 => -20712,
    58400 => -20709,
    58401 => -20707,
    58402 => -20704,
    58403 => -20702,
    58404 => -20700,
    58405 => -20697,
    58406 => -20695,
    58407 => -20692,
    58408 => -20690,
    58409 => -20687,
    58410 => -20685,
    58411 => -20683,
    58412 => -20680,
    58413 => -20678,
    58414 => -20675,
    58415 => -20673,
    58416 => -20670,
    58417 => -20668,
    58418 => -20666,
    58419 => -20663,
    58420 => -20661,
    58421 => -20658,
    58422 => -20656,
    58423 => -20653,
    58424 => -20651,
    58425 => -20648,
    58426 => -20646,
    58427 => -20644,
    58428 => -20641,
    58429 => -20639,
    58430 => -20636,
    58431 => -20634,
    58432 => -20631,
    58433 => -20629,
    58434 => -20626,
    58435 => -20624,
    58436 => -20622,
    58437 => -20619,
    58438 => -20617,
    58439 => -20614,
    58440 => -20612,
    58441 => -20609,
    58442 => -20607,
    58443 => -20604,
    58444 => -20602,
    58445 => -20600,
    58446 => -20597,
    58447 => -20595,
    58448 => -20592,
    58449 => -20590,
    58450 => -20587,
    58451 => -20585,
    58452 => -20583,
    58453 => -20580,
    58454 => -20578,
    58455 => -20575,
    58456 => -20573,
    58457 => -20570,
    58458 => -20568,
    58459 => -20565,
    58460 => -20563,
    58461 => -20560,
    58462 => -20558,
    58463 => -20556,
    58464 => -20553,
    58465 => -20551,
    58466 => -20548,
    58467 => -20546,
    58468 => -20543,
    58469 => -20541,
    58470 => -20538,
    58471 => -20536,
    58472 => -20534,
    58473 => -20531,
    58474 => -20529,
    58475 => -20526,
    58476 => -20524,
    58477 => -20521,
    58478 => -20519,
    58479 => -20516,
    58480 => -20514,
    58481 => -20512,
    58482 => -20509,
    58483 => -20507,
    58484 => -20504,
    58485 => -20502,
    58486 => -20499,
    58487 => -20497,
    58488 => -20494,
    58489 => -20492,
    58490 => -20489,
    58491 => -20487,
    58492 => -20485,
    58493 => -20482,
    58494 => -20480,
    58495 => -20477,
    58496 => -20475,
    58497 => -20472,
    58498 => -20470,
    58499 => -20467,
    58500 => -20465,
    58501 => -20463,
    58502 => -20460,
    58503 => -20458,
    58504 => -20455,
    58505 => -20453,
    58506 => -20450,
    58507 => -20448,
    58508 => -20445,
    58509 => -20443,
    58510 => -20440,
    58511 => -20438,
    58512 => -20436,
    58513 => -20433,
    58514 => -20431,
    58515 => -20428,
    58516 => -20426,
    58517 => -20423,
    58518 => -20421,
    58519 => -20418,
    58520 => -20416,
    58521 => -20413,
    58522 => -20411,
    58523 => -20408,
    58524 => -20406,
    58525 => -20404,
    58526 => -20401,
    58527 => -20399,
    58528 => -20396,
    58529 => -20394,
    58530 => -20391,
    58531 => -20389,
    58532 => -20386,
    58533 => -20384,
    58534 => -20381,
    58535 => -20379,
    58536 => -20377,
    58537 => -20374,
    58538 => -20372,
    58539 => -20369,
    58540 => -20367,
    58541 => -20364,
    58542 => -20362,
    58543 => -20359,
    58544 => -20357,
    58545 => -20354,
    58546 => -20352,
    58547 => -20349,
    58548 => -20347,
    58549 => -20345,
    58550 => -20342,
    58551 => -20340,
    58552 => -20337,
    58553 => -20335,
    58554 => -20332,
    58555 => -20330,
    58556 => -20327,
    58557 => -20325,
    58558 => -20322,
    58559 => -20320,
    58560 => -20317,
    58561 => -20315,
    58562 => -20312,
    58563 => -20310,
    58564 => -20308,
    58565 => -20305,
    58566 => -20303,
    58567 => -20300,
    58568 => -20298,
    58569 => -20295,
    58570 => -20293,
    58571 => -20290,
    58572 => -20288,
    58573 => -20285,
    58574 => -20283,
    58575 => -20280,
    58576 => -20278,
    58577 => -20275,
    58578 => -20273,
    58579 => -20271,
    58580 => -20268,
    58581 => -20266,
    58582 => -20263,
    58583 => -20261,
    58584 => -20258,
    58585 => -20256,
    58586 => -20253,
    58587 => -20251,
    58588 => -20248,
    58589 => -20246,
    58590 => -20243,
    58591 => -20241,
    58592 => -20238,
    58593 => -20236,
    58594 => -20234,
    58595 => -20231,
    58596 => -20229,
    58597 => -20226,
    58598 => -20224,
    58599 => -20221,
    58600 => -20219,
    58601 => -20216,
    58602 => -20214,
    58603 => -20211,
    58604 => -20209,
    58605 => -20206,
    58606 => -20204,
    58607 => -20201,
    58608 => -20199,
    58609 => -20196,
    58610 => -20194,
    58611 => -20191,
    58612 => -20189,
    58613 => -20187,
    58614 => -20184,
    58615 => -20182,
    58616 => -20179,
    58617 => -20177,
    58618 => -20174,
    58619 => -20172,
    58620 => -20169,
    58621 => -20167,
    58622 => -20164,
    58623 => -20162,
    58624 => -20159,
    58625 => -20157,
    58626 => -20154,
    58627 => -20152,
    58628 => -20149,
    58629 => -20147,
    58630 => -20144,
    58631 => -20142,
    58632 => -20139,
    58633 => -20137,
    58634 => -20135,
    58635 => -20132,
    58636 => -20130,
    58637 => -20127,
    58638 => -20125,
    58639 => -20122,
    58640 => -20120,
    58641 => -20117,
    58642 => -20115,
    58643 => -20112,
    58644 => -20110,
    58645 => -20107,
    58646 => -20105,
    58647 => -20102,
    58648 => -20100,
    58649 => -20097,
    58650 => -20095,
    58651 => -20092,
    58652 => -20090,
    58653 => -20087,
    58654 => -20085,
    58655 => -20082,
    58656 => -20080,
    58657 => -20077,
    58658 => -20075,
    58659 => -20072,
    58660 => -20070,
    58661 => -20068,
    58662 => -20065,
    58663 => -20063,
    58664 => -20060,
    58665 => -20058,
    58666 => -20055,
    58667 => -20053,
    58668 => -20050,
    58669 => -20048,
    58670 => -20045,
    58671 => -20043,
    58672 => -20040,
    58673 => -20038,
    58674 => -20035,
    58675 => -20033,
    58676 => -20030,
    58677 => -20028,
    58678 => -20025,
    58679 => -20023,
    58680 => -20020,
    58681 => -20018,
    58682 => -20015,
    58683 => -20013,
    58684 => -20010,
    58685 => -20008,
    58686 => -20005,
    58687 => -20003,
    58688 => -20000,
    58689 => -19998,
    58690 => -19995,
    58691 => -19993,
    58692 => -19990,
    58693 => -19988,
    58694 => -19985,
    58695 => -19983,
    58696 => -19981,
    58697 => -19978,
    58698 => -19976,
    58699 => -19973,
    58700 => -19971,
    58701 => -19968,
    58702 => -19966,
    58703 => -19963,
    58704 => -19961,
    58705 => -19958,
    58706 => -19956,
    58707 => -19953,
    58708 => -19951,
    58709 => -19948,
    58710 => -19946,
    58711 => -19943,
    58712 => -19941,
    58713 => -19938,
    58714 => -19936,
    58715 => -19933,
    58716 => -19931,
    58717 => -19928,
    58718 => -19926,
    58719 => -19923,
    58720 => -19921,
    58721 => -19918,
    58722 => -19916,
    58723 => -19913,
    58724 => -19911,
    58725 => -19908,
    58726 => -19906,
    58727 => -19903,
    58728 => -19901,
    58729 => -19898,
    58730 => -19896,
    58731 => -19893,
    58732 => -19891,
    58733 => -19888,
    58734 => -19886,
    58735 => -19883,
    58736 => -19881,
    58737 => -19878,
    58738 => -19876,
    58739 => -19873,
    58740 => -19871,
    58741 => -19868,
    58742 => -19866,
    58743 => -19863,
    58744 => -19861,
    58745 => -19858,
    58746 => -19856,
    58747 => -19853,
    58748 => -19851,
    58749 => -19848,
    58750 => -19846,
    58751 => -19843,
    58752 => -19841,
    58753 => -19838,
    58754 => -19836,
    58755 => -19833,
    58756 => -19831,
    58757 => -19828,
    58758 => -19826,
    58759 => -19823,
    58760 => -19821,
    58761 => -19818,
    58762 => -19816,
    58763 => -19813,
    58764 => -19811,
    58765 => -19808,
    58766 => -19806,
    58767 => -19803,
    58768 => -19801,
    58769 => -19798,
    58770 => -19796,
    58771 => -19793,
    58772 => -19791,
    58773 => -19788,
    58774 => -19786,
    58775 => -19783,
    58776 => -19781,
    58777 => -19778,
    58778 => -19776,
    58779 => -19773,
    58780 => -19771,
    58781 => -19768,
    58782 => -19766,
    58783 => -19763,
    58784 => -19761,
    58785 => -19758,
    58786 => -19756,
    58787 => -19753,
    58788 => -19751,
    58789 => -19748,
    58790 => -19746,
    58791 => -19743,
    58792 => -19741,
    58793 => -19738,
    58794 => -19736,
    58795 => -19733,
    58796 => -19731,
    58797 => -19728,
    58798 => -19726,
    58799 => -19723,
    58800 => -19721,
    58801 => -19718,
    58802 => -19716,
    58803 => -19713,
    58804 => -19711,
    58805 => -19708,
    58806 => -19706,
    58807 => -19703,
    58808 => -19700,
    58809 => -19698,
    58810 => -19695,
    58811 => -19693,
    58812 => -19690,
    58813 => -19688,
    58814 => -19685,
    58815 => -19683,
    58816 => -19680,
    58817 => -19678,
    58818 => -19675,
    58819 => -19673,
    58820 => -19670,
    58821 => -19668,
    58822 => -19665,
    58823 => -19663,
    58824 => -19660,
    58825 => -19658,
    58826 => -19655,
    58827 => -19653,
    58828 => -19650,
    58829 => -19648,
    58830 => -19645,
    58831 => -19643,
    58832 => -19640,
    58833 => -19638,
    58834 => -19635,
    58835 => -19633,
    58836 => -19630,
    58837 => -19628,
    58838 => -19625,
    58839 => -19623,
    58840 => -19620,
    58841 => -19618,
    58842 => -19615,
    58843 => -19613,
    58844 => -19610,
    58845 => -19607,
    58846 => -19605,
    58847 => -19602,
    58848 => -19600,
    58849 => -19597,
    58850 => -19595,
    58851 => -19592,
    58852 => -19590,
    58853 => -19587,
    58854 => -19585,
    58855 => -19582,
    58856 => -19580,
    58857 => -19577,
    58858 => -19575,
    58859 => -19572,
    58860 => -19570,
    58861 => -19567,
    58862 => -19565,
    58863 => -19562,
    58864 => -19560,
    58865 => -19557,
    58866 => -19555,
    58867 => -19552,
    58868 => -19550,
    58869 => -19547,
    58870 => -19545,
    58871 => -19542,
    58872 => -19539,
    58873 => -19537,
    58874 => -19534,
    58875 => -19532,
    58876 => -19529,
    58877 => -19527,
    58878 => -19524,
    58879 => -19522,
    58880 => -19519,
    58881 => -19517,
    58882 => -19514,
    58883 => -19512,
    58884 => -19509,
    58885 => -19507,
    58886 => -19504,
    58887 => -19502,
    58888 => -19499,
    58889 => -19497,
    58890 => -19494,
    58891 => -19492,
    58892 => -19489,
    58893 => -19486,
    58894 => -19484,
    58895 => -19481,
    58896 => -19479,
    58897 => -19476,
    58898 => -19474,
    58899 => -19471,
    58900 => -19469,
    58901 => -19466,
    58902 => -19464,
    58903 => -19461,
    58904 => -19459,
    58905 => -19456,
    58906 => -19454,
    58907 => -19451,
    58908 => -19449,
    58909 => -19446,
    58910 => -19444,
    58911 => -19441,
    58912 => -19438,
    58913 => -19436,
    58914 => -19433,
    58915 => -19431,
    58916 => -19428,
    58917 => -19426,
    58918 => -19423,
    58919 => -19421,
    58920 => -19418,
    58921 => -19416,
    58922 => -19413,
    58923 => -19411,
    58924 => -19408,
    58925 => -19406,
    58926 => -19403,
    58927 => -19400,
    58928 => -19398,
    58929 => -19395,
    58930 => -19393,
    58931 => -19390,
    58932 => -19388,
    58933 => -19385,
    58934 => -19383,
    58935 => -19380,
    58936 => -19378,
    58937 => -19375,
    58938 => -19373,
    58939 => -19370,
    58940 => -19368,
    58941 => -19365,
    58942 => -19362,
    58943 => -19360,
    58944 => -19357,
    58945 => -19355,
    58946 => -19352,
    58947 => -19350,
    58948 => -19347,
    58949 => -19345,
    58950 => -19342,
    58951 => -19340,
    58952 => -19337,
    58953 => -19335,
    58954 => -19332,
    58955 => -19330,
    58956 => -19327,
    58957 => -19324,
    58958 => -19322,
    58959 => -19319,
    58960 => -19317,
    58961 => -19314,
    58962 => -19312,
    58963 => -19309,
    58964 => -19307,
    58965 => -19304,
    58966 => -19302,
    58967 => -19299,
    58968 => -19297,
    58969 => -19294,
    58970 => -19291,
    58971 => -19289,
    58972 => -19286,
    58973 => -19284,
    58974 => -19281,
    58975 => -19279,
    58976 => -19276,
    58977 => -19274,
    58978 => -19271,
    58979 => -19269,
    58980 => -19266,
    58981 => -19264,
    58982 => -19261,
    58983 => -19258,
    58984 => -19256,
    58985 => -19253,
    58986 => -19251,
    58987 => -19248,
    58988 => -19246,
    58989 => -19243,
    58990 => -19241,
    58991 => -19238,
    58992 => -19236,
    58993 => -19233,
    58994 => -19230,
    58995 => -19228,
    58996 => -19225,
    58997 => -19223,
    58998 => -19220,
    58999 => -19218,
    59000 => -19215,
    59001 => -19213,
    59002 => -19210,
    59003 => -19208,
    59004 => -19205,
    59005 => -19202,
    59006 => -19200,
    59007 => -19197,
    59008 => -19195,
    59009 => -19192,
    59010 => -19190,
    59011 => -19187,
    59012 => -19185,
    59013 => -19182,
    59014 => -19180,
    59015 => -19177,
    59016 => -19174,
    59017 => -19172,
    59018 => -19169,
    59019 => -19167,
    59020 => -19164,
    59021 => -19162,
    59022 => -19159,
    59023 => -19157,
    59024 => -19154,
    59025 => -19152,
    59026 => -19149,
    59027 => -19146,
    59028 => -19144,
    59029 => -19141,
    59030 => -19139,
    59031 => -19136,
    59032 => -19134,
    59033 => -19131,
    59034 => -19129,
    59035 => -19126,
    59036 => -19123,
    59037 => -19121,
    59038 => -19118,
    59039 => -19116,
    59040 => -19113,
    59041 => -19111,
    59042 => -19108,
    59043 => -19106,
    59044 => -19103,
    59045 => -19101,
    59046 => -19098,
    59047 => -19095,
    59048 => -19093,
    59049 => -19090,
    59050 => -19088,
    59051 => -19085,
    59052 => -19083,
    59053 => -19080,
    59054 => -19078,
    59055 => -19075,
    59056 => -19072,
    59057 => -19070,
    59058 => -19067,
    59059 => -19065,
    59060 => -19062,
    59061 => -19060,
    59062 => -19057,
    59063 => -19055,
    59064 => -19052,
    59065 => -19049,
    59066 => -19047,
    59067 => -19044,
    59068 => -19042,
    59069 => -19039,
    59070 => -19037,
    59071 => -19034,
    59072 => -19032,
    59073 => -19029,
    59074 => -19026,
    59075 => -19024,
    59076 => -19021,
    59077 => -19019,
    59078 => -19016,
    59079 => -19014,
    59080 => -19011,
    59081 => -19009,
    59082 => -19006,
    59083 => -19003,
    59084 => -19001,
    59085 => -18998,
    59086 => -18996,
    59087 => -18993,
    59088 => -18991,
    59089 => -18988,
    59090 => -18985,
    59091 => -18983,
    59092 => -18980,
    59093 => -18978,
    59094 => -18975,
    59095 => -18973,
    59096 => -18970,
    59097 => -18968,
    59098 => -18965,
    59099 => -18962,
    59100 => -18960,
    59101 => -18957,
    59102 => -18955,
    59103 => -18952,
    59104 => -18950,
    59105 => -18947,
    59106 => -18944,
    59107 => -18942,
    59108 => -18939,
    59109 => -18937,
    59110 => -18934,
    59111 => -18932,
    59112 => -18929,
    59113 => -18927,
    59114 => -18924,
    59115 => -18921,
    59116 => -18919,
    59117 => -18916,
    59118 => -18914,
    59119 => -18911,
    59120 => -18909,
    59121 => -18906,
    59122 => -18903,
    59123 => -18901,
    59124 => -18898,
    59125 => -18896,
    59126 => -18893,
    59127 => -18891,
    59128 => -18888,
    59129 => -18885,
    59130 => -18883,
    59131 => -18880,
    59132 => -18878,
    59133 => -18875,
    59134 => -18873,
    59135 => -18870,
    59136 => -18868,
    59137 => -18865,
    59138 => -18862,
    59139 => -18860,
    59140 => -18857,
    59141 => -18855,
    59142 => -18852,
    59143 => -18850,
    59144 => -18847,
    59145 => -18844,
    59146 => -18842,
    59147 => -18839,
    59148 => -18837,
    59149 => -18834,
    59150 => -18832,
    59151 => -18829,
    59152 => -18826,
    59153 => -18824,
    59154 => -18821,
    59155 => -18819,
    59156 => -18816,
    59157 => -18814,
    59158 => -18811,
    59159 => -18808,
    59160 => -18806,
    59161 => -18803,
    59162 => -18801,
    59163 => -18798,
    59164 => -18796,
    59165 => -18793,
    59166 => -18790,
    59167 => -18788,
    59168 => -18785,
    59169 => -18783,
    59170 => -18780,
    59171 => -18778,
    59172 => -18775,
    59173 => -18772,
    59174 => -18770,
    59175 => -18767,
    59176 => -18765,
    59177 => -18762,
    59178 => -18759,
    59179 => -18757,
    59180 => -18754,
    59181 => -18752,
    59182 => -18749,
    59183 => -18747,
    59184 => -18744,
    59185 => -18741,
    59186 => -18739,
    59187 => -18736,
    59188 => -18734,
    59189 => -18731,
    59190 => -18729,
    59191 => -18726,
    59192 => -18723,
    59193 => -18721,
    59194 => -18718,
    59195 => -18716,
    59196 => -18713,
    59197 => -18711,
    59198 => -18708,
    59199 => -18705,
    59200 => -18703,
    59201 => -18700,
    59202 => -18698,
    59203 => -18695,
    59204 => -18692,
    59205 => -18690,
    59206 => -18687,
    59207 => -18685,
    59208 => -18682,
    59209 => -18680,
    59210 => -18677,
    59211 => -18674,
    59212 => -18672,
    59213 => -18669,
    59214 => -18667,
    59215 => -18664,
    59216 => -18661,
    59217 => -18659,
    59218 => -18656,
    59219 => -18654,
    59220 => -18651,
    59221 => -18649,
    59222 => -18646,
    59223 => -18643,
    59224 => -18641,
    59225 => -18638,
    59226 => -18636,
    59227 => -18633,
    59228 => -18630,
    59229 => -18628,
    59230 => -18625,
    59231 => -18623,
    59232 => -18620,
    59233 => -18618,
    59234 => -18615,
    59235 => -18612,
    59236 => -18610,
    59237 => -18607,
    59238 => -18605,
    59239 => -18602,
    59240 => -18599,
    59241 => -18597,
    59242 => -18594,
    59243 => -18592,
    59244 => -18589,
    59245 => -18587,
    59246 => -18584,
    59247 => -18581,
    59248 => -18579,
    59249 => -18576,
    59250 => -18574,
    59251 => -18571,
    59252 => -18568,
    59253 => -18566,
    59254 => -18563,
    59255 => -18561,
    59256 => -18558,
    59257 => -18555,
    59258 => -18553,
    59259 => -18550,
    59260 => -18548,
    59261 => -18545,
    59262 => -18543,
    59263 => -18540,
    59264 => -18537,
    59265 => -18535,
    59266 => -18532,
    59267 => -18530,
    59268 => -18527,
    59269 => -18524,
    59270 => -18522,
    59271 => -18519,
    59272 => -18517,
    59273 => -18514,
    59274 => -18511,
    59275 => -18509,
    59276 => -18506,
    59277 => -18504,
    59278 => -18501,
    59279 => -18498,
    59280 => -18496,
    59281 => -18493,
    59282 => -18491,
    59283 => -18488,
    59284 => -18485,
    59285 => -18483,
    59286 => -18480,
    59287 => -18478,
    59288 => -18475,
    59289 => -18473,
    59290 => -18470,
    59291 => -18467,
    59292 => -18465,
    59293 => -18462,
    59294 => -18460,
    59295 => -18457,
    59296 => -18454,
    59297 => -18452,
    59298 => -18449,
    59299 => -18447,
    59300 => -18444,
    59301 => -18441,
    59302 => -18439,
    59303 => -18436,
    59304 => -18434,
    59305 => -18431,
    59306 => -18428,
    59307 => -18426,
    59308 => -18423,
    59309 => -18421,
    59310 => -18418,
    59311 => -18415,
    59312 => -18413,
    59313 => -18410,
    59314 => -18408,
    59315 => -18405,
    59316 => -18402,
    59317 => -18400,
    59318 => -18397,
    59319 => -18395,
    59320 => -18392,
    59321 => -18389,
    59322 => -18387,
    59323 => -18384,
    59324 => -18382,
    59325 => -18379,
    59326 => -18376,
    59327 => -18374,
    59328 => -18371,
    59329 => -18369,
    59330 => -18366,
    59331 => -18363,
    59332 => -18361,
    59333 => -18358,
    59334 => -18356,
    59335 => -18353,
    59336 => -18350,
    59337 => -18348,
    59338 => -18345,
    59339 => -18343,
    59340 => -18340,
    59341 => -18337,
    59342 => -18335,
    59343 => -18332,
    59344 => -18330,
    59345 => -18327,
    59346 => -18324,
    59347 => -18322,
    59348 => -18319,
    59349 => -18317,
    59350 => -18314,
    59351 => -18311,
    59352 => -18309,
    59353 => -18306,
    59354 => -18304,
    59355 => -18301,
    59356 => -18298,
    59357 => -18296,
    59358 => -18293,
    59359 => -18290,
    59360 => -18288,
    59361 => -18285,
    59362 => -18283,
    59363 => -18280,
    59364 => -18277,
    59365 => -18275,
    59366 => -18272,
    59367 => -18270,
    59368 => -18267,
    59369 => -18264,
    59370 => -18262,
    59371 => -18259,
    59372 => -18257,
    59373 => -18254,
    59374 => -18251,
    59375 => -18249,
    59376 => -18246,
    59377 => -18244,
    59378 => -18241,
    59379 => -18238,
    59380 => -18236,
    59381 => -18233,
    59382 => -18230,
    59383 => -18228,
    59384 => -18225,
    59385 => -18223,
    59386 => -18220,
    59387 => -18217,
    59388 => -18215,
    59389 => -18212,
    59390 => -18210,
    59391 => -18207,
    59392 => -18204,
    59393 => -18202,
    59394 => -18199,
    59395 => -18197,
    59396 => -18194,
    59397 => -18191,
    59398 => -18189,
    59399 => -18186,
    59400 => -18183,
    59401 => -18181,
    59402 => -18178,
    59403 => -18176,
    59404 => -18173,
    59405 => -18170,
    59406 => -18168,
    59407 => -18165,
    59408 => -18163,
    59409 => -18160,
    59410 => -18157,
    59411 => -18155,
    59412 => -18152,
    59413 => -18149,
    59414 => -18147,
    59415 => -18144,
    59416 => -18142,
    59417 => -18139,
    59418 => -18136,
    59419 => -18134,
    59420 => -18131,
    59421 => -18129,
    59422 => -18126,
    59423 => -18123,
    59424 => -18121,
    59425 => -18118,
    59426 => -18115,
    59427 => -18113,
    59428 => -18110,
    59429 => -18108,
    59430 => -18105,
    59431 => -18102,
    59432 => -18100,
    59433 => -18097,
    59434 => -18095,
    59435 => -18092,
    59436 => -18089,
    59437 => -18087,
    59438 => -18084,
    59439 => -18081,
    59440 => -18079,
    59441 => -18076,
    59442 => -18074,
    59443 => -18071,
    59444 => -18068,
    59445 => -18066,
    59446 => -18063,
    59447 => -18060,
    59448 => -18058,
    59449 => -18055,
    59450 => -18053,
    59451 => -18050,
    59452 => -18047,
    59453 => -18045,
    59454 => -18042,
    59455 => -18039,
    59456 => -18037,
    59457 => -18034,
    59458 => -18032,
    59459 => -18029,
    59460 => -18026,
    59461 => -18024,
    59462 => -18021,
    59463 => -18018,
    59464 => -18016,
    59465 => -18013,
    59466 => -18011,
    59467 => -18008,
    59468 => -18005,
    59469 => -18003,
    59470 => -18000,
    59471 => -17997,
    59472 => -17995,
    59473 => -17992,
    59474 => -17990,
    59475 => -17987,
    59476 => -17984,
    59477 => -17982,
    59478 => -17979,
    59479 => -17976,
    59480 => -17974,
    59481 => -17971,
    59482 => -17969,
    59483 => -17966,
    59484 => -17963,
    59485 => -17961,
    59486 => -17958,
    59487 => -17955,
    59488 => -17953,
    59489 => -17950,
    59490 => -17948,
    59491 => -17945,
    59492 => -17942,
    59493 => -17940,
    59494 => -17937,
    59495 => -17934,
    59496 => -17932,
    59497 => -17929,
    59498 => -17927,
    59499 => -17924,
    59500 => -17921,
    59501 => -17919,
    59502 => -17916,
    59503 => -17913,
    59504 => -17911,
    59505 => -17908,
    59506 => -17906,
    59507 => -17903,
    59508 => -17900,
    59509 => -17898,
    59510 => -17895,
    59511 => -17892,
    59512 => -17890,
    59513 => -17887,
    59514 => -17884,
    59515 => -17882,
    59516 => -17879,
    59517 => -17877,
    59518 => -17874,
    59519 => -17871,
    59520 => -17869,
    59521 => -17866,
    59522 => -17863,
    59523 => -17861,
    59524 => -17858,
    59525 => -17855,
    59526 => -17853,
    59527 => -17850,
    59528 => -17848,
    59529 => -17845,
    59530 => -17842,
    59531 => -17840,
    59532 => -17837,
    59533 => -17834,
    59534 => -17832,
    59535 => -17829,
    59536 => -17827,
    59537 => -17824,
    59538 => -17821,
    59539 => -17819,
    59540 => -17816,
    59541 => -17813,
    59542 => -17811,
    59543 => -17808,
    59544 => -17805,
    59545 => -17803,
    59546 => -17800,
    59547 => -17798,
    59548 => -17795,
    59549 => -17792,
    59550 => -17790,
    59551 => -17787,
    59552 => -17784,
    59553 => -17782,
    59554 => -17779,
    59555 => -17776,
    59556 => -17774,
    59557 => -17771,
    59558 => -17768,
    59559 => -17766,
    59560 => -17763,
    59561 => -17761,
    59562 => -17758,
    59563 => -17755,
    59564 => -17753,
    59565 => -17750,
    59566 => -17747,
    59567 => -17745,
    59568 => -17742,
    59569 => -17739,
    59570 => -17737,
    59571 => -17734,
    59572 => -17732,
    59573 => -17729,
    59574 => -17726,
    59575 => -17724,
    59576 => -17721,
    59577 => -17718,
    59578 => -17716,
    59579 => -17713,
    59580 => -17710,
    59581 => -17708,
    59582 => -17705,
    59583 => -17702,
    59584 => -17700,
    59585 => -17697,
    59586 => -17695,
    59587 => -17692,
    59588 => -17689,
    59589 => -17687,
    59590 => -17684,
    59591 => -17681,
    59592 => -17679,
    59593 => -17676,
    59594 => -17673,
    59595 => -17671,
    59596 => -17668,
    59597 => -17665,
    59598 => -17663,
    59599 => -17660,
    59600 => -17657,
    59601 => -17655,
    59602 => -17652,
    59603 => -17650,
    59604 => -17647,
    59605 => -17644,
    59606 => -17642,
    59607 => -17639,
    59608 => -17636,
    59609 => -17634,
    59610 => -17631,
    59611 => -17628,
    59612 => -17626,
    59613 => -17623,
    59614 => -17620,
    59615 => -17618,
    59616 => -17615,
    59617 => -17612,
    59618 => -17610,
    59619 => -17607,
    59620 => -17605,
    59621 => -17602,
    59622 => -17599,
    59623 => -17597,
    59624 => -17594,
    59625 => -17591,
    59626 => -17589,
    59627 => -17586,
    59628 => -17583,
    59629 => -17581,
    59630 => -17578,
    59631 => -17575,
    59632 => -17573,
    59633 => -17570,
    59634 => -17567,
    59635 => -17565,
    59636 => -17562,
    59637 => -17559,
    59638 => -17557,
    59639 => -17554,
    59640 => -17551,
    59641 => -17549,
    59642 => -17546,
    59643 => -17544,
    59644 => -17541,
    59645 => -17538,
    59646 => -17536,
    59647 => -17533,
    59648 => -17530,
    59649 => -17528,
    59650 => -17525,
    59651 => -17522,
    59652 => -17520,
    59653 => -17517,
    59654 => -17514,
    59655 => -17512,
    59656 => -17509,
    59657 => -17506,
    59658 => -17504,
    59659 => -17501,
    59660 => -17498,
    59661 => -17496,
    59662 => -17493,
    59663 => -17490,
    59664 => -17488,
    59665 => -17485,
    59666 => -17482,
    59667 => -17480,
    59668 => -17477,
    59669 => -17474,
    59670 => -17472,
    59671 => -17469,
    59672 => -17467,
    59673 => -17464,
    59674 => -17461,
    59675 => -17459,
    59676 => -17456,
    59677 => -17453,
    59678 => -17451,
    59679 => -17448,
    59680 => -17445,
    59681 => -17443,
    59682 => -17440,
    59683 => -17437,
    59684 => -17435,
    59685 => -17432,
    59686 => -17429,
    59687 => -17427,
    59688 => -17424,
    59689 => -17421,
    59690 => -17419,
    59691 => -17416,
    59692 => -17413,
    59693 => -17411,
    59694 => -17408,
    59695 => -17405,
    59696 => -17403,
    59697 => -17400,
    59698 => -17397,
    59699 => -17395,
    59700 => -17392,
    59701 => -17389,
    59702 => -17387,
    59703 => -17384,
    59704 => -17381,
    59705 => -17379,
    59706 => -17376,
    59707 => -17373,
    59708 => -17371,
    59709 => -17368,
    59710 => -17365,
    59711 => -17363,
    59712 => -17360,
    59713 => -17357,
    59714 => -17355,
    59715 => -17352,
    59716 => -17349,
    59717 => -17347,
    59718 => -17344,
    59719 => -17341,
    59720 => -17339,
    59721 => -17336,
    59722 => -17333,
    59723 => -17331,
    59724 => -17328,
    59725 => -17325,
    59726 => -17323,
    59727 => -17320,
    59728 => -17317,
    59729 => -17315,
    59730 => -17312,
    59731 => -17309,
    59732 => -17307,
    59733 => -17304,
    59734 => -17301,
    59735 => -17299,
    59736 => -17296,
    59737 => -17293,
    59738 => -17291,
    59739 => -17288,
    59740 => -17285,
    59741 => -17283,
    59742 => -17280,
    59743 => -17277,
    59744 => -17275,
    59745 => -17272,
    59746 => -17269,
    59747 => -17267,
    59748 => -17264,
    59749 => -17261,
    59750 => -17259,
    59751 => -17256,
    59752 => -17253,
    59753 => -17251,
    59754 => -17248,
    59755 => -17245,
    59756 => -17243,
    59757 => -17240,
    59758 => -17237,
    59759 => -17235,
    59760 => -17232,
    59761 => -17229,
    59762 => -17227,
    59763 => -17224,
    59764 => -17221,
    59765 => -17219,
    59766 => -17216,
    59767 => -17213,
    59768 => -17211,
    59769 => -17208,
    59770 => -17205,
    59771 => -17203,
    59772 => -17200,
    59773 => -17197,
    59774 => -17195,
    59775 => -17192,
    59776 => -17189,
    59777 => -17187,
    59778 => -17184,
    59779 => -17181,
    59780 => -17179,
    59781 => -17176,
    59782 => -17173,
    59783 => -17171,
    59784 => -17168,
    59785 => -17165,
    59786 => -17162,
    59787 => -17160,
    59788 => -17157,
    59789 => -17154,
    59790 => -17152,
    59791 => -17149,
    59792 => -17146,
    59793 => -17144,
    59794 => -17141,
    59795 => -17138,
    59796 => -17136,
    59797 => -17133,
    59798 => -17130,
    59799 => -17128,
    59800 => -17125,
    59801 => -17122,
    59802 => -17120,
    59803 => -17117,
    59804 => -17114,
    59805 => -17112,
    59806 => -17109,
    59807 => -17106,
    59808 => -17104,
    59809 => -17101,
    59810 => -17098,
    59811 => -17096,
    59812 => -17093,
    59813 => -17090,
    59814 => -17087,
    59815 => -17085,
    59816 => -17082,
    59817 => -17079,
    59818 => -17077,
    59819 => -17074,
    59820 => -17071,
    59821 => -17069,
    59822 => -17066,
    59823 => -17063,
    59824 => -17061,
    59825 => -17058,
    59826 => -17055,
    59827 => -17053,
    59828 => -17050,
    59829 => -17047,
    59830 => -17045,
    59831 => -17042,
    59832 => -17039,
    59833 => -17037,
    59834 => -17034,
    59835 => -17031,
    59836 => -17028,
    59837 => -17026,
    59838 => -17023,
    59839 => -17020,
    59840 => -17018,
    59841 => -17015,
    59842 => -17012,
    59843 => -17010,
    59844 => -17007,
    59845 => -17004,
    59846 => -17002,
    59847 => -16999,
    59848 => -16996,
    59849 => -16994,
    59850 => -16991,
    59851 => -16988,
    59852 => -16986,
    59853 => -16983,
    59854 => -16980,
    59855 => -16977,
    59856 => -16975,
    59857 => -16972,
    59858 => -16969,
    59859 => -16967,
    59860 => -16964,
    59861 => -16961,
    59862 => -16959,
    59863 => -16956,
    59864 => -16953,
    59865 => -16951,
    59866 => -16948,
    59867 => -16945,
    59868 => -16943,
    59869 => -16940,
    59870 => -16937,
    59871 => -16934,
    59872 => -16932,
    59873 => -16929,
    59874 => -16926,
    59875 => -16924,
    59876 => -16921,
    59877 => -16918,
    59878 => -16916,
    59879 => -16913,
    59880 => -16910,
    59881 => -16908,
    59882 => -16905,
    59883 => -16902,
    59884 => -16899,
    59885 => -16897,
    59886 => -16894,
    59887 => -16891,
    59888 => -16889,
    59889 => -16886,
    59890 => -16883,
    59891 => -16881,
    59892 => -16878,
    59893 => -16875,
    59894 => -16873,
    59895 => -16870,
    59896 => -16867,
    59897 => -16864,
    59898 => -16862,
    59899 => -16859,
    59900 => -16856,
    59901 => -16854,
    59902 => -16851,
    59903 => -16848,
    59904 => -16846,
    59905 => -16843,
    59906 => -16840,
    59907 => -16838,
    59908 => -16835,
    59909 => -16832,
    59910 => -16829,
    59911 => -16827,
    59912 => -16824,
    59913 => -16821,
    59914 => -16819,
    59915 => -16816,
    59916 => -16813,
    59917 => -16811,
    59918 => -16808,
    59919 => -16805,
    59920 => -16802,
    59921 => -16800,
    59922 => -16797,
    59923 => -16794,
    59924 => -16792,
    59925 => -16789,
    59926 => -16786,
    59927 => -16784,
    59928 => -16781,
    59929 => -16778,
    59930 => -16775,
    59931 => -16773,
    59932 => -16770,
    59933 => -16767,
    59934 => -16765,
    59935 => -16762,
    59936 => -16759,
    59937 => -16757,
    59938 => -16754,
    59939 => -16751,
    59940 => -16749,
    59941 => -16746,
    59942 => -16743,
    59943 => -16740,
    59944 => -16738,
    59945 => -16735,
    59946 => -16732,
    59947 => -16730,
    59948 => -16727,
    59949 => -16724,
    59950 => -16721,
    59951 => -16719,
    59952 => -16716,
    59953 => -16713,
    59954 => -16711,
    59955 => -16708,
    59956 => -16705,
    59957 => -16703,
    59958 => -16700,
    59959 => -16697,
    59960 => -16694,
    59961 => -16692,
    59962 => -16689,
    59963 => -16686,
    59964 => -16684,
    59965 => -16681,
    59966 => -16678,
    59967 => -16676,
    59968 => -16673,
    59969 => -16670,
    59970 => -16667,
    59971 => -16665,
    59972 => -16662,
    59973 => -16659,
    59974 => -16657,
    59975 => -16654,
    59976 => -16651,
    59977 => -16648,
    59978 => -16646,
    59979 => -16643,
    59980 => -16640,
    59981 => -16638,
    59982 => -16635,
    59983 => -16632,
    59984 => -16630,
    59985 => -16627,
    59986 => -16624,
    59987 => -16621,
    59988 => -16619,
    59989 => -16616,
    59990 => -16613,
    59991 => -16611,
    59992 => -16608,
    59993 => -16605,
    59994 => -16602,
    59995 => -16600,
    59996 => -16597,
    59997 => -16594,
    59998 => -16592,
    59999 => -16589,
    60000 => -16586,
    60001 => -16584,
    60002 => -16581,
    60003 => -16578,
    60004 => -16575,
    60005 => -16573,
    60006 => -16570,
    60007 => -16567,
    60008 => -16565,
    60009 => -16562,
    60010 => -16559,
    60011 => -16556,
    60012 => -16554,
    60013 => -16551,
    60014 => -16548,
    60015 => -16546,
    60016 => -16543,
    60017 => -16540,
    60018 => -16537,
    60019 => -16535,
    60020 => -16532,
    60021 => -16529,
    60022 => -16527,
    60023 => -16524,
    60024 => -16521,
    60025 => -16518,
    60026 => -16516,
    60027 => -16513,
    60028 => -16510,
    60029 => -16508,
    60030 => -16505,
    60031 => -16502,
    60032 => -16499,
    60033 => -16497,
    60034 => -16494,
    60035 => -16491,
    60036 => -16489,
    60037 => -16486,
    60038 => -16483,
    60039 => -16480,
    60040 => -16478,
    60041 => -16475,
    60042 => -16472,
    60043 => -16470,
    60044 => -16467,
    60045 => -16464,
    60046 => -16461,
    60047 => -16459,
    60048 => -16456,
    60049 => -16453,
    60050 => -16451,
    60051 => -16448,
    60052 => -16445,
    60053 => -16442,
    60054 => -16440,
    60055 => -16437,
    60056 => -16434,
    60057 => -16432,
    60058 => -16429,
    60059 => -16426,
    60060 => -16423,
    60061 => -16421,
    60062 => -16418,
    60063 => -16415,
    60064 => -16413,
    60065 => -16410,
    60066 => -16407,
    60067 => -16404,
    60068 => -16402,
    60069 => -16399,
    60070 => -16396,
    60071 => -16393,
    60072 => -16391,
    60073 => -16388,
    60074 => -16385,
    60075 => -16383,
    60076 => -16380,
    60077 => -16377,
    60078 => -16374,
    60079 => -16372,
    60080 => -16369,
    60081 => -16366,
    60082 => -16364,
    60083 => -16361,
    60084 => -16358,
    60085 => -16355,
    60086 => -16353,
    60087 => -16350,
    60088 => -16347,
    60089 => -16344,
    60090 => -16342,
    60091 => -16339,
    60092 => -16336,
    60093 => -16334,
    60094 => -16331,
    60095 => -16328,
    60096 => -16325,
    60097 => -16323,
    60098 => -16320,
    60099 => -16317,
    60100 => -16315,
    60101 => -16312,
    60102 => -16309,
    60103 => -16306,
    60104 => -16304,
    60105 => -16301,
    60106 => -16298,
    60107 => -16295,
    60108 => -16293,
    60109 => -16290,
    60110 => -16287,
    60111 => -16285,
    60112 => -16282,
    60113 => -16279,
    60114 => -16276,
    60115 => -16274,
    60116 => -16271,
    60117 => -16268,
    60118 => -16265,
    60119 => -16263,
    60120 => -16260,
    60121 => -16257,
    60122 => -16255,
    60123 => -16252,
    60124 => -16249,
    60125 => -16246,
    60126 => -16244,
    60127 => -16241,
    60128 => -16238,
    60129 => -16235,
    60130 => -16233,
    60131 => -16230,
    60132 => -16227,
    60133 => -16225,
    60134 => -16222,
    60135 => -16219,
    60136 => -16216,
    60137 => -16214,
    60138 => -16211,
    60139 => -16208,
    60140 => -16205,
    60141 => -16203,
    60142 => -16200,
    60143 => -16197,
    60144 => -16195,
    60145 => -16192,
    60146 => -16189,
    60147 => -16186,
    60148 => -16184,
    60149 => -16181,
    60150 => -16178,
    60151 => -16175,
    60152 => -16173,
    60153 => -16170,
    60154 => -16167,
    60155 => -16164,
    60156 => -16162,
    60157 => -16159,
    60158 => -16156,
    60159 => -16154,
    60160 => -16151,
    60161 => -16148,
    60162 => -16145,
    60163 => -16143,
    60164 => -16140,
    60165 => -16137,
    60166 => -16134,
    60167 => -16132,
    60168 => -16129,
    60169 => -16126,
    60170 => -16123,
    60171 => -16121,
    60172 => -16118,
    60173 => -16115,
    60174 => -16113,
    60175 => -16110,
    60176 => -16107,
    60177 => -16104,
    60178 => -16102,
    60179 => -16099,
    60180 => -16096,
    60181 => -16093,
    60182 => -16091,
    60183 => -16088,
    60184 => -16085,
    60185 => -16082,
    60186 => -16080,
    60187 => -16077,
    60188 => -16074,
    60189 => -16071,
    60190 => -16069,
    60191 => -16066,
    60192 => -16063,
    60193 => -16061,
    60194 => -16058,
    60195 => -16055,
    60196 => -16052,
    60197 => -16050,
    60198 => -16047,
    60199 => -16044,
    60200 => -16041,
    60201 => -16039,
    60202 => -16036,
    60203 => -16033,
    60204 => -16030,
    60205 => -16028,
    60206 => -16025,
    60207 => -16022,
    60208 => -16019,
    60209 => -16017,
    60210 => -16014,
    60211 => -16011,
    60212 => -16008,
    60213 => -16006,
    60214 => -16003,
    60215 => -16000,
    60216 => -15997,
    60217 => -15995,
    60218 => -15992,
    60219 => -15989,
    60220 => -15987,
    60221 => -15984,
    60222 => -15981,
    60223 => -15978,
    60224 => -15976,
    60225 => -15973,
    60226 => -15970,
    60227 => -15967,
    60228 => -15965,
    60229 => -15962,
    60230 => -15959,
    60231 => -15956,
    60232 => -15954,
    60233 => -15951,
    60234 => -15948,
    60235 => -15945,
    60236 => -15943,
    60237 => -15940,
    60238 => -15937,
    60239 => -15934,
    60240 => -15932,
    60241 => -15929,
    60242 => -15926,
    60243 => -15923,
    60244 => -15921,
    60245 => -15918,
    60246 => -15915,
    60247 => -15912,
    60248 => -15910,
    60249 => -15907,
    60250 => -15904,
    60251 => -15901,
    60252 => -15899,
    60253 => -15896,
    60254 => -15893,
    60255 => -15890,
    60256 => -15888,
    60257 => -15885,
    60258 => -15882,
    60259 => -15879,
    60260 => -15877,
    60261 => -15874,
    60262 => -15871,
    60263 => -15868,
    60264 => -15866,
    60265 => -15863,
    60266 => -15860,
    60267 => -15857,
    60268 => -15855,
    60269 => -15852,
    60270 => -15849,
    60271 => -15846,
    60272 => -15844,
    60273 => -15841,
    60274 => -15838,
    60275 => -15835,
    60276 => -15833,
    60277 => -15830,
    60278 => -15827,
    60279 => -15824,
    60280 => -15822,
    60281 => -15819,
    60282 => -15816,
    60283 => -15813,
    60284 => -15811,
    60285 => -15808,
    60286 => -15805,
    60287 => -15802,
    60288 => -15800,
    60289 => -15797,
    60290 => -15794,
    60291 => -15791,
    60292 => -15789,
    60293 => -15786,
    60294 => -15783,
    60295 => -15780,
    60296 => -15778,
    60297 => -15775,
    60298 => -15772,
    60299 => -15769,
    60300 => -15767,
    60301 => -15764,
    60302 => -15761,
    60303 => -15758,
    60304 => -15756,
    60305 => -15753,
    60306 => -15750,
    60307 => -15747,
    60308 => -15745,
    60309 => -15742,
    60310 => -15739,
    60311 => -15736,
    60312 => -15734,
    60313 => -15731,
    60314 => -15728,
    60315 => -15725,
    60316 => -15723,
    60317 => -15720,
    60318 => -15717,
    60319 => -15714,
    60320 => -15712,
    60321 => -15709,
    60322 => -15706,
    60323 => -15703,
    60324 => -15701,
    60325 => -15698,
    60326 => -15695,
    60327 => -15692,
    60328 => -15690,
    60329 => -15687,
    60330 => -15684,
    60331 => -15681,
    60332 => -15678,
    60333 => -15676,
    60334 => -15673,
    60335 => -15670,
    60336 => -15667,
    60337 => -15665,
    60338 => -15662,
    60339 => -15659,
    60340 => -15656,
    60341 => -15654,
    60342 => -15651,
    60343 => -15648,
    60344 => -15645,
    60345 => -15643,
    60346 => -15640,
    60347 => -15637,
    60348 => -15634,
    60349 => -15632,
    60350 => -15629,
    60351 => -15626,
    60352 => -15623,
    60353 => -15621,
    60354 => -15618,
    60355 => -15615,
    60356 => -15612,
    60357 => -15609,
    60358 => -15607,
    60359 => -15604,
    60360 => -15601,
    60361 => -15598,
    60362 => -15596,
    60363 => -15593,
    60364 => -15590,
    60365 => -15587,
    60366 => -15585,
    60367 => -15582,
    60368 => -15579,
    60369 => -15576,
    60370 => -15574,
    60371 => -15571,
    60372 => -15568,
    60373 => -15565,
    60374 => -15562,
    60375 => -15560,
    60376 => -15557,
    60377 => -15554,
    60378 => -15551,
    60379 => -15549,
    60380 => -15546,
    60381 => -15543,
    60382 => -15540,
    60383 => -15538,
    60384 => -15535,
    60385 => -15532,
    60386 => -15529,
    60387 => -15527,
    60388 => -15524,
    60389 => -15521,
    60390 => -15518,
    60391 => -15515,
    60392 => -15513,
    60393 => -15510,
    60394 => -15507,
    60395 => -15504,
    60396 => -15502,
    60397 => -15499,
    60398 => -15496,
    60399 => -15493,
    60400 => -15491,
    60401 => -15488,
    60402 => -15485,
    60403 => -15482,
    60404 => -15479,
    60405 => -15477,
    60406 => -15474,
    60407 => -15471,
    60408 => -15468,
    60409 => -15466,
    60410 => -15463,
    60411 => -15460,
    60412 => -15457,
    60413 => -15455,
    60414 => -15452,
    60415 => -15449,
    60416 => -15446,
    60417 => -15443,
    60418 => -15441,
    60419 => -15438,
    60420 => -15435,
    60421 => -15432,
    60422 => -15430,
    60423 => -15427,
    60424 => -15424,
    60425 => -15421,
    60426 => -15419,
    60427 => -15416,
    60428 => -15413,
    60429 => -15410,
    60430 => -15407,
    60431 => -15405,
    60432 => -15402,
    60433 => -15399,
    60434 => -15396,
    60435 => -15394,
    60436 => -15391,
    60437 => -15388,
    60438 => -15385,
    60439 => -15382,
    60440 => -15380,
    60441 => -15377,
    60442 => -15374,
    60443 => -15371,
    60444 => -15369,
    60445 => -15366,
    60446 => -15363,
    60447 => -15360,
    60448 => -15358,
    60449 => -15355,
    60450 => -15352,
    60451 => -15349,
    60452 => -15346,
    60453 => -15344,
    60454 => -15341,
    60455 => -15338,
    60456 => -15335,
    60457 => -15333,
    60458 => -15330,
    60459 => -15327,
    60460 => -15324,
    60461 => -15321,
    60462 => -15319,
    60463 => -15316,
    60464 => -15313,
    60465 => -15310,
    60466 => -15308,
    60467 => -15305,
    60468 => -15302,
    60469 => -15299,
    60470 => -15296,
    60471 => -15294,
    60472 => -15291,
    60473 => -15288,
    60474 => -15285,
    60475 => -15283,
    60476 => -15280,
    60477 => -15277,
    60478 => -15274,
    60479 => -15271,
    60480 => -15269,
    60481 => -15266,
    60482 => -15263,
    60483 => -15260,
    60484 => -15258,
    60485 => -15255,
    60486 => -15252,
    60487 => -15249,
    60488 => -15246,
    60489 => -15244,
    60490 => -15241,
    60491 => -15238,
    60492 => -15235,
    60493 => -15233,
    60494 => -15230,
    60495 => -15227,
    60496 => -15224,
    60497 => -15221,
    60498 => -15219,
    60499 => -15216,
    60500 => -15213,
    60501 => -15210,
    60502 => -15207,
    60503 => -15205,
    60504 => -15202,
    60505 => -15199,
    60506 => -15196,
    60507 => -15194,
    60508 => -15191,
    60509 => -15188,
    60510 => -15185,
    60511 => -15182,
    60512 => -15180,
    60513 => -15177,
    60514 => -15174,
    60515 => -15171,
    60516 => -15168,
    60517 => -15166,
    60518 => -15163,
    60519 => -15160,
    60520 => -15157,
    60521 => -15155,
    60522 => -15152,
    60523 => -15149,
    60524 => -15146,
    60525 => -15143,
    60526 => -15141,
    60527 => -15138,
    60528 => -15135,
    60529 => -15132,
    60530 => -15129,
    60531 => -15127,
    60532 => -15124,
    60533 => -15121,
    60534 => -15118,
    60535 => -15116,
    60536 => -15113,
    60537 => -15110,
    60538 => -15107,
    60539 => -15104,
    60540 => -15102,
    60541 => -15099,
    60542 => -15096,
    60543 => -15093,
    60544 => -15090,
    60545 => -15088,
    60546 => -15085,
    60547 => -15082,
    60548 => -15079,
    60549 => -15077,
    60550 => -15074,
    60551 => -15071,
    60552 => -15068,
    60553 => -15065,
    60554 => -15063,
    60555 => -15060,
    60556 => -15057,
    60557 => -15054,
    60558 => -15051,
    60559 => -15049,
    60560 => -15046,
    60561 => -15043,
    60562 => -15040,
    60563 => -15037,
    60564 => -15035,
    60565 => -15032,
    60566 => -15029,
    60567 => -15026,
    60568 => -15024,
    60569 => -15021,
    60570 => -15018,
    60571 => -15015,
    60572 => -15012,
    60573 => -15010,
    60574 => -15007,
    60575 => -15004,
    60576 => -15001,
    60577 => -14998,
    60578 => -14996,
    60579 => -14993,
    60580 => -14990,
    60581 => -14987,
    60582 => -14984,
    60583 => -14982,
    60584 => -14979,
    60585 => -14976,
    60586 => -14973,
    60587 => -14970,
    60588 => -14968,
    60589 => -14965,
    60590 => -14962,
    60591 => -14959,
    60592 => -14956,
    60593 => -14954,
    60594 => -14951,
    60595 => -14948,
    60596 => -14945,
    60597 => -14942,
    60598 => -14940,
    60599 => -14937,
    60600 => -14934,
    60601 => -14931,
    60602 => -14929,
    60603 => -14926,
    60604 => -14923,
    60605 => -14920,
    60606 => -14917,
    60607 => -14915,
    60608 => -14912,
    60609 => -14909,
    60610 => -14906,
    60611 => -14903,
    60612 => -14901,
    60613 => -14898,
    60614 => -14895,
    60615 => -14892,
    60616 => -14889,
    60617 => -14887,
    60618 => -14884,
    60619 => -14881,
    60620 => -14878,
    60621 => -14875,
    60622 => -14873,
    60623 => -14870,
    60624 => -14867,
    60625 => -14864,
    60626 => -14861,
    60627 => -14859,
    60628 => -14856,
    60629 => -14853,
    60630 => -14850,
    60631 => -14847,
    60632 => -14845,
    60633 => -14842,
    60634 => -14839,
    60635 => -14836,
    60636 => -14833,
    60637 => -14831,
    60638 => -14828,
    60639 => -14825,
    60640 => -14822,
    60641 => -14819,
    60642 => -14817,
    60643 => -14814,
    60644 => -14811,
    60645 => -14808,
    60646 => -14805,
    60647 => -14803,
    60648 => -14800,
    60649 => -14797,
    60650 => -14794,
    60651 => -14791,
    60652 => -14789,
    60653 => -14786,
    60654 => -14783,
    60655 => -14780,
    60656 => -14777,
    60657 => -14774,
    60658 => -14772,
    60659 => -14769,
    60660 => -14766,
    60661 => -14763,
    60662 => -14760,
    60663 => -14758,
    60664 => -14755,
    60665 => -14752,
    60666 => -14749,
    60667 => -14746,
    60668 => -14744,
    60669 => -14741,
    60670 => -14738,
    60671 => -14735,
    60672 => -14732,
    60673 => -14730,
    60674 => -14727,
    60675 => -14724,
    60676 => -14721,
    60677 => -14718,
    60678 => -14716,
    60679 => -14713,
    60680 => -14710,
    60681 => -14707,
    60682 => -14704,
    60683 => -14702,
    60684 => -14699,
    60685 => -14696,
    60686 => -14693,
    60687 => -14690,
    60688 => -14688,
    60689 => -14685,
    60690 => -14682,
    60691 => -14679,
    60692 => -14676,
    60693 => -14673,
    60694 => -14671,
    60695 => -14668,
    60696 => -14665,
    60697 => -14662,
    60698 => -14659,
    60699 => -14657,
    60700 => -14654,
    60701 => -14651,
    60702 => -14648,
    60703 => -14645,
    60704 => -14643,
    60705 => -14640,
    60706 => -14637,
    60707 => -14634,
    60708 => -14631,
    60709 => -14628,
    60710 => -14626,
    60711 => -14623,
    60712 => -14620,
    60713 => -14617,
    60714 => -14614,
    60715 => -14612,
    60716 => -14609,
    60717 => -14606,
    60718 => -14603,
    60719 => -14600,
    60720 => -14598,
    60721 => -14595,
    60722 => -14592,
    60723 => -14589,
    60724 => -14586,
    60725 => -14584,
    60726 => -14581,
    60727 => -14578,
    60728 => -14575,
    60729 => -14572,
    60730 => -14569,
    60731 => -14567,
    60732 => -14564,
    60733 => -14561,
    60734 => -14558,
    60735 => -14555,
    60736 => -14553,
    60737 => -14550,
    60738 => -14547,
    60739 => -14544,
    60740 => -14541,
    60741 => -14538,
    60742 => -14536,
    60743 => -14533,
    60744 => -14530,
    60745 => -14527,
    60746 => -14524,
    60747 => -14522,
    60748 => -14519,
    60749 => -14516,
    60750 => -14513,
    60751 => -14510,
    60752 => -14507,
    60753 => -14505,
    60754 => -14502,
    60755 => -14499,
    60756 => -14496,
    60757 => -14493,
    60758 => -14491,
    60759 => -14488,
    60760 => -14485,
    60761 => -14482,
    60762 => -14479,
    60763 => -14477,
    60764 => -14474,
    60765 => -14471,
    60766 => -14468,
    60767 => -14465,
    60768 => -14462,
    60769 => -14460,
    60770 => -14457,
    60771 => -14454,
    60772 => -14451,
    60773 => -14448,
    60774 => -14445,
    60775 => -14443,
    60776 => -14440,
    60777 => -14437,
    60778 => -14434,
    60779 => -14431,
    60780 => -14429,
    60781 => -14426,
    60782 => -14423,
    60783 => -14420,
    60784 => -14417,
    60785 => -14414,
    60786 => -14412,
    60787 => -14409,
    60788 => -14406,
    60789 => -14403,
    60790 => -14400,
    60791 => -14398,
    60792 => -14395,
    60793 => -14392,
    60794 => -14389,
    60795 => -14386,
    60796 => -14383,
    60797 => -14381,
    60798 => -14378,
    60799 => -14375,
    60800 => -14372,
    60801 => -14369,
    60802 => -14366,
    60803 => -14364,
    60804 => -14361,
    60805 => -14358,
    60806 => -14355,
    60807 => -14352,
    60808 => -14350,
    60809 => -14347,
    60810 => -14344,
    60811 => -14341,
    60812 => -14338,
    60813 => -14335,
    60814 => -14333,
    60815 => -14330,
    60816 => -14327,
    60817 => -14324,
    60818 => -14321,
    60819 => -14318,
    60820 => -14316,
    60821 => -14313,
    60822 => -14310,
    60823 => -14307,
    60824 => -14304,
    60825 => -14302,
    60826 => -14299,
    60827 => -14296,
    60828 => -14293,
    60829 => -14290,
    60830 => -14287,
    60831 => -14285,
    60832 => -14282,
    60833 => -14279,
    60834 => -14276,
    60835 => -14273,
    60836 => -14270,
    60837 => -14268,
    60838 => -14265,
    60839 => -14262,
    60840 => -14259,
    60841 => -14256,
    60842 => -14253,
    60843 => -14251,
    60844 => -14248,
    60845 => -14245,
    60846 => -14242,
    60847 => -14239,
    60848 => -14236,
    60849 => -14234,
    60850 => -14231,
    60851 => -14228,
    60852 => -14225,
    60853 => -14222,
    60854 => -14219,
    60855 => -14217,
    60856 => -14214,
    60857 => -14211,
    60858 => -14208,
    60859 => -14205,
    60860 => -14203,
    60861 => -14200,
    60862 => -14197,
    60863 => -14194,
    60864 => -14191,
    60865 => -14188,
    60866 => -14186,
    60867 => -14183,
    60868 => -14180,
    60869 => -14177,
    60870 => -14174,
    60871 => -14171,
    60872 => -14169,
    60873 => -14166,
    60874 => -14163,
    60875 => -14160,
    60876 => -14157,
    60877 => -14154,
    60878 => -14152,
    60879 => -14149,
    60880 => -14146,
    60881 => -14143,
    60882 => -14140,
    60883 => -14137,
    60884 => -14135,
    60885 => -14132,
    60886 => -14129,
    60887 => -14126,
    60888 => -14123,
    60889 => -14120,
    60890 => -14118,
    60891 => -14115,
    60892 => -14112,
    60893 => -14109,
    60894 => -14106,
    60895 => -14103,
    60896 => -14101,
    60897 => -14098,
    60898 => -14095,
    60899 => -14092,
    60900 => -14089,
    60901 => -14086,
    60902 => -14083,
    60903 => -14081,
    60904 => -14078,
    60905 => -14075,
    60906 => -14072,
    60907 => -14069,
    60908 => -14066,
    60909 => -14064,
    60910 => -14061,
    60911 => -14058,
    60912 => -14055,
    60913 => -14052,
    60914 => -14049,
    60915 => -14047,
    60916 => -14044,
    60917 => -14041,
    60918 => -14038,
    60919 => -14035,
    60920 => -14032,
    60921 => -14030,
    60922 => -14027,
    60923 => -14024,
    60924 => -14021,
    60925 => -14018,
    60926 => -14015,
    60927 => -14013,
    60928 => -14010,
    60929 => -14007,
    60930 => -14004,
    60931 => -14001,
    60932 => -13998,
    60933 => -13995,
    60934 => -13993,
    60935 => -13990,
    60936 => -13987,
    60937 => -13984,
    60938 => -13981,
    60939 => -13978,
    60940 => -13976,
    60941 => -13973,
    60942 => -13970,
    60943 => -13967,
    60944 => -13964,
    60945 => -13961,
    60946 => -13959,
    60947 => -13956,
    60948 => -13953,
    60949 => -13950,
    60950 => -13947,
    60951 => -13944,
    60952 => -13942,
    60953 => -13939,
    60954 => -13936,
    60955 => -13933,
    60956 => -13930,
    60957 => -13927,
    60958 => -13924,
    60959 => -13922,
    60960 => -13919,
    60961 => -13916,
    60962 => -13913,
    60963 => -13910,
    60964 => -13907,
    60965 => -13905,
    60966 => -13902,
    60967 => -13899,
    60968 => -13896,
    60969 => -13893,
    60970 => -13890,
    60971 => -13887,
    60972 => -13885,
    60973 => -13882,
    60974 => -13879,
    60975 => -13876,
    60976 => -13873,
    60977 => -13870,
    60978 => -13868,
    60979 => -13865,
    60980 => -13862,
    60981 => -13859,
    60982 => -13856,
    60983 => -13853,
    60984 => -13850,
    60985 => -13848,
    60986 => -13845,
    60987 => -13842,
    60988 => -13839,
    60989 => -13836,
    60990 => -13833,
    60991 => -13831,
    60992 => -13828,
    60993 => -13825,
    60994 => -13822,
    60995 => -13819,
    60996 => -13816,
    60997 => -13813,
    60998 => -13811,
    60999 => -13808,
    61000 => -13805,
    61001 => -13802,
    61002 => -13799,
    61003 => -13796,
    61004 => -13793,
    61005 => -13791,
    61006 => -13788,
    61007 => -13785,
    61008 => -13782,
    61009 => -13779,
    61010 => -13776,
    61011 => -13774,
    61012 => -13771,
    61013 => -13768,
    61014 => -13765,
    61015 => -13762,
    61016 => -13759,
    61017 => -13756,
    61018 => -13754,
    61019 => -13751,
    61020 => -13748,
    61021 => -13745,
    61022 => -13742,
    61023 => -13739,
    61024 => -13736,
    61025 => -13734,
    61026 => -13731,
    61027 => -13728,
    61028 => -13725,
    61029 => -13722,
    61030 => -13719,
    61031 => -13717,
    61032 => -13714,
    61033 => -13711,
    61034 => -13708,
    61035 => -13705,
    61036 => -13702,
    61037 => -13699,
    61038 => -13697,
    61039 => -13694,
    61040 => -13691,
    61041 => -13688,
    61042 => -13685,
    61043 => -13682,
    61044 => -13679,
    61045 => -13677,
    61046 => -13674,
    61047 => -13671,
    61048 => -13668,
    61049 => -13665,
    61050 => -13662,
    61051 => -13659,
    61052 => -13657,
    61053 => -13654,
    61054 => -13651,
    61055 => -13648,
    61056 => -13645,
    61057 => -13642,
    61058 => -13639,
    61059 => -13637,
    61060 => -13634,
    61061 => -13631,
    61062 => -13628,
    61063 => -13625,
    61064 => -13622,
    61065 => -13619,
    61066 => -13617,
    61067 => -13614,
    61068 => -13611,
    61069 => -13608,
    61070 => -13605,
    61071 => -13602,
    61072 => -13599,
    61073 => -13597,
    61074 => -13594,
    61075 => -13591,
    61076 => -13588,
    61077 => -13585,
    61078 => -13582,
    61079 => -13579,
    61080 => -13577,
    61081 => -13574,
    61082 => -13571,
    61083 => -13568,
    61084 => -13565,
    61085 => -13562,
    61086 => -13559,
    61087 => -13557,
    61088 => -13554,
    61089 => -13551,
    61090 => -13548,
    61091 => -13545,
    61092 => -13542,
    61093 => -13539,
    61094 => -13537,
    61095 => -13534,
    61096 => -13531,
    61097 => -13528,
    61098 => -13525,
    61099 => -13522,
    61100 => -13519,
    61101 => -13516,
    61102 => -13514,
    61103 => -13511,
    61104 => -13508,
    61105 => -13505,
    61106 => -13502,
    61107 => -13499,
    61108 => -13496,
    61109 => -13494,
    61110 => -13491,
    61111 => -13488,
    61112 => -13485,
    61113 => -13482,
    61114 => -13479,
    61115 => -13476,
    61116 => -13474,
    61117 => -13471,
    61118 => -13468,
    61119 => -13465,
    61120 => -13462,
    61121 => -13459,
    61122 => -13456,
    61123 => -13454,
    61124 => -13451,
    61125 => -13448,
    61126 => -13445,
    61127 => -13442,
    61128 => -13439,
    61129 => -13436,
    61130 => -13433,
    61131 => -13431,
    61132 => -13428,
    61133 => -13425,
    61134 => -13422,
    61135 => -13419,
    61136 => -13416,
    61137 => -13413,
    61138 => -13411,
    61139 => -13408,
    61140 => -13405,
    61141 => -13402,
    61142 => -13399,
    61143 => -13396,
    61144 => -13393,
    61145 => -13390,
    61146 => -13388,
    61147 => -13385,
    61148 => -13382,
    61149 => -13379,
    61150 => -13376,
    61151 => -13373,
    61152 => -13370,
    61153 => -13368,
    61154 => -13365,
    61155 => -13362,
    61156 => -13359,
    61157 => -13356,
    61158 => -13353,
    61159 => -13350,
    61160 => -13347,
    61161 => -13345,
    61162 => -13342,
    61163 => -13339,
    61164 => -13336,
    61165 => -13333,
    61166 => -13330,
    61167 => -13327,
    61168 => -13324,
    61169 => -13322,
    61170 => -13319,
    61171 => -13316,
    61172 => -13313,
    61173 => -13310,
    61174 => -13307,
    61175 => -13304,
    61176 => -13302,
    61177 => -13299,
    61178 => -13296,
    61179 => -13293,
    61180 => -13290,
    61181 => -13287,
    61182 => -13284,
    61183 => -13281,
    61184 => -13279,
    61185 => -13276,
    61186 => -13273,
    61187 => -13270,
    61188 => -13267,
    61189 => -13264,
    61190 => -13261,
    61191 => -13258,
    61192 => -13256,
    61193 => -13253,
    61194 => -13250,
    61195 => -13247,
    61196 => -13244,
    61197 => -13241,
    61198 => -13238,
    61199 => -13235,
    61200 => -13233,
    61201 => -13230,
    61202 => -13227,
    61203 => -13224,
    61204 => -13221,
    61205 => -13218,
    61206 => -13215,
    61207 => -13212,
    61208 => -13210,
    61209 => -13207,
    61210 => -13204,
    61211 => -13201,
    61212 => -13198,
    61213 => -13195,
    61214 => -13192,
    61215 => -13189,
    61216 => -13187,
    61217 => -13184,
    61218 => -13181,
    61219 => -13178,
    61220 => -13175,
    61221 => -13172,
    61222 => -13169,
    61223 => -13166,
    61224 => -13164,
    61225 => -13161,
    61226 => -13158,
    61227 => -13155,
    61228 => -13152,
    61229 => -13149,
    61230 => -13146,
    61231 => -13143,
    61232 => -13141,
    61233 => -13138,
    61234 => -13135,
    61235 => -13132,
    61236 => -13129,
    61237 => -13126,
    61238 => -13123,
    61239 => -13120,
    61240 => -13118,
    61241 => -13115,
    61242 => -13112,
    61243 => -13109,
    61244 => -13106,
    61245 => -13103,
    61246 => -13100,
    61247 => -13097,
    61248 => -13094,
    61249 => -13092,
    61250 => -13089,
    61251 => -13086,
    61252 => -13083,
    61253 => -13080,
    61254 => -13077,
    61255 => -13074,
    61256 => -13071,
    61257 => -13069,
    61258 => -13066,
    61259 => -13063,
    61260 => -13060,
    61261 => -13057,
    61262 => -13054,
    61263 => -13051,
    61264 => -13048,
    61265 => -13046,
    61266 => -13043,
    61267 => -13040,
    61268 => -13037,
    61269 => -13034,
    61270 => -13031,
    61271 => -13028,
    61272 => -13025,
    61273 => -13022,
    61274 => -13020,
    61275 => -13017,
    61276 => -13014,
    61277 => -13011,
    61278 => -13008,
    61279 => -13005,
    61280 => -13002,
    61281 => -12999,
    61282 => -12997,
    61283 => -12994,
    61284 => -12991,
    61285 => -12988,
    61286 => -12985,
    61287 => -12982,
    61288 => -12979,
    61289 => -12976,
    61290 => -12973,
    61291 => -12971,
    61292 => -12968,
    61293 => -12965,
    61294 => -12962,
    61295 => -12959,
    61296 => -12956,
    61297 => -12953,
    61298 => -12950,
    61299 => -12947,
    61300 => -12945,
    61301 => -12942,
    61302 => -12939,
    61303 => -12936,
    61304 => -12933,
    61305 => -12930,
    61306 => -12927,
    61307 => -12924,
    61308 => -12921,
    61309 => -12919,
    61310 => -12916,
    61311 => -12913,
    61312 => -12910,
    61313 => -12907,
    61314 => -12904,
    61315 => -12901,
    61316 => -12898,
    61317 => -12895,
    61318 => -12893,
    61319 => -12890,
    61320 => -12887,
    61321 => -12884,
    61322 => -12881,
    61323 => -12878,
    61324 => -12875,
    61325 => -12872,
    61326 => -12870,
    61327 => -12867,
    61328 => -12864,
    61329 => -12861,
    61330 => -12858,
    61331 => -12855,
    61332 => -12852,
    61333 => -12849,
    61334 => -12846,
    61335 => -12843,
    61336 => -12841,
    61337 => -12838,
    61338 => -12835,
    61339 => -12832,
    61340 => -12829,
    61341 => -12826,
    61342 => -12823,
    61343 => -12820,
    61344 => -12817,
    61345 => -12815,
    61346 => -12812,
    61347 => -12809,
    61348 => -12806,
    61349 => -12803,
    61350 => -12800,
    61351 => -12797,
    61352 => -12794,
    61353 => -12791,
    61354 => -12789,
    61355 => -12786,
    61356 => -12783,
    61357 => -12780,
    61358 => -12777,
    61359 => -12774,
    61360 => -12771,
    61361 => -12768,
    61362 => -12765,
    61363 => -12763,
    61364 => -12760,
    61365 => -12757,
    61366 => -12754,
    61367 => -12751,
    61368 => -12748,
    61369 => -12745,
    61370 => -12742,
    61371 => -12739,
    61372 => -12736,
    61373 => -12734,
    61374 => -12731,
    61375 => -12728,
    61376 => -12725,
    61377 => -12722,
    61378 => -12719,
    61379 => -12716,
    61380 => -12713,
    61381 => -12710,
    61382 => -12708,
    61383 => -12705,
    61384 => -12702,
    61385 => -12699,
    61386 => -12696,
    61387 => -12693,
    61388 => -12690,
    61389 => -12687,
    61390 => -12684,
    61391 => -12681,
    61392 => -12679,
    61393 => -12676,
    61394 => -12673,
    61395 => -12670,
    61396 => -12667,
    61397 => -12664,
    61398 => -12661,
    61399 => -12658,
    61400 => -12655,
    61401 => -12652,
    61402 => -12650,
    61403 => -12647,
    61404 => -12644,
    61405 => -12641,
    61406 => -12638,
    61407 => -12635,
    61408 => -12632,
    61409 => -12629,
    61410 => -12626,
    61411 => -12624,
    61412 => -12621,
    61413 => -12618,
    61414 => -12615,
    61415 => -12612,
    61416 => -12609,
    61417 => -12606,
    61418 => -12603,
    61419 => -12600,
    61420 => -12597,
    61421 => -12595,
    61422 => -12592,
    61423 => -12589,
    61424 => -12586,
    61425 => -12583,
    61426 => -12580,
    61427 => -12577,
    61428 => -12574,
    61429 => -12571,
    61430 => -12568,
    61431 => -12566,
    61432 => -12563,
    61433 => -12560,
    61434 => -12557,
    61435 => -12554,
    61436 => -12551,
    61437 => -12548,
    61438 => -12545,
    61439 => -12542,
    61440 => -12539,
    61441 => -12536,
    61442 => -12534,
    61443 => -12531,
    61444 => -12528,
    61445 => -12525,
    61446 => -12522,
    61447 => -12519,
    61448 => -12516,
    61449 => -12513,
    61450 => -12510,
    61451 => -12507,
    61452 => -12505,
    61453 => -12502,
    61454 => -12499,
    61455 => -12496,
    61456 => -12493,
    61457 => -12490,
    61458 => -12487,
    61459 => -12484,
    61460 => -12481,
    61461 => -12478,
    61462 => -12476,
    61463 => -12473,
    61464 => -12470,
    61465 => -12467,
    61466 => -12464,
    61467 => -12461,
    61468 => -12458,
    61469 => -12455,
    61470 => -12452,
    61471 => -12449,
    61472 => -12446,
    61473 => -12444,
    61474 => -12441,
    61475 => -12438,
    61476 => -12435,
    61477 => -12432,
    61478 => -12429,
    61479 => -12426,
    61480 => -12423,
    61481 => -12420,
    61482 => -12417,
    61483 => -12414,
    61484 => -12412,
    61485 => -12409,
    61486 => -12406,
    61487 => -12403,
    61488 => -12400,
    61489 => -12397,
    61490 => -12394,
    61491 => -12391,
    61492 => -12388,
    61493 => -12385,
    61494 => -12382,
    61495 => -12380,
    61496 => -12377,
    61497 => -12374,
    61498 => -12371,
    61499 => -12368,
    61500 => -12365,
    61501 => -12362,
    61502 => -12359,
    61503 => -12356,
    61504 => -12353,
    61505 => -12350,
    61506 => -12348,
    61507 => -12345,
    61508 => -12342,
    61509 => -12339,
    61510 => -12336,
    61511 => -12333,
    61512 => -12330,
    61513 => -12327,
    61514 => -12324,
    61515 => -12321,
    61516 => -12318,
    61517 => -12316,
    61518 => -12313,
    61519 => -12310,
    61520 => -12307,
    61521 => -12304,
    61522 => -12301,
    61523 => -12298,
    61524 => -12295,
    61525 => -12292,
    61526 => -12289,
    61527 => -12286,
    61528 => -12284,
    61529 => -12281,
    61530 => -12278,
    61531 => -12275,
    61532 => -12272,
    61533 => -12269,
    61534 => -12266,
    61535 => -12263,
    61536 => -12260,
    61537 => -12257,
    61538 => -12254,
    61539 => -12251,
    61540 => -12249,
    61541 => -12246,
    61542 => -12243,
    61543 => -12240,
    61544 => -12237,
    61545 => -12234,
    61546 => -12231,
    61547 => -12228,
    61548 => -12225,
    61549 => -12222,
    61550 => -12219,
    61551 => -12217,
    61552 => -12214,
    61553 => -12211,
    61554 => -12208,
    61555 => -12205,
    61556 => -12202,
    61557 => -12199,
    61558 => -12196,
    61559 => -12193,
    61560 => -12190,
    61561 => -12187,
    61562 => -12184,
    61563 => -12182,
    61564 => -12179,
    61565 => -12176,
    61566 => -12173,
    61567 => -12170,
    61568 => -12167,
    61569 => -12164,
    61570 => -12161,
    61571 => -12158,
    61572 => -12155,
    61573 => -12152,
    61574 => -12149,
    61575 => -12147,
    61576 => -12144,
    61577 => -12141,
    61578 => -12138,
    61579 => -12135,
    61580 => -12132,
    61581 => -12129,
    61582 => -12126,
    61583 => -12123,
    61584 => -12120,
    61585 => -12117,
    61586 => -12114,
    61587 => -12112,
    61588 => -12109,
    61589 => -12106,
    61590 => -12103,
    61591 => -12100,
    61592 => -12097,
    61593 => -12094,
    61594 => -12091,
    61595 => -12088,
    61596 => -12085,
    61597 => -12082,
    61598 => -12079,
    61599 => -12076,
    61600 => -12074,
    61601 => -12071,
    61602 => -12068,
    61603 => -12065,
    61604 => -12062,
    61605 => -12059,
    61606 => -12056,
    61607 => -12053,
    61608 => -12050,
    61609 => -12047,
    61610 => -12044,
    61611 => -12041,
    61612 => -12038,
    61613 => -12036,
    61614 => -12033,
    61615 => -12030,
    61616 => -12027,
    61617 => -12024,
    61618 => -12021,
    61619 => -12018,
    61620 => -12015,
    61621 => -12012,
    61622 => -12009,
    61623 => -12006,
    61624 => -12003,
    61625 => -12001,
    61626 => -11998,
    61627 => -11995,
    61628 => -11992,
    61629 => -11989,
    61630 => -11986,
    61631 => -11983,
    61632 => -11980,
    61633 => -11977,
    61634 => -11974,
    61635 => -11971,
    61636 => -11968,
    61637 => -11965,
    61638 => -11962,
    61639 => -11960,
    61640 => -11957,
    61641 => -11954,
    61642 => -11951,
    61643 => -11948,
    61644 => -11945,
    61645 => -11942,
    61646 => -11939,
    61647 => -11936,
    61648 => -11933,
    61649 => -11930,
    61650 => -11927,
    61651 => -11924,
    61652 => -11922,
    61653 => -11919,
    61654 => -11916,
    61655 => -11913,
    61656 => -11910,
    61657 => -11907,
    61658 => -11904,
    61659 => -11901,
    61660 => -11898,
    61661 => -11895,
    61662 => -11892,
    61663 => -11889,
    61664 => -11886,
    61665 => -11883,
    61666 => -11881,
    61667 => -11878,
    61668 => -11875,
    61669 => -11872,
    61670 => -11869,
    61671 => -11866,
    61672 => -11863,
    61673 => -11860,
    61674 => -11857,
    61675 => -11854,
    61676 => -11851,
    61677 => -11848,
    61678 => -11845,
    61679 => -11842,
    61680 => -11840,
    61681 => -11837,
    61682 => -11834,
    61683 => -11831,
    61684 => -11828,
    61685 => -11825,
    61686 => -11822,
    61687 => -11819,
    61688 => -11816,
    61689 => -11813,
    61690 => -11810,
    61691 => -11807,
    61692 => -11804,
    61693 => -11801,
    61694 => -11799,
    61695 => -11796,
    61696 => -11793,
    61697 => -11790,
    61698 => -11787,
    61699 => -11784,
    61700 => -11781,
    61701 => -11778,
    61702 => -11775,
    61703 => -11772,
    61704 => -11769,
    61705 => -11766,
    61706 => -11763,
    61707 => -11760,
    61708 => -11758,
    61709 => -11755,
    61710 => -11752,
    61711 => -11749,
    61712 => -11746,
    61713 => -11743,
    61714 => -11740,
    61715 => -11737,
    61716 => -11734,
    61717 => -11731,
    61718 => -11728,
    61719 => -11725,
    61720 => -11722,
    61721 => -11719,
    61722 => -11716,
    61723 => -11714,
    61724 => -11711,
    61725 => -11708,
    61726 => -11705,
    61727 => -11702,
    61728 => -11699,
    61729 => -11696,
    61730 => -11693,
    61731 => -11690,
    61732 => -11687,
    61733 => -11684,
    61734 => -11681,
    61735 => -11678,
    61736 => -11675,
    61737 => -11672,
    61738 => -11669,
    61739 => -11667,
    61740 => -11664,
    61741 => -11661,
    61742 => -11658,
    61743 => -11655,
    61744 => -11652,
    61745 => -11649,
    61746 => -11646,
    61747 => -11643,
    61748 => -11640,
    61749 => -11637,
    61750 => -11634,
    61751 => -11631,
    61752 => -11628,
    61753 => -11625,
    61754 => -11623,
    61755 => -11620,
    61756 => -11617,
    61757 => -11614,
    61758 => -11611,
    61759 => -11608,
    61760 => -11605,
    61761 => -11602,
    61762 => -11599,
    61763 => -11596,
    61764 => -11593,
    61765 => -11590,
    61766 => -11587,
    61767 => -11584,
    61768 => -11581,
    61769 => -11578,
    61770 => -11575,
    61771 => -11573,
    61772 => -11570,
    61773 => -11567,
    61774 => -11564,
    61775 => -11561,
    61776 => -11558,
    61777 => -11555,
    61778 => -11552,
    61779 => -11549,
    61780 => -11546,
    61781 => -11543,
    61782 => -11540,
    61783 => -11537,
    61784 => -11534,
    61785 => -11531,
    61786 => -11528,
    61787 => -11526,
    61788 => -11523,
    61789 => -11520,
    61790 => -11517,
    61791 => -11514,
    61792 => -11511,
    61793 => -11508,
    61794 => -11505,
    61795 => -11502,
    61796 => -11499,
    61797 => -11496,
    61798 => -11493,
    61799 => -11490,
    61800 => -11487,
    61801 => -11484,
    61802 => -11481,
    61803 => -11478,
    61804 => -11476,
    61805 => -11473,
    61806 => -11470,
    61807 => -11467,
    61808 => -11464,
    61809 => -11461,
    61810 => -11458,
    61811 => -11455,
    61812 => -11452,
    61813 => -11449,
    61814 => -11446,
    61815 => -11443,
    61816 => -11440,
    61817 => -11437,
    61818 => -11434,
    61819 => -11431,
    61820 => -11428,
    61821 => -11425,
    61822 => -11423,
    61823 => -11420,
    61824 => -11417,
    61825 => -11414,
    61826 => -11411,
    61827 => -11408,
    61828 => -11405,
    61829 => -11402,
    61830 => -11399,
    61831 => -11396,
    61832 => -11393,
    61833 => -11390,
    61834 => -11387,
    61835 => -11384,
    61836 => -11381,
    61837 => -11378,
    61838 => -11375,
    61839 => -11372,
    61840 => -11370,
    61841 => -11367,
    61842 => -11364,
    61843 => -11361,
    61844 => -11358,
    61845 => -11355,
    61846 => -11352,
    61847 => -11349,
    61848 => -11346,
    61849 => -11343,
    61850 => -11340,
    61851 => -11337,
    61852 => -11334,
    61853 => -11331,
    61854 => -11328,
    61855 => -11325,
    61856 => -11322,
    61857 => -11319,
    61858 => -11316,
    61859 => -11314,
    61860 => -11311,
    61861 => -11308,
    61862 => -11305,
    61863 => -11302,
    61864 => -11299,
    61865 => -11296,
    61866 => -11293,
    61867 => -11290,
    61868 => -11287,
    61869 => -11284,
    61870 => -11281,
    61871 => -11278,
    61872 => -11275,
    61873 => -11272,
    61874 => -11269,
    61875 => -11266,
    61876 => -11263,
    61877 => -11260,
    61878 => -11257,
    61879 => -11255,
    61880 => -11252,
    61881 => -11249,
    61882 => -11246,
    61883 => -11243,
    61884 => -11240,
    61885 => -11237,
    61886 => -11234,
    61887 => -11231,
    61888 => -11228,
    61889 => -11225,
    61890 => -11222,
    61891 => -11219,
    61892 => -11216,
    61893 => -11213,
    61894 => -11210,
    61895 => -11207,
    61896 => -11204,
    61897 => -11201,
    61898 => -11198,
    61899 => -11195,
    61900 => -11193,
    61901 => -11190,
    61902 => -11187,
    61903 => -11184,
    61904 => -11181,
    61905 => -11178,
    61906 => -11175,
    61907 => -11172,
    61908 => -11169,
    61909 => -11166,
    61910 => -11163,
    61911 => -11160,
    61912 => -11157,
    61913 => -11154,
    61914 => -11151,
    61915 => -11148,
    61916 => -11145,
    61917 => -11142,
    61918 => -11139,
    61919 => -11136,
    61920 => -11133,
    61921 => -11131,
    61922 => -11128,
    61923 => -11125,
    61924 => -11122,
    61925 => -11119,
    61926 => -11116,
    61927 => -11113,
    61928 => -11110,
    61929 => -11107,
    61930 => -11104,
    61931 => -11101,
    61932 => -11098,
    61933 => -11095,
    61934 => -11092,
    61935 => -11089,
    61936 => -11086,
    61937 => -11083,
    61938 => -11080,
    61939 => -11077,
    61940 => -11074,
    61941 => -11071,
    61942 => -11068,
    61943 => -11065,
    61944 => -11063,
    61945 => -11060,
    61946 => -11057,
    61947 => -11054,
    61948 => -11051,
    61949 => -11048,
    61950 => -11045,
    61951 => -11042,
    61952 => -11039,
    61953 => -11036,
    61954 => -11033,
    61955 => -11030,
    61956 => -11027,
    61957 => -11024,
    61958 => -11021,
    61959 => -11018,
    61960 => -11015,
    61961 => -11012,
    61962 => -11009,
    61963 => -11006,
    61964 => -11003,
    61965 => -11000,
    61966 => -10997,
    61967 => -10994,
    61968 => -10992,
    61969 => -10989,
    61970 => -10986,
    61971 => -10983,
    61972 => -10980,
    61973 => -10977,
    61974 => -10974,
    61975 => -10971,
    61976 => -10968,
    61977 => -10965,
    61978 => -10962,
    61979 => -10959,
    61980 => -10956,
    61981 => -10953,
    61982 => -10950,
    61983 => -10947,
    61984 => -10944,
    61985 => -10941,
    61986 => -10938,
    61987 => -10935,
    61988 => -10932,
    61989 => -10929,
    61990 => -10926,
    61991 => -10923,
    61992 => -10920,
    61993 => -10918,
    61994 => -10915,
    61995 => -10912,
    61996 => -10909,
    61997 => -10906,
    61998 => -10903,
    61999 => -10900,
    62000 => -10897,
    62001 => -10894,
    62002 => -10891,
    62003 => -10888,
    62004 => -10885,
    62005 => -10882,
    62006 => -10879,
    62007 => -10876,
    62008 => -10873,
    62009 => -10870,
    62010 => -10867,
    62011 => -10864,
    62012 => -10861,
    62013 => -10858,
    62014 => -10855,
    62015 => -10852,
    62016 => -10849,
    62017 => -10846,
    62018 => -10843,
    62019 => -10840,
    62020 => -10838,
    62021 => -10835,
    62022 => -10832,
    62023 => -10829,
    62024 => -10826,
    62025 => -10823,
    62026 => -10820,
    62027 => -10817,
    62028 => -10814,
    62029 => -10811,
    62030 => -10808,
    62031 => -10805,
    62032 => -10802,
    62033 => -10799,
    62034 => -10796,
    62035 => -10793,
    62036 => -10790,
    62037 => -10787,
    62038 => -10784,
    62039 => -10781,
    62040 => -10778,
    62041 => -10775,
    62042 => -10772,
    62043 => -10769,
    62044 => -10766,
    62045 => -10763,
    62046 => -10760,
    62047 => -10757,
    62048 => -10754,
    62049 => -10751,
    62050 => -10749,
    62051 => -10746,
    62052 => -10743,
    62053 => -10740,
    62054 => -10737,
    62055 => -10734,
    62056 => -10731,
    62057 => -10728,
    62058 => -10725,
    62059 => -10722,
    62060 => -10719,
    62061 => -10716,
    62062 => -10713,
    62063 => -10710,
    62064 => -10707,
    62065 => -10704,
    62066 => -10701,
    62067 => -10698,
    62068 => -10695,
    62069 => -10692,
    62070 => -10689,
    62071 => -10686,
    62072 => -10683,
    62073 => -10680,
    62074 => -10677,
    62075 => -10674,
    62076 => -10671,
    62077 => -10668,
    62078 => -10665,
    62079 => -10662,
    62080 => -10659,
    62081 => -10656,
    62082 => -10654,
    62083 => -10651,
    62084 => -10648,
    62085 => -10645,
    62086 => -10642,
    62087 => -10639,
    62088 => -10636,
    62089 => -10633,
    62090 => -10630,
    62091 => -10627,
    62092 => -10624,
    62093 => -10621,
    62094 => -10618,
    62095 => -10615,
    62096 => -10612,
    62097 => -10609,
    62098 => -10606,
    62099 => -10603,
    62100 => -10600,
    62101 => -10597,
    62102 => -10594,
    62103 => -10591,
    62104 => -10588,
    62105 => -10585,
    62106 => -10582,
    62107 => -10579,
    62108 => -10576,
    62109 => -10573,
    62110 => -10570,
    62111 => -10567,
    62112 => -10564,
    62113 => -10561,
    62114 => -10558,
    62115 => -10555,
    62116 => -10552,
    62117 => -10549,
    62118 => -10546,
    62119 => -10544,
    62120 => -10541,
    62121 => -10538,
    62122 => -10535,
    62123 => -10532,
    62124 => -10529,
    62125 => -10526,
    62126 => -10523,
    62127 => -10520,
    62128 => -10517,
    62129 => -10514,
    62130 => -10511,
    62131 => -10508,
    62132 => -10505,
    62133 => -10502,
    62134 => -10499,
    62135 => -10496,
    62136 => -10493,
    62137 => -10490,
    62138 => -10487,
    62139 => -10484,
    62140 => -10481,
    62141 => -10478,
    62142 => -10475,
    62143 => -10472,
    62144 => -10469,
    62145 => -10466,
    62146 => -10463,
    62147 => -10460,
    62148 => -10457,
    62149 => -10454,
    62150 => -10451,
    62151 => -10448,
    62152 => -10445,
    62153 => -10442,
    62154 => -10439,
    62155 => -10436,
    62156 => -10433,
    62157 => -10430,
    62158 => -10427,
    62159 => -10424,
    62160 => -10421,
    62161 => -10419,
    62162 => -10416,
    62163 => -10413,
    62164 => -10410,
    62165 => -10407,
    62166 => -10404,
    62167 => -10401,
    62168 => -10398,
    62169 => -10395,
    62170 => -10392,
    62171 => -10389,
    62172 => -10386,
    62173 => -10383,
    62174 => -10380,
    62175 => -10377,
    62176 => -10374,
    62177 => -10371,
    62178 => -10368,
    62179 => -10365,
    62180 => -10362,
    62181 => -10359,
    62182 => -10356,
    62183 => -10353,
    62184 => -10350,
    62185 => -10347,
    62186 => -10344,
    62187 => -10341,
    62188 => -10338,
    62189 => -10335,
    62190 => -10332,
    62191 => -10329,
    62192 => -10326,
    62193 => -10323,
    62194 => -10320,
    62195 => -10317,
    62196 => -10314,
    62197 => -10311,
    62198 => -10308,
    62199 => -10305,
    62200 => -10302,
    62201 => -10299,
    62202 => -10296,
    62203 => -10293,
    62204 => -10290,
    62205 => -10287,
    62206 => -10284,
    62207 => -10281,
    62208 => -10278,
    62209 => -10275,
    62210 => -10272,
    62211 => -10269,
    62212 => -10266,
    62213 => -10263,
    62214 => -10261,
    62215 => -10258,
    62216 => -10255,
    62217 => -10252,
    62218 => -10249,
    62219 => -10246,
    62220 => -10243,
    62221 => -10240,
    62222 => -10237,
    62223 => -10234,
    62224 => -10231,
    62225 => -10228,
    62226 => -10225,
    62227 => -10222,
    62228 => -10219,
    62229 => -10216,
    62230 => -10213,
    62231 => -10210,
    62232 => -10207,
    62233 => -10204,
    62234 => -10201,
    62235 => -10198,
    62236 => -10195,
    62237 => -10192,
    62238 => -10189,
    62239 => -10186,
    62240 => -10183,
    62241 => -10180,
    62242 => -10177,
    62243 => -10174,
    62244 => -10171,
    62245 => -10168,
    62246 => -10165,
    62247 => -10162,
    62248 => -10159,
    62249 => -10156,
    62250 => -10153,
    62251 => -10150,
    62252 => -10147,
    62253 => -10144,
    62254 => -10141,
    62255 => -10138,
    62256 => -10135,
    62257 => -10132,
    62258 => -10129,
    62259 => -10126,
    62260 => -10123,
    62261 => -10120,
    62262 => -10117,
    62263 => -10114,
    62264 => -10111,
    62265 => -10108,
    62266 => -10105,
    62267 => -10102,
    62268 => -10099,
    62269 => -10096,
    62270 => -10093,
    62271 => -10090,
    62272 => -10087,
    62273 => -10084,
    62274 => -10081,
    62275 => -10078,
    62276 => -10075,
    62277 => -10072,
    62278 => -10069,
    62279 => -10066,
    62280 => -10063,
    62281 => -10060,
    62282 => -10057,
    62283 => -10054,
    62284 => -10051,
    62285 => -10048,
    62286 => -10045,
    62287 => -10042,
    62288 => -10039,
    62289 => -10036,
    62290 => -10033,
    62291 => -10031,
    62292 => -10028,
    62293 => -10025,
    62294 => -10022,
    62295 => -10019,
    62296 => -10016,
    62297 => -10013,
    62298 => -10010,
    62299 => -10007,
    62300 => -10004,
    62301 => -10001,
    62302 => -9998,
    62303 => -9995,
    62304 => -9992,
    62305 => -9989,
    62306 => -9986,
    62307 => -9983,
    62308 => -9980,
    62309 => -9977,
    62310 => -9974,
    62311 => -9971,
    62312 => -9968,
    62313 => -9965,
    62314 => -9962,
    62315 => -9959,
    62316 => -9956,
    62317 => -9953,
    62318 => -9950,
    62319 => -9947,
    62320 => -9944,
    62321 => -9941,
    62322 => -9938,
    62323 => -9935,
    62324 => -9932,
    62325 => -9929,
    62326 => -9926,
    62327 => -9923,
    62328 => -9920,
    62329 => -9917,
    62330 => -9914,
    62331 => -9911,
    62332 => -9908,
    62333 => -9905,
    62334 => -9902,
    62335 => -9899,
    62336 => -9896,
    62337 => -9893,
    62338 => -9890,
    62339 => -9887,
    62340 => -9884,
    62341 => -9881,
    62342 => -9878,
    62343 => -9875,
    62344 => -9872,
    62345 => -9869,
    62346 => -9866,
    62347 => -9863,
    62348 => -9860,
    62349 => -9857,
    62350 => -9854,
    62351 => -9851,
    62352 => -9848,
    62353 => -9845,
    62354 => -9842,
    62355 => -9839,
    62356 => -9836,
    62357 => -9833,
    62358 => -9830,
    62359 => -9827,
    62360 => -9824,
    62361 => -9821,
    62362 => -9818,
    62363 => -9815,
    62364 => -9812,
    62365 => -9809,
    62366 => -9806,
    62367 => -9803,
    62368 => -9800,
    62369 => -9797,
    62370 => -9794,
    62371 => -9791,
    62372 => -9788,
    62373 => -9785,
    62374 => -9782,
    62375 => -9779,
    62376 => -9776,
    62377 => -9773,
    62378 => -9770,
    62379 => -9767,
    62380 => -9764,
    62381 => -9761,
    62382 => -9758,
    62383 => -9755,
    62384 => -9752,
    62385 => -9749,
    62386 => -9746,
    62387 => -9743,
    62388 => -9740,
    62389 => -9737,
    62390 => -9734,
    62391 => -9731,
    62392 => -9728,
    62393 => -9725,
    62394 => -9722,
    62395 => -9719,
    62396 => -9716,
    62397 => -9713,
    62398 => -9710,
    62399 => -9707,
    62400 => -9704,
    62401 => -9701,
    62402 => -9698,
    62403 => -9695,
    62404 => -9692,
    62405 => -9689,
    62406 => -9686,
    62407 => -9683,
    62408 => -9680,
    62409 => -9677,
    62410 => -9674,
    62411 => -9671,
    62412 => -9668,
    62413 => -9665,
    62414 => -9662,
    62415 => -9659,
    62416 => -9656,
    62417 => -9653,
    62418 => -9650,
    62419 => -9647,
    62420 => -9644,
    62421 => -9641,
    62422 => -9638,
    62423 => -9635,
    62424 => -9632,
    62425 => -9629,
    62426 => -9626,
    62427 => -9623,
    62428 => -9620,
    62429 => -9617,
    62430 => -9614,
    62431 => -9611,
    62432 => -9608,
    62433 => -9605,
    62434 => -9602,
    62435 => -9599,
    62436 => -9596,
    62437 => -9593,
    62438 => -9590,
    62439 => -9587,
    62440 => -9584,
    62441 => -9581,
    62442 => -9578,
    62443 => -9575,
    62444 => -9572,
    62445 => -9569,
    62446 => -9566,
    62447 => -9563,
    62448 => -9560,
    62449 => -9557,
    62450 => -9554,
    62451 => -9551,
    62452 => -9548,
    62453 => -9545,
    62454 => -9542,
    62455 => -9539,
    62456 => -9536,
    62457 => -9533,
    62458 => -9530,
    62459 => -9527,
    62460 => -9524,
    62461 => -9521,
    62462 => -9518,
    62463 => -9515,
    62464 => -9512,
    62465 => -9509,
    62466 => -9506,
    62467 => -9503,
    62468 => -9500,
    62469 => -9497,
    62470 => -9494,
    62471 => -9491,
    62472 => -9488,
    62473 => -9485,
    62474 => -9482,
    62475 => -9479,
    62476 => -9476,
    62477 => -9473,
    62478 => -9470,
    62479 => -9467,
    62480 => -9464,
    62481 => -9461,
    62482 => -9458,
    62483 => -9455,
    62484 => -9452,
    62485 => -9449,
    62486 => -9446,
    62487 => -9443,
    62488 => -9440,
    62489 => -9437,
    62490 => -9434,
    62491 => -9431,
    62492 => -9428,
    62493 => -9425,
    62494 => -9422,
    62495 => -9419,
    62496 => -9416,
    62497 => -9413,
    62498 => -9409,
    62499 => -9406,
    62500 => -9403,
    62501 => -9400,
    62502 => -9397,
    62503 => -9394,
    62504 => -9391,
    62505 => -9388,
    62506 => -9385,
    62507 => -9382,
    62508 => -9379,
    62509 => -9376,
    62510 => -9373,
    62511 => -9370,
    62512 => -9367,
    62513 => -9364,
    62514 => -9361,
    62515 => -9358,
    62516 => -9355,
    62517 => -9352,
    62518 => -9349,
    62519 => -9346,
    62520 => -9343,
    62521 => -9340,
    62522 => -9337,
    62523 => -9334,
    62524 => -9331,
    62525 => -9328,
    62526 => -9325,
    62527 => -9322,
    62528 => -9319,
    62529 => -9316,
    62530 => -9313,
    62531 => -9310,
    62532 => -9307,
    62533 => -9304,
    62534 => -9301,
    62535 => -9298,
    62536 => -9295,
    62537 => -9292,
    62538 => -9289,
    62539 => -9286,
    62540 => -9283,
    62541 => -9280,
    62542 => -9277,
    62543 => -9274,
    62544 => -9271,
    62545 => -9268,
    62546 => -9265,
    62547 => -9262,
    62548 => -9259,
    62549 => -9256,
    62550 => -9253,
    62551 => -9250,
    62552 => -9247,
    62553 => -9244,
    62554 => -9241,
    62555 => -9238,
    62556 => -9235,
    62557 => -9232,
    62558 => -9229,
    62559 => -9226,
    62560 => -9223,
    62561 => -9220,
    62562 => -9217,
    62563 => -9214,
    62564 => -9211,
    62565 => -9208,
    62566 => -9205,
    62567 => -9202,
    62568 => -9199,
    62569 => -9196,
    62570 => -9193,
    62571 => -9190,
    62572 => -9187,
    62573 => -9184,
    62574 => -9181,
    62575 => -9178,
    62576 => -9175,
    62577 => -9172,
    62578 => -9168,
    62579 => -9165,
    62580 => -9162,
    62581 => -9159,
    62582 => -9156,
    62583 => -9153,
    62584 => -9150,
    62585 => -9147,
    62586 => -9144,
    62587 => -9141,
    62588 => -9138,
    62589 => -9135,
    62590 => -9132,
    62591 => -9129,
    62592 => -9126,
    62593 => -9123,
    62594 => -9120,
    62595 => -9117,
    62596 => -9114,
    62597 => -9111,
    62598 => -9108,
    62599 => -9105,
    62600 => -9102,
    62601 => -9099,
    62602 => -9096,
    62603 => -9093,
    62604 => -9090,
    62605 => -9087,
    62606 => -9084,
    62607 => -9081,
    62608 => -9078,
    62609 => -9075,
    62610 => -9072,
    62611 => -9069,
    62612 => -9066,
    62613 => -9063,
    62614 => -9060,
    62615 => -9057,
    62616 => -9054,
    62617 => -9051,
    62618 => -9048,
    62619 => -9045,
    62620 => -9042,
    62621 => -9039,
    62622 => -9036,
    62623 => -9033,
    62624 => -9030,
    62625 => -9027,
    62626 => -9024,
    62627 => -9021,
    62628 => -9018,
    62629 => -9015,
    62630 => -9012,
    62631 => -9009,
    62632 => -9006,
    62633 => -9002,
    62634 => -8999,
    62635 => -8996,
    62636 => -8993,
    62637 => -8990,
    62638 => -8987,
    62639 => -8984,
    62640 => -8981,
    62641 => -8978,
    62642 => -8975,
    62643 => -8972,
    62644 => -8969,
    62645 => -8966,
    62646 => -8963,
    62647 => -8960,
    62648 => -8957,
    62649 => -8954,
    62650 => -8951,
    62651 => -8948,
    62652 => -8945,
    62653 => -8942,
    62654 => -8939,
    62655 => -8936,
    62656 => -8933,
    62657 => -8930,
    62658 => -8927,
    62659 => -8924,
    62660 => -8921,
    62661 => -8918,
    62662 => -8915,
    62663 => -8912,
    62664 => -8909,
    62665 => -8906,
    62666 => -8903,
    62667 => -8900,
    62668 => -8897,
    62669 => -8894,
    62670 => -8891,
    62671 => -8888,
    62672 => -8885,
    62673 => -8882,
    62674 => -8879,
    62675 => -8876,
    62676 => -8873,
    62677 => -8869,
    62678 => -8866,
    62679 => -8863,
    62680 => -8860,
    62681 => -8857,
    62682 => -8854,
    62683 => -8851,
    62684 => -8848,
    62685 => -8845,
    62686 => -8842,
    62687 => -8839,
    62688 => -8836,
    62689 => -8833,
    62690 => -8830,
    62691 => -8827,
    62692 => -8824,
    62693 => -8821,
    62694 => -8818,
    62695 => -8815,
    62696 => -8812,
    62697 => -8809,
    62698 => -8806,
    62699 => -8803,
    62700 => -8800,
    62701 => -8797,
    62702 => -8794,
    62703 => -8791,
    62704 => -8788,
    62705 => -8785,
    62706 => -8782,
    62707 => -8779,
    62708 => -8776,
    62709 => -8773,
    62710 => -8770,
    62711 => -8767,
    62712 => -8764,
    62713 => -8761,
    62714 => -8758,
    62715 => -8755,
    62716 => -8751,
    62717 => -8748,
    62718 => -8745,
    62719 => -8742,
    62720 => -8739,
    62721 => -8736,
    62722 => -8733,
    62723 => -8730,
    62724 => -8727,
    62725 => -8724,
    62726 => -8721,
    62727 => -8718,
    62728 => -8715,
    62729 => -8712,
    62730 => -8709,
    62731 => -8706,
    62732 => -8703,
    62733 => -8700,
    62734 => -8697,
    62735 => -8694,
    62736 => -8691,
    62737 => -8688,
    62738 => -8685,
    62739 => -8682,
    62740 => -8679,
    62741 => -8676,
    62742 => -8673,
    62743 => -8670,
    62744 => -8667,
    62745 => -8664,
    62746 => -8661,
    62747 => -8658,
    62748 => -8655,
    62749 => -8652,
    62750 => -8649,
    62751 => -8645,
    62752 => -8642,
    62753 => -8639,
    62754 => -8636,
    62755 => -8633,
    62756 => -8630,
    62757 => -8627,
    62758 => -8624,
    62759 => -8621,
    62760 => -8618,
    62761 => -8615,
    62762 => -8612,
    62763 => -8609,
    62764 => -8606,
    62765 => -8603,
    62766 => -8600,
    62767 => -8597,
    62768 => -8594,
    62769 => -8591,
    62770 => -8588,
    62771 => -8585,
    62772 => -8582,
    62773 => -8579,
    62774 => -8576,
    62775 => -8573,
    62776 => -8570,
    62777 => -8567,
    62778 => -8564,
    62779 => -8561,
    62780 => -8558,
    62781 => -8555,
    62782 => -8552,
    62783 => -8548,
    62784 => -8545,
    62785 => -8542,
    62786 => -8539,
    62787 => -8536,
    62788 => -8533,
    62789 => -8530,
    62790 => -8527,
    62791 => -8524,
    62792 => -8521,
    62793 => -8518,
    62794 => -8515,
    62795 => -8512,
    62796 => -8509,
    62797 => -8506,
    62798 => -8503,
    62799 => -8500,
    62800 => -8497,
    62801 => -8494,
    62802 => -8491,
    62803 => -8488,
    62804 => -8485,
    62805 => -8482,
    62806 => -8479,
    62807 => -8476,
    62808 => -8473,
    62809 => -8470,
    62810 => -8467,
    62811 => -8464,
    62812 => -8460,
    62813 => -8457,
    62814 => -8454,
    62815 => -8451,
    62816 => -8448,
    62817 => -8445,
    62818 => -8442,
    62819 => -8439,
    62820 => -8436,
    62821 => -8433,
    62822 => -8430,
    62823 => -8427,
    62824 => -8424,
    62825 => -8421,
    62826 => -8418,
    62827 => -8415,
    62828 => -8412,
    62829 => -8409,
    62830 => -8406,
    62831 => -8403,
    62832 => -8400,
    62833 => -8397,
    62834 => -8394,
    62835 => -8391,
    62836 => -8388,
    62837 => -8385,
    62838 => -8382,
    62839 => -8379,
    62840 => -8375,
    62841 => -8372,
    62842 => -8369,
    62843 => -8366,
    62844 => -8363,
    62845 => -8360,
    62846 => -8357,
    62847 => -8354,
    62848 => -8351,
    62849 => -8348,
    62850 => -8345,
    62851 => -8342,
    62852 => -8339,
    62853 => -8336,
    62854 => -8333,
    62855 => -8330,
    62856 => -8327,
    62857 => -8324,
    62858 => -8321,
    62859 => -8318,
    62860 => -8315,
    62861 => -8312,
    62862 => -8309,
    62863 => -8306,
    62864 => -8303,
    62865 => -8300,
    62866 => -8296,
    62867 => -8293,
    62868 => -8290,
    62869 => -8287,
    62870 => -8284,
    62871 => -8281,
    62872 => -8278,
    62873 => -8275,
    62874 => -8272,
    62875 => -8269,
    62876 => -8266,
    62877 => -8263,
    62878 => -8260,
    62879 => -8257,
    62880 => -8254,
    62881 => -8251,
    62882 => -8248,
    62883 => -8245,
    62884 => -8242,
    62885 => -8239,
    62886 => -8236,
    62887 => -8233,
    62888 => -8230,
    62889 => -8227,
    62890 => -8224,
    62891 => -8220,
    62892 => -8217,
    62893 => -8214,
    62894 => -8211,
    62895 => -8208,
    62896 => -8205,
    62897 => -8202,
    62898 => -8199,
    62899 => -8196,
    62900 => -8193,
    62901 => -8190,
    62902 => -8187,
    62903 => -8184,
    62904 => -8181,
    62905 => -8178,
    62906 => -8175,
    62907 => -8172,
    62908 => -8169,
    62909 => -8166,
    62910 => -8163,
    62911 => -8160,
    62912 => -8157,
    62913 => -8154,
    62914 => -8151,
    62915 => -8147,
    62916 => -8144,
    62917 => -8141,
    62918 => -8138,
    62919 => -8135,
    62920 => -8132,
    62921 => -8129,
    62922 => -8126,
    62923 => -8123,
    62924 => -8120,
    62925 => -8117,
    62926 => -8114,
    62927 => -8111,
    62928 => -8108,
    62929 => -8105,
    62930 => -8102,
    62931 => -8099,
    62932 => -8096,
    62933 => -8093,
    62934 => -8090,
    62935 => -8087,
    62936 => -8084,
    62937 => -8081,
    62938 => -8077,
    62939 => -8074,
    62940 => -8071,
    62941 => -8068,
    62942 => -8065,
    62943 => -8062,
    62944 => -8059,
    62945 => -8056,
    62946 => -8053,
    62947 => -8050,
    62948 => -8047,
    62949 => -8044,
    62950 => -8041,
    62951 => -8038,
    62952 => -8035,
    62953 => -8032,
    62954 => -8029,
    62955 => -8026,
    62956 => -8023,
    62957 => -8020,
    62958 => -8017,
    62959 => -8014,
    62960 => -8010,
    62961 => -8007,
    62962 => -8004,
    62963 => -8001,
    62964 => -7998,
    62965 => -7995,
    62966 => -7992,
    62967 => -7989,
    62968 => -7986,
    62969 => -7983,
    62970 => -7980,
    62971 => -7977,
    62972 => -7974,
    62973 => -7971,
    62974 => -7968,
    62975 => -7965,
    62976 => -7962,
    62977 => -7959,
    62978 => -7956,
    62979 => -7953,
    62980 => -7950,
    62981 => -7946,
    62982 => -7943,
    62983 => -7940,
    62984 => -7937,
    62985 => -7934,
    62986 => -7931,
    62987 => -7928,
    62988 => -7925,
    62989 => -7922,
    62990 => -7919,
    62991 => -7916,
    62992 => -7913,
    62993 => -7910,
    62994 => -7907,
    62995 => -7904,
    62996 => -7901,
    62997 => -7898,
    62998 => -7895,
    62999 => -7892,
    63000 => -7889,
    63001 => -7886,
    63002 => -7882,
    63003 => -7879,
    63004 => -7876,
    63005 => -7873,
    63006 => -7870,
    63007 => -7867,
    63008 => -7864,
    63009 => -7861,
    63010 => -7858,
    63011 => -7855,
    63012 => -7852,
    63013 => -7849,
    63014 => -7846,
    63015 => -7843,
    63016 => -7840,
    63017 => -7837,
    63018 => -7834,
    63019 => -7831,
    63020 => -7828,
    63021 => -7825,
    63022 => -7821,
    63023 => -7818,
    63024 => -7815,
    63025 => -7812,
    63026 => -7809,
    63027 => -7806,
    63028 => -7803,
    63029 => -7800,
    63030 => -7797,
    63031 => -7794,
    63032 => -7791,
    63033 => -7788,
    63034 => -7785,
    63035 => -7782,
    63036 => -7779,
    63037 => -7776,
    63038 => -7773,
    63039 => -7770,
    63040 => -7767,
    63041 => -7764,
    63042 => -7760,
    63043 => -7757,
    63044 => -7754,
    63045 => -7751,
    63046 => -7748,
    63047 => -7745,
    63048 => -7742,
    63049 => -7739,
    63050 => -7736,
    63051 => -7733,
    63052 => -7730,
    63053 => -7727,
    63054 => -7724,
    63055 => -7721,
    63056 => -7718,
    63057 => -7715,
    63058 => -7712,
    63059 => -7709,
    63060 => -7705,
    63061 => -7702,
    63062 => -7699,
    63063 => -7696,
    63064 => -7693,
    63065 => -7690,
    63066 => -7687,
    63067 => -7684,
    63068 => -7681,
    63069 => -7678,
    63070 => -7675,
    63071 => -7672,
    63072 => -7669,
    63073 => -7666,
    63074 => -7663,
    63075 => -7660,
    63076 => -7657,
    63077 => -7654,
    63078 => -7651,
    63079 => -7647,
    63080 => -7644,
    63081 => -7641,
    63082 => -7638,
    63083 => -7635,
    63084 => -7632,
    63085 => -7629,
    63086 => -7626,
    63087 => -7623,
    63088 => -7620,
    63089 => -7617,
    63090 => -7614,
    63091 => -7611,
    63092 => -7608,
    63093 => -7605,
    63094 => -7602,
    63095 => -7599,
    63096 => -7596,
    63097 => -7592,
    63098 => -7589,
    63099 => -7586,
    63100 => -7583,
    63101 => -7580,
    63102 => -7577,
    63103 => -7574,
    63104 => -7571,
    63105 => -7568,
    63106 => -7565,
    63107 => -7562,
    63108 => -7559,
    63109 => -7556,
    63110 => -7553,
    63111 => -7550,
    63112 => -7547,
    63113 => -7544,
    63114 => -7541,
    63115 => -7537,
    63116 => -7534,
    63117 => -7531,
    63118 => -7528,
    63119 => -7525,
    63120 => -7522,
    63121 => -7519,
    63122 => -7516,
    63123 => -7513,
    63124 => -7510,
    63125 => -7507,
    63126 => -7504,
    63127 => -7501,
    63128 => -7498,
    63129 => -7495,
    63130 => -7492,
    63131 => -7489,
    63132 => -7485,
    63133 => -7482,
    63134 => -7479,
    63135 => -7476,
    63136 => -7473,
    63137 => -7470,
    63138 => -7467,
    63139 => -7464,
    63140 => -7461,
    63141 => -7458,
    63142 => -7455,
    63143 => -7452,
    63144 => -7449,
    63145 => -7446,
    63146 => -7443,
    63147 => -7440,
    63148 => -7437,
    63149 => -7433,
    63150 => -7430,
    63151 => -7427,
    63152 => -7424,
    63153 => -7421,
    63154 => -7418,
    63155 => -7415,
    63156 => -7412,
    63157 => -7409,
    63158 => -7406,
    63159 => -7403,
    63160 => -7400,
    63161 => -7397,
    63162 => -7394,
    63163 => -7391,
    63164 => -7388,
    63165 => -7385,
    63166 => -7381,
    63167 => -7378,
    63168 => -7375,
    63169 => -7372,
    63170 => -7369,
    63171 => -7366,
    63172 => -7363,
    63173 => -7360,
    63174 => -7357,
    63175 => -7354,
    63176 => -7351,
    63177 => -7348,
    63178 => -7345,
    63179 => -7342,
    63180 => -7339,
    63181 => -7336,
    63182 => -7332,
    63183 => -7329,
    63184 => -7326,
    63185 => -7323,
    63186 => -7320,
    63187 => -7317,
    63188 => -7314,
    63189 => -7311,
    63190 => -7308,
    63191 => -7305,
    63192 => -7302,
    63193 => -7299,
    63194 => -7296,
    63195 => -7293,
    63196 => -7290,
    63197 => -7287,
    63198 => -7283,
    63199 => -7280,
    63200 => -7277,
    63201 => -7274,
    63202 => -7271,
    63203 => -7268,
    63204 => -7265,
    63205 => -7262,
    63206 => -7259,
    63207 => -7256,
    63208 => -7253,
    63209 => -7250,
    63210 => -7247,
    63211 => -7244,
    63212 => -7241,
    63213 => -7238,
    63214 => -7234,
    63215 => -7231,
    63216 => -7228,
    63217 => -7225,
    63218 => -7222,
    63219 => -7219,
    63220 => -7216,
    63221 => -7213,
    63222 => -7210,
    63223 => -7207,
    63224 => -7204,
    63225 => -7201,
    63226 => -7198,
    63227 => -7195,
    63228 => -7192,
    63229 => -7188,
    63230 => -7185,
    63231 => -7182,
    63232 => -7179,
    63233 => -7176,
    63234 => -7173,
    63235 => -7170,
    63236 => -7167,
    63237 => -7164,
    63238 => -7161,
    63239 => -7158,
    63240 => -7155,
    63241 => -7152,
    63242 => -7149,
    63243 => -7146,
    63244 => -7143,
    63245 => -7139,
    63246 => -7136,
    63247 => -7133,
    63248 => -7130,
    63249 => -7127,
    63250 => -7124,
    63251 => -7121,
    63252 => -7118,
    63253 => -7115,
    63254 => -7112,
    63255 => -7109,
    63256 => -7106,
    63257 => -7103,
    63258 => -7100,
    63259 => -7097,
    63260 => -7093,
    63261 => -7090,
    63262 => -7087,
    63263 => -7084,
    63264 => -7081,
    63265 => -7078,
    63266 => -7075,
    63267 => -7072,
    63268 => -7069,
    63269 => -7066,
    63270 => -7063,
    63271 => -7060,
    63272 => -7057,
    63273 => -7054,
    63274 => -7050,
    63275 => -7047,
    63276 => -7044,
    63277 => -7041,
    63278 => -7038,
    63279 => -7035,
    63280 => -7032,
    63281 => -7029,
    63282 => -7026,
    63283 => -7023,
    63284 => -7020,
    63285 => -7017,
    63286 => -7014,
    63287 => -7011,
    63288 => -7008,
    63289 => -7004,
    63290 => -7001,
    63291 => -6998,
    63292 => -6995,
    63293 => -6992,
    63294 => -6989,
    63295 => -6986,
    63296 => -6983,
    63297 => -6980,
    63298 => -6977,
    63299 => -6974,
    63300 => -6971,
    63301 => -6968,
    63302 => -6965,
    63303 => -6961,
    63304 => -6958,
    63305 => -6955,
    63306 => -6952,
    63307 => -6949,
    63308 => -6946,
    63309 => -6943,
    63310 => -6940,
    63311 => -6937,
    63312 => -6934,
    63313 => -6931,
    63314 => -6928,
    63315 => -6925,
    63316 => -6922,
    63317 => -6919,
    63318 => -6915,
    63319 => -6912,
    63320 => -6909,
    63321 => -6906,
    63322 => -6903,
    63323 => -6900,
    63324 => -6897,
    63325 => -6894,
    63326 => -6891,
    63327 => -6888,
    63328 => -6885,
    63329 => -6882,
    63330 => -6879,
    63331 => -6876,
    63332 => -6872,
    63333 => -6869,
    63334 => -6866,
    63335 => -6863,
    63336 => -6860,
    63337 => -6857,
    63338 => -6854,
    63339 => -6851,
    63340 => -6848,
    63341 => -6845,
    63342 => -6842,
    63343 => -6839,
    63344 => -6836,
    63345 => -6833,
    63346 => -6829,
    63347 => -6826,
    63348 => -6823,
    63349 => -6820,
    63350 => -6817,
    63351 => -6814,
    63352 => -6811,
    63353 => -6808,
    63354 => -6805,
    63355 => -6802,
    63356 => -6799,
    63357 => -6796,
    63358 => -6793,
    63359 => -6789,
    63360 => -6786,
    63361 => -6783,
    63362 => -6780,
    63363 => -6777,
    63364 => -6774,
    63365 => -6771,
    63366 => -6768,
    63367 => -6765,
    63368 => -6762,
    63369 => -6759,
    63370 => -6756,
    63371 => -6753,
    63372 => -6750,
    63373 => -6746,
    63374 => -6743,
    63375 => -6740,
    63376 => -6737,
    63377 => -6734,
    63378 => -6731,
    63379 => -6728,
    63380 => -6725,
    63381 => -6722,
    63382 => -6719,
    63383 => -6716,
    63384 => -6713,
    63385 => -6710,
    63386 => -6706,
    63387 => -6703,
    63388 => -6700,
    63389 => -6697,
    63390 => -6694,
    63391 => -6691,
    63392 => -6688,
    63393 => -6685,
    63394 => -6682,
    63395 => -6679,
    63396 => -6676,
    63397 => -6673,
    63398 => -6670,
    63399 => -6667,
    63400 => -6663,
    63401 => -6660,
    63402 => -6657,
    63403 => -6654,
    63404 => -6651,
    63405 => -6648,
    63406 => -6645,
    63407 => -6642,
    63408 => -6639,
    63409 => -6636,
    63410 => -6633,
    63411 => -6630,
    63412 => -6627,
    63413 => -6623,
    63414 => -6620,
    63415 => -6617,
    63416 => -6614,
    63417 => -6611,
    63418 => -6608,
    63419 => -6605,
    63420 => -6602,
    63421 => -6599,
    63422 => -6596,
    63423 => -6593,
    63424 => -6590,
    63425 => -6587,
    63426 => -6583,
    63427 => -6580,
    63428 => -6577,
    63429 => -6574,
    63430 => -6571,
    63431 => -6568,
    63432 => -6565,
    63433 => -6562,
    63434 => -6559,
    63435 => -6556,
    63436 => -6553,
    63437 => -6550,
    63438 => -6547,
    63439 => -6543,
    63440 => -6540,
    63441 => -6537,
    63442 => -6534,
    63443 => -6531,
    63444 => -6528,
    63445 => -6525,
    63446 => -6522,
    63447 => -6519,
    63448 => -6516,
    63449 => -6513,
    63450 => -6510,
    63451 => -6506,
    63452 => -6503,
    63453 => -6500,
    63454 => -6497,
    63455 => -6494,
    63456 => -6491,
    63457 => -6488,
    63458 => -6485,
    63459 => -6482,
    63460 => -6479,
    63461 => -6476,
    63462 => -6473,
    63463 => -6470,
    63464 => -6466,
    63465 => -6463,
    63466 => -6460,
    63467 => -6457,
    63468 => -6454,
    63469 => -6451,
    63470 => -6448,
    63471 => -6445,
    63472 => -6442,
    63473 => -6439,
    63474 => -6436,
    63475 => -6433,
    63476 => -6429,
    63477 => -6426,
    63478 => -6423,
    63479 => -6420,
    63480 => -6417,
    63481 => -6414,
    63482 => -6411,
    63483 => -6408,
    63484 => -6405,
    63485 => -6402,
    63486 => -6399,
    63487 => -6396,
    63488 => -6393,
    63489 => -6389,
    63490 => -6386,
    63491 => -6383,
    63492 => -6380,
    63493 => -6377,
    63494 => -6374,
    63495 => -6371,
    63496 => -6368,
    63497 => -6365,
    63498 => -6362,
    63499 => -6359,
    63500 => -6356,
    63501 => -6352,
    63502 => -6349,
    63503 => -6346,
    63504 => -6343,
    63505 => -6340,
    63506 => -6337,
    63507 => -6334,
    63508 => -6331,
    63509 => -6328,
    63510 => -6325,
    63511 => -6322,
    63512 => -6319,
    63513 => -6315,
    63514 => -6312,
    63515 => -6309,
    63516 => -6306,
    63517 => -6303,
    63518 => -6300,
    63519 => -6297,
    63520 => -6294,
    63521 => -6291,
    63522 => -6288,
    63523 => -6285,
    63524 => -6282,
    63525 => -6278,
    63526 => -6275,
    63527 => -6272,
    63528 => -6269,
    63529 => -6266,
    63530 => -6263,
    63531 => -6260,
    63532 => -6257,
    63533 => -6254,
    63534 => -6251,
    63535 => -6248,
    63536 => -6245,
    63537 => -6241,
    63538 => -6238,
    63539 => -6235,
    63540 => -6232,
    63541 => -6229,
    63542 => -6226,
    63543 => -6223,
    63544 => -6220,
    63545 => -6217,
    63546 => -6214,
    63547 => -6211,
    63548 => -6208,
    63549 => -6204,
    63550 => -6201,
    63551 => -6198,
    63552 => -6195,
    63553 => -6192,
    63554 => -6189,
    63555 => -6186,
    63556 => -6183,
    63557 => -6180,
    63558 => -6177,
    63559 => -6174,
    63560 => -6171,
    63561 => -6167,
    63562 => -6164,
    63563 => -6161,
    63564 => -6158,
    63565 => -6155,
    63566 => -6152,
    63567 => -6149,
    63568 => -6146,
    63569 => -6143,
    63570 => -6140,
    63571 => -6137,
    63572 => -6134,
    63573 => -6130,
    63574 => -6127,
    63575 => -6124,
    63576 => -6121,
    63577 => -6118,
    63578 => -6115,
    63579 => -6112,
    63580 => -6109,
    63581 => -6106,
    63582 => -6103,
    63583 => -6100,
    63584 => -6096,
    63585 => -6093,
    63586 => -6090,
    63587 => -6087,
    63588 => -6084,
    63589 => -6081,
    63590 => -6078,
    63591 => -6075,
    63592 => -6072,
    63593 => -6069,
    63594 => -6066,
    63595 => -6063,
    63596 => -6059,
    63597 => -6056,
    63598 => -6053,
    63599 => -6050,
    63600 => -6047,
    63601 => -6044,
    63602 => -6041,
    63603 => -6038,
    63604 => -6035,
    63605 => -6032,
    63606 => -6029,
    63607 => -6025,
    63608 => -6022,
    63609 => -6019,
    63610 => -6016,
    63611 => -6013,
    63612 => -6010,
    63613 => -6007,
    63614 => -6004,
    63615 => -6001,
    63616 => -5998,
    63617 => -5995,
    63618 => -5991,
    63619 => -5988,
    63620 => -5985,
    63621 => -5982,
    63622 => -5979,
    63623 => -5976,
    63624 => -5973,
    63625 => -5970,
    63626 => -5967,
    63627 => -5964,
    63628 => -5961,
    63629 => -5958,
    63630 => -5954,
    63631 => -5951,
    63632 => -5948,
    63633 => -5945,
    63634 => -5942,
    63635 => -5939,
    63636 => -5936,
    63637 => -5933,
    63638 => -5930,
    63639 => -5927,
    63640 => -5924,
    63641 => -5920,
    63642 => -5917,
    63643 => -5914,
    63644 => -5911,
    63645 => -5908,
    63646 => -5905,
    63647 => -5902,
    63648 => -5899,
    63649 => -5896,
    63650 => -5893,
    63651 => -5890,
    63652 => -5886,
    63653 => -5883,
    63654 => -5880,
    63655 => -5877,
    63656 => -5874,
    63657 => -5871,
    63658 => -5868,
    63659 => -5865,
    63660 => -5862,
    63661 => -5859,
    63662 => -5856,
    63663 => -5852,
    63664 => -5849,
    63665 => -5846,
    63666 => -5843,
    63667 => -5840,
    63668 => -5837,
    63669 => -5834,
    63670 => -5831,
    63671 => -5828,
    63672 => -5825,
    63673 => -5822,
    63674 => -5818,
    63675 => -5815,
    63676 => -5812,
    63677 => -5809,
    63678 => -5806,
    63679 => -5803,
    63680 => -5800,
    63681 => -5797,
    63682 => -5794,
    63683 => -5791,
    63684 => -5788,
    63685 => -5784,
    63686 => -5781,
    63687 => -5778,
    63688 => -5775,
    63689 => -5772,
    63690 => -5769,
    63691 => -5766,
    63692 => -5763,
    63693 => -5760,
    63694 => -5757,
    63695 => -5754,
    63696 => -5750,
    63697 => -5747,
    63698 => -5744,
    63699 => -5741,
    63700 => -5738,
    63701 => -5735,
    63702 => -5732,
    63703 => -5729,
    63704 => -5726,
    63705 => -5723,
    63706 => -5719,
    63707 => -5716,
    63708 => -5713,
    63709 => -5710,
    63710 => -5707,
    63711 => -5704,
    63712 => -5701,
    63713 => -5698,
    63714 => -5695,
    63715 => -5692,
    63716 => -5689,
    63717 => -5685,
    63718 => -5682,
    63719 => -5679,
    63720 => -5676,
    63721 => -5673,
    63722 => -5670,
    63723 => -5667,
    63724 => -5664,
    63725 => -5661,
    63726 => -5658,
    63727 => -5655,
    63728 => -5651,
    63729 => -5648,
    63730 => -5645,
    63731 => -5642,
    63732 => -5639,
    63733 => -5636,
    63734 => -5633,
    63735 => -5630,
    63736 => -5627,
    63737 => -5624,
    63738 => -5620,
    63739 => -5617,
    63740 => -5614,
    63741 => -5611,
    63742 => -5608,
    63743 => -5605,
    63744 => -5602,
    63745 => -5599,
    63746 => -5596,
    63747 => -5593,
    63748 => -5590,
    63749 => -5586,
    63750 => -5583,
    63751 => -5580,
    63752 => -5577,
    63753 => -5574,
    63754 => -5571,
    63755 => -5568,
    63756 => -5565,
    63757 => -5562,
    63758 => -5559,
    63759 => -5555,
    63760 => -5552,
    63761 => -5549,
    63762 => -5546,
    63763 => -5543,
    63764 => -5540,
    63765 => -5537,
    63766 => -5534,
    63767 => -5531,
    63768 => -5528,
    63769 => -5525,
    63770 => -5521,
    63771 => -5518,
    63772 => -5515,
    63773 => -5512,
    63774 => -5509,
    63775 => -5506,
    63776 => -5503,
    63777 => -5500,
    63778 => -5497,
    63779 => -5494,
    63780 => -5490,
    63781 => -5487,
    63782 => -5484,
    63783 => -5481,
    63784 => -5478,
    63785 => -5475,
    63786 => -5472,
    63787 => -5469,
    63788 => -5466,
    63789 => -5463,
    63790 => -5459,
    63791 => -5456,
    63792 => -5453,
    63793 => -5450,
    63794 => -5447,
    63795 => -5444,
    63796 => -5441,
    63797 => -5438,
    63798 => -5435,
    63799 => -5432,
    63800 => -5428,
    63801 => -5425,
    63802 => -5422,
    63803 => -5419,
    63804 => -5416,
    63805 => -5413,
    63806 => -5410,
    63807 => -5407,
    63808 => -5404,
    63809 => -5401,
    63810 => -5398,
    63811 => -5394,
    63812 => -5391,
    63813 => -5388,
    63814 => -5385,
    63815 => -5382,
    63816 => -5379,
    63817 => -5376,
    63818 => -5373,
    63819 => -5370,
    63820 => -5367,
    63821 => -5363,
    63822 => -5360,
    63823 => -5357,
    63824 => -5354,
    63825 => -5351,
    63826 => -5348,
    63827 => -5345,
    63828 => -5342,
    63829 => -5339,
    63830 => -5336,
    63831 => -5332,
    63832 => -5329,
    63833 => -5326,
    63834 => -5323,
    63835 => -5320,
    63836 => -5317,
    63837 => -5314,
    63838 => -5311,
    63839 => -5308,
    63840 => -5305,
    63841 => -5301,
    63842 => -5298,
    63843 => -5295,
    63844 => -5292,
    63845 => -5289,
    63846 => -5286,
    63847 => -5283,
    63848 => -5280,
    63849 => -5277,
    63850 => -5274,
    63851 => -5270,
    63852 => -5267,
    63853 => -5264,
    63854 => -5261,
    63855 => -5258,
    63856 => -5255,
    63857 => -5252,
    63858 => -5249,
    63859 => -5246,
    63860 => -5243,
    63861 => -5239,
    63862 => -5236,
    63863 => -5233,
    63864 => -5230,
    63865 => -5227,
    63866 => -5224,
    63867 => -5221,
    63868 => -5218,
    63869 => -5215,
    63870 => -5212,
    63871 => -5208,
    63872 => -5205,
    63873 => -5202,
    63874 => -5199,
    63875 => -5196,
    63876 => -5193,
    63877 => -5190,
    63878 => -5187,
    63879 => -5184,
    63880 => -5180,
    63881 => -5177,
    63882 => -5174,
    63883 => -5171,
    63884 => -5168,
    63885 => -5165,
    63886 => -5162,
    63887 => -5159,
    63888 => -5156,
    63889 => -5153,
    63890 => -5149,
    63891 => -5146,
    63892 => -5143,
    63893 => -5140,
    63894 => -5137,
    63895 => -5134,
    63896 => -5131,
    63897 => -5128,
    63898 => -5125,
    63899 => -5122,
    63900 => -5118,
    63901 => -5115,
    63902 => -5112,
    63903 => -5109,
    63904 => -5106,
    63905 => -5103,
    63906 => -5100,
    63907 => -5097,
    63908 => -5094,
    63909 => -5091,
    63910 => -5087,
    63911 => -5084,
    63912 => -5081,
    63913 => -5078,
    63914 => -5075,
    63915 => -5072,
    63916 => -5069,
    63917 => -5066,
    63918 => -5063,
    63919 => -5059,
    63920 => -5056,
    63921 => -5053,
    63922 => -5050,
    63923 => -5047,
    63924 => -5044,
    63925 => -5041,
    63926 => -5038,
    63927 => -5035,
    63928 => -5032,
    63929 => -5028,
    63930 => -5025,
    63931 => -5022,
    63932 => -5019,
    63933 => -5016,
    63934 => -5013,
    63935 => -5010,
    63936 => -5007,
    63937 => -5004,
    63938 => -5000,
    63939 => -4997,
    63940 => -4994,
    63941 => -4991,
    63942 => -4988,
    63943 => -4985,
    63944 => -4982,
    63945 => -4979,
    63946 => -4976,
    63947 => -4973,
    63948 => -4969,
    63949 => -4966,
    63950 => -4963,
    63951 => -4960,
    63952 => -4957,
    63953 => -4954,
    63954 => -4951,
    63955 => -4948,
    63956 => -4945,
    63957 => -4941,
    63958 => -4938,
    63959 => -4935,
    63960 => -4932,
    63961 => -4929,
    63962 => -4926,
    63963 => -4923,
    63964 => -4920,
    63965 => -4917,
    63966 => -4914,
    63967 => -4910,
    63968 => -4907,
    63969 => -4904,
    63970 => -4901,
    63971 => -4898,
    63972 => -4895,
    63973 => -4892,
    63974 => -4889,
    63975 => -4886,
    63976 => -4882,
    63977 => -4879,
    63978 => -4876,
    63979 => -4873,
    63980 => -4870,
    63981 => -4867,
    63982 => -4864,
    63983 => -4861,
    63984 => -4858,
    63985 => -4855,
    63986 => -4851,
    63987 => -4848,
    63988 => -4845,
    63989 => -4842,
    63990 => -4839,
    63991 => -4836,
    63992 => -4833,
    63993 => -4830,
    63994 => -4827,
    63995 => -4823,
    63996 => -4820,
    63997 => -4817,
    63998 => -4814,
    63999 => -4811,
    64000 => -4808,
    64001 => -4805,
    64002 => -4802,
    64003 => -4799,
    64004 => -4795,
    64005 => -4792,
    64006 => -4789,
    64007 => -4786,
    64008 => -4783,
    64009 => -4780,
    64010 => -4777,
    64011 => -4774,
    64012 => -4771,
    64013 => -4768,
    64014 => -4764,
    64015 => -4761,
    64016 => -4758,
    64017 => -4755,
    64018 => -4752,
    64019 => -4749,
    64020 => -4746,
    64021 => -4743,
    64022 => -4740,
    64023 => -4736,
    64024 => -4733,
    64025 => -4730,
    64026 => -4727,
    64027 => -4724,
    64028 => -4721,
    64029 => -4718,
    64030 => -4715,
    64031 => -4712,
    64032 => -4708,
    64033 => -4705,
    64034 => -4702,
    64035 => -4699,
    64036 => -4696,
    64037 => -4693,
    64038 => -4690,
    64039 => -4687,
    64040 => -4684,
    64041 => -4680,
    64042 => -4677,
    64043 => -4674,
    64044 => -4671,
    64045 => -4668,
    64046 => -4665,
    64047 => -4662,
    64048 => -4659,
    64049 => -4656,
    64050 => -4652,
    64051 => -4649,
    64052 => -4646,
    64053 => -4643,
    64054 => -4640,
    64055 => -4637,
    64056 => -4634,
    64057 => -4631,
    64058 => -4628,
    64059 => -4624,
    64060 => -4621,
    64061 => -4618,
    64062 => -4615,
    64063 => -4612,
    64064 => -4609,
    64065 => -4606,
    64066 => -4603,
    64067 => -4600,
    64068 => -4597,
    64069 => -4593,
    64070 => -4590,
    64071 => -4587,
    64072 => -4584,
    64073 => -4581,
    64074 => -4578,
    64075 => -4575,
    64076 => -4572,
    64077 => -4569,
    64078 => -4565,
    64079 => -4562,
    64080 => -4559,
    64081 => -4556,
    64082 => -4553,
    64083 => -4550,
    64084 => -4547,
    64085 => -4544,
    64086 => -4541,
    64087 => -4537,
    64088 => -4534,
    64089 => -4531,
    64090 => -4528,
    64091 => -4525,
    64092 => -4522,
    64093 => -4519,
    64094 => -4516,
    64095 => -4513,
    64096 => -4509,
    64097 => -4506,
    64098 => -4503,
    64099 => -4500,
    64100 => -4497,
    64101 => -4494,
    64102 => -4491,
    64103 => -4488,
    64104 => -4485,
    64105 => -4481,
    64106 => -4478,
    64107 => -4475,
    64108 => -4472,
    64109 => -4469,
    64110 => -4466,
    64111 => -4463,
    64112 => -4460,
    64113 => -4456,
    64114 => -4453,
    64115 => -4450,
    64116 => -4447,
    64117 => -4444,
    64118 => -4441,
    64119 => -4438,
    64120 => -4435,
    64121 => -4432,
    64122 => -4428,
    64123 => -4425,
    64124 => -4422,
    64125 => -4419,
    64126 => -4416,
    64127 => -4413,
    64128 => -4410,
    64129 => -4407,
    64130 => -4404,
    64131 => -4400,
    64132 => -4397,
    64133 => -4394,
    64134 => -4391,
    64135 => -4388,
    64136 => -4385,
    64137 => -4382,
    64138 => -4379,
    64139 => -4376,
    64140 => -4372,
    64141 => -4369,
    64142 => -4366,
    64143 => -4363,
    64144 => -4360,
    64145 => -4357,
    64146 => -4354,
    64147 => -4351,
    64148 => -4348,
    64149 => -4344,
    64150 => -4341,
    64151 => -4338,
    64152 => -4335,
    64153 => -4332,
    64154 => -4329,
    64155 => -4326,
    64156 => -4323,
    64157 => -4320,
    64158 => -4316,
    64159 => -4313,
    64160 => -4310,
    64161 => -4307,
    64162 => -4304,
    64163 => -4301,
    64164 => -4298,
    64165 => -4295,
    64166 => -4291,
    64167 => -4288,
    64168 => -4285,
    64169 => -4282,
    64170 => -4279,
    64171 => -4276,
    64172 => -4273,
    64173 => -4270,
    64174 => -4267,
    64175 => -4263,
    64176 => -4260,
    64177 => -4257,
    64178 => -4254,
    64179 => -4251,
    64180 => -4248,
    64181 => -4245,
    64182 => -4242,
    64183 => -4239,
    64184 => -4235,
    64185 => -4232,
    64186 => -4229,
    64187 => -4226,
    64188 => -4223,
    64189 => -4220,
    64190 => -4217,
    64191 => -4214,
    64192 => -4210,
    64193 => -4207,
    64194 => -4204,
    64195 => -4201,
    64196 => -4198,
    64197 => -4195,
    64198 => -4192,
    64199 => -4189,
    64200 => -4186,
    64201 => -4182,
    64202 => -4179,
    64203 => -4176,
    64204 => -4173,
    64205 => -4170,
    64206 => -4167,
    64207 => -4164,
    64208 => -4161,
    64209 => -4158,
    64210 => -4154,
    64211 => -4151,
    64212 => -4148,
    64213 => -4145,
    64214 => -4142,
    64215 => -4139,
    64216 => -4136,
    64217 => -4133,
    64218 => -4129,
    64219 => -4126,
    64220 => -4123,
    64221 => -4120,
    64222 => -4117,
    64223 => -4114,
    64224 => -4111,
    64225 => -4108,
    64226 => -4105,
    64227 => -4101,
    64228 => -4098,
    64229 => -4095,
    64230 => -4092,
    64231 => -4089,
    64232 => -4086,
    64233 => -4083,
    64234 => -4080,
    64235 => -4076,
    64236 => -4073,
    64237 => -4070,
    64238 => -4067,
    64239 => -4064,
    64240 => -4061,
    64241 => -4058,
    64242 => -4055,
    64243 => -4052,
    64244 => -4048,
    64245 => -4045,
    64246 => -4042,
    64247 => -4039,
    64248 => -4036,
    64249 => -4033,
    64250 => -4030,
    64251 => -4027,
    64252 => -4024,
    64253 => -4020,
    64254 => -4017,
    64255 => -4014,
    64256 => -4011,
    64257 => -4008,
    64258 => -4005,
    64259 => -4002,
    64260 => -3999,
    64261 => -3995,
    64262 => -3992,
    64263 => -3989,
    64264 => -3986,
    64265 => -3983,
    64266 => -3980,
    64267 => -3977,
    64268 => -3974,
    64269 => -3970,
    64270 => -3967,
    64271 => -3964,
    64272 => -3961,
    64273 => -3958,
    64274 => -3955,
    64275 => -3952,
    64276 => -3949,
    64277 => -3946,
    64278 => -3942,
    64279 => -3939,
    64280 => -3936,
    64281 => -3933,
    64282 => -3930,
    64283 => -3927,
    64284 => -3924,
    64285 => -3921,
    64286 => -3917,
    64287 => -3914,
    64288 => -3911,
    64289 => -3908,
    64290 => -3905,
    64291 => -3902,
    64292 => -3899,
    64293 => -3896,
    64294 => -3893,
    64295 => -3889,
    64296 => -3886,
    64297 => -3883,
    64298 => -3880,
    64299 => -3877,
    64300 => -3874,
    64301 => -3871,
    64302 => -3868,
    64303 => -3864,
    64304 => -3861,
    64305 => -3858,
    64306 => -3855,
    64307 => -3852,
    64308 => -3849,
    64309 => -3846,
    64310 => -3843,
    64311 => -3839,
    64312 => -3836,
    64313 => -3833,
    64314 => -3830,
    64315 => -3827,
    64316 => -3824,
    64317 => -3821,
    64318 => -3818,
    64319 => -3815,
    64320 => -3811,
    64321 => -3808,
    64322 => -3805,
    64323 => -3802,
    64324 => -3799,
    64325 => -3796,
    64326 => -3793,
    64327 => -3790,
    64328 => -3786,
    64329 => -3783,
    64330 => -3780,
    64331 => -3777,
    64332 => -3774,
    64333 => -3771,
    64334 => -3768,
    64335 => -3765,
    64336 => -3761,
    64337 => -3758,
    64338 => -3755,
    64339 => -3752,
    64340 => -3749,
    64341 => -3746,
    64342 => -3743,
    64343 => -3740,
    64344 => -3737,
    64345 => -3733,
    64346 => -3730,
    64347 => -3727,
    64348 => -3724,
    64349 => -3721,
    64350 => -3718,
    64351 => -3715,
    64352 => -3712,
    64353 => -3708,
    64354 => -3705,
    64355 => -3702,
    64356 => -3699,
    64357 => -3696,
    64358 => -3693,
    64359 => -3690,
    64360 => -3687,
    64361 => -3683,
    64362 => -3680,
    64363 => -3677,
    64364 => -3674,
    64365 => -3671,
    64366 => -3668,
    64367 => -3665,
    64368 => -3662,
    64369 => -3658,
    64370 => -3655,
    64371 => -3652,
    64372 => -3649,
    64373 => -3646,
    64374 => -3643,
    64375 => -3640,
    64376 => -3637,
    64377 => -3634,
    64378 => -3630,
    64379 => -3627,
    64380 => -3624,
    64381 => -3621,
    64382 => -3618,
    64383 => -3615,
    64384 => -3612,
    64385 => -3609,
    64386 => -3605,
    64387 => -3602,
    64388 => -3599,
    64389 => -3596,
    64390 => -3593,
    64391 => -3590,
    64392 => -3587,
    64393 => -3584,
    64394 => -3580,
    64395 => -3577,
    64396 => -3574,
    64397 => -3571,
    64398 => -3568,
    64399 => -3565,
    64400 => -3562,
    64401 => -3559,
    64402 => -3555,
    64403 => -3552,
    64404 => -3549,
    64405 => -3546,
    64406 => -3543,
    64407 => -3540,
    64408 => -3537,
    64409 => -3534,
    64410 => -3530,
    64411 => -3527,
    64412 => -3524,
    64413 => -3521,
    64414 => -3518,
    64415 => -3515,
    64416 => -3512,
    64417 => -3509,
    64418 => -3505,
    64419 => -3502,
    64420 => -3499,
    64421 => -3496,
    64422 => -3493,
    64423 => -3490,
    64424 => -3487,
    64425 => -3484,
    64426 => -3480,
    64427 => -3477,
    64428 => -3474,
    64429 => -3471,
    64430 => -3468,
    64431 => -3465,
    64432 => -3462,
    64433 => -3459,
    64434 => -3455,
    64435 => -3452,
    64436 => -3449,
    64437 => -3446,
    64438 => -3443,
    64439 => -3440,
    64440 => -3437,
    64441 => -3434,
    64442 => -3430,
    64443 => -3427,
    64444 => -3424,
    64445 => -3421,
    64446 => -3418,
    64447 => -3415,
    64448 => -3412,
    64449 => -3409,
    64450 => -3406,
    64451 => -3402,
    64452 => -3399,
    64453 => -3396,
    64454 => -3393,
    64455 => -3390,
    64456 => -3387,
    64457 => -3384,
    64458 => -3381,
    64459 => -3377,
    64460 => -3374,
    64461 => -3371,
    64462 => -3368,
    64463 => -3365,
    64464 => -3362,
    64465 => -3359,
    64466 => -3356,
    64467 => -3352,
    64468 => -3349,
    64469 => -3346,
    64470 => -3343,
    64471 => -3340,
    64472 => -3337,
    64473 => -3334,
    64474 => -3331,
    64475 => -3327,
    64476 => -3324,
    64477 => -3321,
    64478 => -3318,
    64479 => -3315,
    64480 => -3312,
    64481 => -3309,
    64482 => -3306,
    64483 => -3302,
    64484 => -3299,
    64485 => -3296,
    64486 => -3293,
    64487 => -3290,
    64488 => -3287,
    64489 => -3284,
    64490 => -3281,
    64491 => -3277,
    64492 => -3274,
    64493 => -3271,
    64494 => -3268,
    64495 => -3265,
    64496 => -3262,
    64497 => -3259,
    64498 => -3255,
    64499 => -3252,
    64500 => -3249,
    64501 => -3246,
    64502 => -3243,
    64503 => -3240,
    64504 => -3237,
    64505 => -3234,
    64506 => -3230,
    64507 => -3227,
    64508 => -3224,
    64509 => -3221,
    64510 => -3218,
    64511 => -3215,
    64512 => -3212,
    64513 => -3209,
    64514 => -3205,
    64515 => -3202,
    64516 => -3199,
    64517 => -3196,
    64518 => -3193,
    64519 => -3190,
    64520 => -3187,
    64521 => -3184,
    64522 => -3180,
    64523 => -3177,
    64524 => -3174,
    64525 => -3171,
    64526 => -3168,
    64527 => -3165,
    64528 => -3162,
    64529 => -3159,
    64530 => -3155,
    64531 => -3152,
    64532 => -3149,
    64533 => -3146,
    64534 => -3143,
    64535 => -3140,
    64536 => -3137,
    64537 => -3134,
    64538 => -3130,
    64539 => -3127,
    64540 => -3124,
    64541 => -3121,
    64542 => -3118,
    64543 => -3115,
    64544 => -3112,
    64545 => -3109,
    64546 => -3105,
    64547 => -3102,
    64548 => -3099,
    64549 => -3096,
    64550 => -3093,
    64551 => -3090,
    64552 => -3087,
    64553 => -3084,
    64554 => -3080,
    64555 => -3077,
    64556 => -3074,
    64557 => -3071,
    64558 => -3068,
    64559 => -3065,
    64560 => -3062,
    64561 => -3059,
    64562 => -3055,
    64563 => -3052,
    64564 => -3049,
    64565 => -3046,
    64566 => -3043,
    64567 => -3040,
    64568 => -3037,
    64569 => -3033,
    64570 => -3030,
    64571 => -3027,
    64572 => -3024,
    64573 => -3021,
    64574 => -3018,
    64575 => -3015,
    64576 => -3012,
    64577 => -3008,
    64578 => -3005,
    64579 => -3002,
    64580 => -2999,
    64581 => -2996,
    64582 => -2993,
    64583 => -2990,
    64584 => -2987,
    64585 => -2983,
    64586 => -2980,
    64587 => -2977,
    64588 => -2974,
    64589 => -2971,
    64590 => -2968,
    64591 => -2965,
    64592 => -2962,
    64593 => -2958,
    64594 => -2955,
    64595 => -2952,
    64596 => -2949,
    64597 => -2946,
    64598 => -2943,
    64599 => -2940,
    64600 => -2936,
    64601 => -2933,
    64602 => -2930,
    64603 => -2927,
    64604 => -2924,
    64605 => -2921,
    64606 => -2918,
    64607 => -2915,
    64608 => -2911,
    64609 => -2908,
    64610 => -2905,
    64611 => -2902,
    64612 => -2899,
    64613 => -2896,
    64614 => -2893,
    64615 => -2890,
    64616 => -2886,
    64617 => -2883,
    64618 => -2880,
    64619 => -2877,
    64620 => -2874,
    64621 => -2871,
    64622 => -2868,
    64623 => -2865,
    64624 => -2861,
    64625 => -2858,
    64626 => -2855,
    64627 => -2852,
    64628 => -2849,
    64629 => -2846,
    64630 => -2843,
    64631 => -2839,
    64632 => -2836,
    64633 => -2833,
    64634 => -2830,
    64635 => -2827,
    64636 => -2824,
    64637 => -2821,
    64638 => -2818,
    64639 => -2814,
    64640 => -2811,
    64641 => -2808,
    64642 => -2805,
    64643 => -2802,
    64644 => -2799,
    64645 => -2796,
    64646 => -2793,
    64647 => -2789,
    64648 => -2786,
    64649 => -2783,
    64650 => -2780,
    64651 => -2777,
    64652 => -2774,
    64653 => -2771,
    64654 => -2767,
    64655 => -2764,
    64656 => -2761,
    64657 => -2758,
    64658 => -2755,
    64659 => -2752,
    64660 => -2749,
    64661 => -2746,
    64662 => -2742,
    64663 => -2739,
    64664 => -2736,
    64665 => -2733,
    64666 => -2730,
    64667 => -2727,
    64668 => -2724,
    64669 => -2721,
    64670 => -2717,
    64671 => -2714,
    64672 => -2711,
    64673 => -2708,
    64674 => -2705,
    64675 => -2702,
    64676 => -2699,
    64677 => -2695,
    64678 => -2692,
    64679 => -2689,
    64680 => -2686,
    64681 => -2683,
    64682 => -2680,
    64683 => -2677,
    64684 => -2674,
    64685 => -2670,
    64686 => -2667,
    64687 => -2664,
    64688 => -2661,
    64689 => -2658,
    64690 => -2655,
    64691 => -2652,
    64692 => -2649,
    64693 => -2645,
    64694 => -2642,
    64695 => -2639,
    64696 => -2636,
    64697 => -2633,
    64698 => -2630,
    64699 => -2627,
    64700 => -2623,
    64701 => -2620,
    64702 => -2617,
    64703 => -2614,
    64704 => -2611,
    64705 => -2608,
    64706 => -2605,
    64707 => -2602,
    64708 => -2598,
    64709 => -2595,
    64710 => -2592,
    64711 => -2589,
    64712 => -2586,
    64713 => -2583,
    64714 => -2580,
    64715 => -2577,
    64716 => -2573,
    64717 => -2570,
    64718 => -2567,
    64719 => -2564,
    64720 => -2561,
    64721 => -2558,
    64722 => -2555,
    64723 => -2551,
    64724 => -2548,
    64725 => -2545,
    64726 => -2542,
    64727 => -2539,
    64728 => -2536,
    64729 => -2533,
    64730 => -2530,
    64731 => -2526,
    64732 => -2523,
    64733 => -2520,
    64734 => -2517,
    64735 => -2514,
    64736 => -2511,
    64737 => -2508,
    64738 => -2504,
    64739 => -2501,
    64740 => -2498,
    64741 => -2495,
    64742 => -2492,
    64743 => -2489,
    64744 => -2486,
    64745 => -2483,
    64746 => -2479,
    64747 => -2476,
    64748 => -2473,
    64749 => -2470,
    64750 => -2467,
    64751 => -2464,
    64752 => -2461,
    64753 => -2457,
    64754 => -2454,
    64755 => -2451,
    64756 => -2448,
    64757 => -2445,
    64758 => -2442,
    64759 => -2439,
    64760 => -2436,
    64761 => -2432,
    64762 => -2429,
    64763 => -2426,
    64764 => -2423,
    64765 => -2420,
    64766 => -2417,
    64767 => -2414,
    64768 => -2410,
    64769 => -2407,
    64770 => -2404,
    64771 => -2401,
    64772 => -2398,
    64773 => -2395,
    64774 => -2392,
    64775 => -2389,
    64776 => -2385,
    64777 => -2382,
    64778 => -2379,
    64779 => -2376,
    64780 => -2373,
    64781 => -2370,
    64782 => -2367,
    64783 => -2363,
    64784 => -2360,
    64785 => -2357,
    64786 => -2354,
    64787 => -2351,
    64788 => -2348,
    64789 => -2345,
    64790 => -2342,
    64791 => -2338,
    64792 => -2335,
    64793 => -2332,
    64794 => -2329,
    64795 => -2326,
    64796 => -2323,
    64797 => -2320,
    64798 => -2316,
    64799 => -2313,
    64800 => -2310,
    64801 => -2307,
    64802 => -2304,
    64803 => -2301,
    64804 => -2298,
    64805 => -2295,
    64806 => -2291,
    64807 => -2288,
    64808 => -2285,
    64809 => -2282,
    64810 => -2279,
    64811 => -2276,
    64812 => -2273,
    64813 => -2269,
    64814 => -2266,
    64815 => -2263,
    64816 => -2260,
    64817 => -2257,
    64818 => -2254,
    64819 => -2251,
    64820 => -2248,
    64821 => -2244,
    64822 => -2241,
    64823 => -2238,
    64824 => -2235,
    64825 => -2232,
    64826 => -2229,
    64827 => -2226,
    64828 => -2222,
    64829 => -2219,
    64830 => -2216,
    64831 => -2213,
    64832 => -2210,
    64833 => -2207,
    64834 => -2204,
    64835 => -2201,
    64836 => -2197,
    64837 => -2194,
    64838 => -2191,
    64839 => -2188,
    64840 => -2185,
    64841 => -2182,
    64842 => -2179,
    64843 => -2175,
    64844 => -2172,
    64845 => -2169,
    64846 => -2166,
    64847 => -2163,
    64848 => -2160,
    64849 => -2157,
    64850 => -2154,
    64851 => -2150,
    64852 => -2147,
    64853 => -2144,
    64854 => -2141,
    64855 => -2138,
    64856 => -2135,
    64857 => -2132,
    64858 => -2128,
    64859 => -2125,
    64860 => -2122,
    64861 => -2119,
    64862 => -2116,
    64863 => -2113,
    64864 => -2110,
    64865 => -2106,
    64866 => -2103,
    64867 => -2100,
    64868 => -2097,
    64869 => -2094,
    64870 => -2091,
    64871 => -2088,
    64872 => -2085,
    64873 => -2081,
    64874 => -2078,
    64875 => -2075,
    64876 => -2072,
    64877 => -2069,
    64878 => -2066,
    64879 => -2063,
    64880 => -2059,
    64881 => -2056,
    64882 => -2053,
    64883 => -2050,
    64884 => -2047,
    64885 => -2044,
    64886 => -2041,
    64887 => -2038,
    64888 => -2034,
    64889 => -2031,
    64890 => -2028,
    64891 => -2025,
    64892 => -2022,
    64893 => -2019,
    64894 => -2016,
    64895 => -2012,
    64896 => -2009,
    64897 => -2006,
    64898 => -2003,
    64899 => -2000,
    64900 => -1997,
    64901 => -1994,
    64902 => -1990,
    64903 => -1987,
    64904 => -1984,
    64905 => -1981,
    64906 => -1978,
    64907 => -1975,
    64908 => -1972,
    64909 => -1969,
    64910 => -1965,
    64911 => -1962,
    64912 => -1959,
    64913 => -1956,
    64914 => -1953,
    64915 => -1950,
    64916 => -1947,
    64917 => -1943,
    64918 => -1940,
    64919 => -1937,
    64920 => -1934,
    64921 => -1931,
    64922 => -1928,
    64923 => -1925,
    64924 => -1921,
    64925 => -1918,
    64926 => -1915,
    64927 => -1912,
    64928 => -1909,
    64929 => -1906,
    64930 => -1903,
    64931 => -1900,
    64932 => -1896,
    64933 => -1893,
    64934 => -1890,
    64935 => -1887,
    64936 => -1884,
    64937 => -1881,
    64938 => -1878,
    64939 => -1874,
    64940 => -1871,
    64941 => -1868,
    64942 => -1865,
    64943 => -1862,
    64944 => -1859,
    64945 => -1856,
    64946 => -1852,
    64947 => -1849,
    64948 => -1846,
    64949 => -1843,
    64950 => -1840,
    64951 => -1837,
    64952 => -1834,
    64953 => -1831,
    64954 => -1827,
    64955 => -1824,
    64956 => -1821,
    64957 => -1818,
    64958 => -1815,
    64959 => -1812,
    64960 => -1809,
    64961 => -1805,
    64962 => -1802,
    64963 => -1799,
    64964 => -1796,
    64965 => -1793,
    64966 => -1790,
    64967 => -1787,
    64968 => -1783,
    64969 => -1780,
    64970 => -1777,
    64971 => -1774,
    64972 => -1771,
    64973 => -1768,
    64974 => -1765,
    64975 => -1762,
    64976 => -1758,
    64977 => -1755,
    64978 => -1752,
    64979 => -1749,
    64980 => -1746,
    64981 => -1743,
    64982 => -1740,
    64983 => -1736,
    64984 => -1733,
    64985 => -1730,
    64986 => -1727,
    64987 => -1724,
    64988 => -1721,
    64989 => -1718,
    64990 => -1714,
    64991 => -1711,
    64992 => -1708,
    64993 => -1705,
    64994 => -1702,
    64995 => -1699,
    64996 => -1696,
    64997 => -1693,
    64998 => -1689,
    64999 => -1686,
    65000 => -1683,
    65001 => -1680,
    65002 => -1677,
    65003 => -1674,
    65004 => -1671,
    65005 => -1667,
    65006 => -1664,
    65007 => -1661,
    65008 => -1658,
    65009 => -1655,
    65010 => -1652,
    65011 => -1649,
    65012 => -1645,
    65013 => -1642,
    65014 => -1639,
    65015 => -1636,
    65016 => -1633,
    65017 => -1630,
    65018 => -1627,
    65019 => -1623,
    65020 => -1620,
    65021 => -1617,
    65022 => -1614,
    65023 => -1611,
    65024 => -1608,
    65025 => -1605,
    65026 => -1602,
    65027 => -1598,
    65028 => -1595,
    65029 => -1592,
    65030 => -1589,
    65031 => -1586,
    65032 => -1583,
    65033 => -1580,
    65034 => -1576,
    65035 => -1573,
    65036 => -1570,
    65037 => -1567,
    65038 => -1564,
    65039 => -1561,
    65040 => -1558,
    65041 => -1554,
    65042 => -1551,
    65043 => -1548,
    65044 => -1545,
    65045 => -1542,
    65046 => -1539,
    65047 => -1536,
    65048 => -1532,
    65049 => -1529,
    65050 => -1526,
    65051 => -1523,
    65052 => -1520,
    65053 => -1517,
    65054 => -1514,
    65055 => -1511,
    65056 => -1507,
    65057 => -1504,
    65058 => -1501,
    65059 => -1498,
    65060 => -1495,
    65061 => -1492,
    65062 => -1489,
    65063 => -1485,
    65064 => -1482,
    65065 => -1479,
    65066 => -1476,
    65067 => -1473,
    65068 => -1470,
    65069 => -1467,
    65070 => -1463,
    65071 => -1460,
    65072 => -1457,
    65073 => -1454,
    65074 => -1451,
    65075 => -1448,
    65076 => -1445,
    65077 => -1441,
    65078 => -1438,
    65079 => -1435,
    65080 => -1432,
    65081 => -1429,
    65082 => -1426,
    65083 => -1423,
    65084 => -1420,
    65085 => -1416,
    65086 => -1413,
    65087 => -1410,
    65088 => -1407,
    65089 => -1404,
    65090 => -1401,
    65091 => -1398,
    65092 => -1394,
    65093 => -1391,
    65094 => -1388,
    65095 => -1385,
    65096 => -1382,
    65097 => -1379,
    65098 => -1376,
    65099 => -1372,
    65100 => -1369,
    65101 => -1366,
    65102 => -1363,
    65103 => -1360,
    65104 => -1357,
    65105 => -1354,
    65106 => -1350,
    65107 => -1347,
    65108 => -1344,
    65109 => -1341,
    65110 => -1338,
    65111 => -1335,
    65112 => -1332,
    65113 => -1328,
    65114 => -1325,
    65115 => -1322,
    65116 => -1319,
    65117 => -1316,
    65118 => -1313,
    65119 => -1310,
    65120 => -1307,
    65121 => -1303,
    65122 => -1300,
    65123 => -1297,
    65124 => -1294,
    65125 => -1291,
    65126 => -1288,
    65127 => -1285,
    65128 => -1281,
    65129 => -1278,
    65130 => -1275,
    65131 => -1272,
    65132 => -1269,
    65133 => -1266,
    65134 => -1263,
    65135 => -1259,
    65136 => -1256,
    65137 => -1253,
    65138 => -1250,
    65139 => -1247,
    65140 => -1244,
    65141 => -1241,
    65142 => -1237,
    65143 => -1234,
    65144 => -1231,
    65145 => -1228,
    65146 => -1225,
    65147 => -1222,
    65148 => -1219,
    65149 => -1215,
    65150 => -1212,
    65151 => -1209,
    65152 => -1206,
    65153 => -1203,
    65154 => -1200,
    65155 => -1197,
    65156 => -1194,
    65157 => -1190,
    65158 => -1187,
    65159 => -1184,
    65160 => -1181,
    65161 => -1178,
    65162 => -1175,
    65163 => -1172,
    65164 => -1168,
    65165 => -1165,
    65166 => -1162,
    65167 => -1159,
    65168 => -1156,
    65169 => -1153,
    65170 => -1150,
    65171 => -1146,
    65172 => -1143,
    65173 => -1140,
    65174 => -1137,
    65175 => -1134,
    65176 => -1131,
    65177 => -1128,
    65178 => -1124,
    65179 => -1121,
    65180 => -1118,
    65181 => -1115,
    65182 => -1112,
    65183 => -1109,
    65184 => -1106,
    65185 => -1102,
    65186 => -1099,
    65187 => -1096,
    65188 => -1093,
    65189 => -1090,
    65190 => -1087,
    65191 => -1084,
    65192 => -1080,
    65193 => -1077,
    65194 => -1074,
    65195 => -1071,
    65196 => -1068,
    65197 => -1065,
    65198 => -1062,
    65199 => -1059,
    65200 => -1055,
    65201 => -1052,
    65202 => -1049,
    65203 => -1046,
    65204 => -1043,
    65205 => -1040,
    65206 => -1037,
    65207 => -1033,
    65208 => -1030,
    65209 => -1027,
    65210 => -1024,
    65211 => -1021,
    65212 => -1018,
    65213 => -1015,
    65214 => -1011,
    65215 => -1008,
    65216 => -1005,
    65217 => -1002,
    65218 => -999,
    65219 => -996,
    65220 => -993,
    65221 => -989,
    65222 => -986,
    65223 => -983,
    65224 => -980,
    65225 => -977,
    65226 => -974,
    65227 => -971,
    65228 => -967,
    65229 => -964,
    65230 => -961,
    65231 => -958,
    65232 => -955,
    65233 => -952,
    65234 => -949,
    65235 => -945,
    65236 => -942,
    65237 => -939,
    65238 => -936,
    65239 => -933,
    65240 => -930,
    65241 => -927,
    65242 => -923,
    65243 => -920,
    65244 => -917,
    65245 => -914,
    65246 => -911,
    65247 => -908,
    65248 => -905,
    65249 => -901,
    65250 => -898,
    65251 => -895,
    65252 => -892,
    65253 => -889,
    65254 => -886,
    65255 => -883,
    65256 => -880,
    65257 => -876,
    65258 => -873,
    65259 => -870,
    65260 => -867,
    65261 => -864,
    65262 => -861,
    65263 => -858,
    65264 => -854,
    65265 => -851,
    65266 => -848,
    65267 => -845,
    65268 => -842,
    65269 => -839,
    65270 => -836,
    65271 => -832,
    65272 => -829,
    65273 => -826,
    65274 => -823,
    65275 => -820,
    65276 => -817,
    65277 => -814,
    65278 => -810,
    65279 => -807,
    65280 => -804,
    65281 => -801,
    65282 => -798,
    65283 => -795,
    65284 => -792,
    65285 => -788,
    65286 => -785,
    65287 => -782,
    65288 => -779,
    65289 => -776,
    65290 => -773,
    65291 => -770,
    65292 => -766,
    65293 => -763,
    65294 => -760,
    65295 => -757,
    65296 => -754,
    65297 => -751,
    65298 => -748,
    65299 => -744,
    65300 => -741,
    65301 => -738,
    65302 => -735,
    65303 => -732,
    65304 => -729,
    65305 => -726,
    65306 => -722,
    65307 => -719,
    65308 => -716,
    65309 => -713,
    65310 => -710,
    65311 => -707,
    65312 => -704,
    65313 => -701,
    65314 => -697,
    65315 => -694,
    65316 => -691,
    65317 => -688,
    65318 => -685,
    65319 => -682,
    65320 => -679,
    65321 => -675,
    65322 => -672,
    65323 => -669,
    65324 => -666,
    65325 => -663,
    65326 => -660,
    65327 => -657,
    65328 => -653,
    65329 => -650,
    65330 => -647,
    65331 => -644,
    65332 => -641,
    65333 => -638,
    65334 => -635,
    65335 => -631,
    65336 => -628,
    65337 => -625,
    65338 => -622,
    65339 => -619,
    65340 => -616,
    65341 => -613,
    65342 => -609,
    65343 => -606,
    65344 => -603,
    65345 => -600,
    65346 => -597,
    65347 => -594,
    65348 => -591,
    65349 => -587,
    65350 => -584,
    65351 => -581,
    65352 => -578,
    65353 => -575,
    65354 => -572,
    65355 => -569,
    65356 => -565,
    65357 => -562,
    65358 => -559,
    65359 => -556,
    65360 => -553,
    65361 => -550,
    65362 => -547,
    65363 => -543,
    65364 => -540,
    65365 => -537,
    65366 => -534,
    65367 => -531,
    65368 => -528,
    65369 => -525,
    65370 => -521,
    65371 => -518,
    65372 => -515,
    65373 => -512,
    65374 => -509,
    65375 => -506,
    65376 => -503,
    65377 => -499,
    65378 => -496,
    65379 => -493,
    65380 => -490,
    65381 => -487,
    65382 => -484,
    65383 => -481,
    65384 => -477,
    65385 => -474,
    65386 => -471,
    65387 => -468,
    65388 => -465,
    65389 => -462,
    65390 => -459,
    65391 => -456,
    65392 => -452,
    65393 => -449,
    65394 => -446,
    65395 => -443,
    65396 => -440,
    65397 => -437,
    65398 => -434,
    65399 => -430,
    65400 => -427,
    65401 => -424,
    65402 => -421,
    65403 => -418,
    65404 => -415,
    65405 => -412,
    65406 => -408,
    65407 => -405,
    65408 => -402,
    65409 => -399,
    65410 => -396,
    65411 => -393,
    65412 => -390,
    65413 => -386,
    65414 => -383,
    65415 => -380,
    65416 => -377,
    65417 => -374,
    65418 => -371,
    65419 => -368,
    65420 => -364,
    65421 => -361,
    65422 => -358,
    65423 => -355,
    65424 => -352,
    65425 => -349,
    65426 => -346,
    65427 => -342,
    65428 => -339,
    65429 => -336,
    65430 => -333,
    65431 => -330,
    65432 => -327,
    65433 => -324,
    65434 => -320,
    65435 => -317,
    65436 => -314,
    65437 => -311,
    65438 => -308,
    65439 => -305,
    65440 => -302,
    65441 => -298,
    65442 => -295,
    65443 => -292,
    65444 => -289,
    65445 => -286,
    65446 => -283,
    65447 => -280,
    65448 => -276,
    65449 => -273,
    65450 => -270,
    65451 => -267,
    65452 => -264,
    65453 => -261,
    65454 => -258,
    65455 => -254,
    65456 => -251,
    65457 => -248,
    65458 => -245,
    65459 => -242,
    65460 => -239,
    65461 => -236,
    65462 => -232,
    65463 => -229,
    65464 => -226,
    65465 => -223,
    65466 => -220,
    65467 => -217,
    65468 => -214,
    65469 => -210,
    65470 => -207,
    65471 => -204,
    65472 => -201,
    65473 => -198,
    65474 => -195,
    65475 => -192,
    65476 => -188,
    65477 => -185,
    65478 => -182,
    65479 => -179,
    65480 => -176,
    65481 => -173,
    65482 => -170,
    65483 => -166,
    65484 => -163,
    65485 => -160,
    65486 => -157,
    65487 => -154,
    65488 => -151,
    65489 => -148,
    65490 => -145,
    65491 => -141,
    65492 => -138,
    65493 => -135,
    65494 => -132,
    65495 => -129,
    65496 => -126,
    65497 => -123,
    65498 => -119,
    65499 => -116,
    65500 => -113,
    65501 => -110,
    65502 => -107,
    65503 => -104,
    65504 => -101,
    65505 => -97,
    65506 => -94,
    65507 => -91,
    65508 => -88,
    65509 => -85,
    65510 => -82,
    65511 => -79,
    65512 => -75,
    65513 => -72,
    65514 => -69,
    65515 => -66,
    65516 => -63,
    65517 => -60,
    65518 => -57,
    65519 => -53,
    65520 => -50,
    65521 => -47,
    65522 => -44,
    65523 => -41,
    65524 => -38,
    65525 => -35,
    65526 => -31,
    65527 => -28,
    65528 => -25,
    65529 => -22,
    65530 => -19,
    65531 => -16,
    65532 => -13,
    65533 => -9,
    65534 => -6,
    65535 => -3
  );

begin
  ddfs_out <= std_logic_vector(to_signed(LUT(to_integer(unsigned(address))),16));
end architecture;
