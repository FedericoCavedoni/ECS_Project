library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity qlut_table_16384_7bit is
  generic (
    N : integer := 14;   -- Address width (log2 of 16384)
    P : integer := 7     -- Output width
  );
  port (
    address  : in  std_logic_vector(N-1 downto 0);  -- Address input
    lut_out  : out std_logic_vector(P-1 downto 0)   -- Output data
  );
end entity;

architecture rtl of qlut_table_16384_7bit is
  -- Type declaration for LUT
  type LUT_t is array (natural range 0 to 16383) of integer;
  -- LUT initialization with data
  constant LUT: LUT_t := (
    0 => 0,
    1 => 0,
    2 => 0,
    3 => 0,
    4 => 0,
    5 => 0,
    6 => 0,
    7 => 0,
    8 => 0,
    9 => 0,
    10 => 0,
    11 => 0,
    12 => 0,
    13 => 0,
    14 => 0,
    15 => 0,
    16 => 0,
    17 => 0,
    18 => 0,
    19 => 0,
    20 => 0,
    21 => 0,
    22 => 0,
    23 => 0,
    24 => 0,
    25 => 0,
    26 => 0,
    27 => 0,
    28 => 0,
    29 => 0,
    30 => 0,
    31 => 0,
    32 => 0,
    33 => 0,
    34 => 0,
    35 => 0,
    36 => 0,
    37 => 0,
    38 => 0,
    39 => 0,
    40 => 0,
    41 => 0,
    42 => 0,
    43 => 0,
    44 => 0,
    45 => 0,
    46 => 0,
    47 => 0,
    48 => 0,
    49 => 0,
    50 => 0,
    51 => 0,
    52 => 0,
    53 => 0,
    54 => 0,
    55 => 0,
    56 => 0,
    57 => 0,
    58 => 0,
    59 => 0,
    60 => 0,
    61 => 0,
    62 => 0,
    63 => 0,
    64 => 0,
    65 => 0,
    66 => 0,
    67 => 0,
    68 => 0,
    69 => 0,
    70 => 0,
    71 => 0,
    72 => 0,
    73 => 0,
    74 => 0,
    75 => 0,
    76 => 0,
    77 => 0,
    78 => 0,
    79 => 0,
    80 => 0,
    81 => 0,
    82 => 0,
    83 => 1,
    84 => 1,
    85 => 1,
    86 => 1,
    87 => 1,
    88 => 1,
    89 => 1,
    90 => 1,
    91 => 1,
    92 => 1,
    93 => 1,
    94 => 1,
    95 => 1,
    96 => 1,
    97 => 1,
    98 => 1,
    99 => 1,
    100 => 1,
    101 => 1,
    102 => 1,
    103 => 1,
    104 => 1,
    105 => 1,
    106 => 1,
    107 => 1,
    108 => 1,
    109 => 1,
    110 => 1,
    111 => 1,
    112 => 1,
    113 => 1,
    114 => 1,
    115 => 1,
    116 => 1,
    117 => 1,
    118 => 1,
    119 => 1,
    120 => 1,
    121 => 1,
    122 => 1,
    123 => 1,
    124 => 1,
    125 => 1,
    126 => 1,
    127 => 1,
    128 => 1,
    129 => 1,
    130 => 1,
    131 => 1,
    132 => 1,
    133 => 1,
    134 => 1,
    135 => 1,
    136 => 1,
    137 => 1,
    138 => 1,
    139 => 1,
    140 => 1,
    141 => 1,
    142 => 1,
    143 => 1,
    144 => 1,
    145 => 1,
    146 => 1,
    147 => 1,
    148 => 1,
    149 => 1,
    150 => 1,
    151 => 1,
    152 => 1,
    153 => 1,
    154 => 1,
    155 => 1,
    156 => 1,
    157 => 1,
    158 => 1,
    159 => 1,
    160 => 1,
    161 => 1,
    162 => 1,
    163 => 1,
    164 => 1,
    165 => 1,
    166 => 1,
    167 => 1,
    168 => 1,
    169 => 1,
    170 => 1,
    171 => 1,
    172 => 1,
    173 => 1,
    174 => 1,
    175 => 1,
    176 => 1,
    177 => 1,
    178 => 1,
    179 => 1,
    180 => 1,
    181 => 1,
    182 => 1,
    183 => 1,
    184 => 1,
    185 => 1,
    186 => 1,
    187 => 1,
    188 => 1,
    189 => 1,
    190 => 1,
    191 => 1,
    192 => 1,
    193 => 1,
    194 => 1,
    195 => 1,
    196 => 1,
    197 => 1,
    198 => 1,
    199 => 1,
    200 => 1,
    201 => 1,
    202 => 1,
    203 => 1,
    204 => 1,
    205 => 1,
    206 => 1,
    207 => 1,
    208 => 1,
    209 => 1,
    210 => 1,
    211 => 1,
    212 => 1,
    213 => 1,
    214 => 1,
    215 => 1,
    216 => 1,
    217 => 1,
    218 => 1,
    219 => 1,
    220 => 1,
    221 => 1,
    222 => 1,
    223 => 1,
    224 => 1,
    225 => 1,
    226 => 1,
    227 => 1,
    228 => 1,
    229 => 1,
    230 => 1,
    231 => 1,
    232 => 1,
    233 => 1,
    234 => 1,
    235 => 1,
    236 => 1,
    237 => 1,
    238 => 1,
    239 => 1,
    240 => 1,
    241 => 1,
    242 => 1,
    243 => 1,
    244 => 1,
    245 => 1,
    246 => 1,
    247 => 1,
    248 => 1,
    249 => 2,
    250 => 2,
    251 => 2,
    252 => 2,
    253 => 2,
    254 => 2,
    255 => 2,
    256 => 2,
    257 => 2,
    258 => 2,
    259 => 2,
    260 => 2,
    261 => 2,
    262 => 2,
    263 => 2,
    264 => 2,
    265 => 2,
    266 => 2,
    267 => 2,
    268 => 2,
    269 => 2,
    270 => 2,
    271 => 2,
    272 => 2,
    273 => 2,
    274 => 2,
    275 => 2,
    276 => 2,
    277 => 2,
    278 => 2,
    279 => 2,
    280 => 2,
    281 => 2,
    282 => 2,
    283 => 2,
    284 => 2,
    285 => 2,
    286 => 2,
    287 => 2,
    288 => 2,
    289 => 2,
    290 => 2,
    291 => 2,
    292 => 2,
    293 => 2,
    294 => 2,
    295 => 2,
    296 => 2,
    297 => 2,
    298 => 2,
    299 => 2,
    300 => 2,
    301 => 2,
    302 => 2,
    303 => 2,
    304 => 2,
    305 => 2,
    306 => 2,
    307 => 2,
    308 => 2,
    309 => 2,
    310 => 2,
    311 => 2,
    312 => 2,
    313 => 2,
    314 => 2,
    315 => 2,
    316 => 2,
    317 => 2,
    318 => 2,
    319 => 2,
    320 => 2,
    321 => 2,
    322 => 2,
    323 => 2,
    324 => 2,
    325 => 2,
    326 => 2,
    327 => 2,
    328 => 2,
    329 => 2,
    330 => 2,
    331 => 2,
    332 => 2,
    333 => 2,
    334 => 2,
    335 => 2,
    336 => 2,
    337 => 2,
    338 => 2,
    339 => 2,
    340 => 2,
    341 => 2,
    342 => 2,
    343 => 2,
    344 => 2,
    345 => 2,
    346 => 2,
    347 => 2,
    348 => 2,
    349 => 2,
    350 => 2,
    351 => 2,
    352 => 2,
    353 => 2,
    354 => 2,
    355 => 2,
    356 => 2,
    357 => 2,
    358 => 2,
    359 => 2,
    360 => 2,
    361 => 2,
    362 => 2,
    363 => 2,
    364 => 2,
    365 => 2,
    366 => 2,
    367 => 2,
    368 => 2,
    369 => 2,
    370 => 2,
    371 => 2,
    372 => 2,
    373 => 2,
    374 => 2,
    375 => 2,
    376 => 2,
    377 => 2,
    378 => 2,
    379 => 2,
    380 => 2,
    381 => 2,
    382 => 2,
    383 => 2,
    384 => 2,
    385 => 2,
    386 => 2,
    387 => 2,
    388 => 2,
    389 => 2,
    390 => 2,
    391 => 2,
    392 => 2,
    393 => 2,
    394 => 2,
    395 => 2,
    396 => 2,
    397 => 2,
    398 => 2,
    399 => 2,
    400 => 2,
    401 => 2,
    402 => 2,
    403 => 2,
    404 => 2,
    405 => 2,
    406 => 2,
    407 => 2,
    408 => 2,
    409 => 2,
    410 => 2,
    411 => 2,
    412 => 2,
    413 => 2,
    414 => 2,
    415 => 3,
    416 => 3,
    417 => 3,
    418 => 3,
    419 => 3,
    420 => 3,
    421 => 3,
    422 => 3,
    423 => 3,
    424 => 3,
    425 => 3,
    426 => 3,
    427 => 3,
    428 => 3,
    429 => 3,
    430 => 3,
    431 => 3,
    432 => 3,
    433 => 3,
    434 => 3,
    435 => 3,
    436 => 3,
    437 => 3,
    438 => 3,
    439 => 3,
    440 => 3,
    441 => 3,
    442 => 3,
    443 => 3,
    444 => 3,
    445 => 3,
    446 => 3,
    447 => 3,
    448 => 3,
    449 => 3,
    450 => 3,
    451 => 3,
    452 => 3,
    453 => 3,
    454 => 3,
    455 => 3,
    456 => 3,
    457 => 3,
    458 => 3,
    459 => 3,
    460 => 3,
    461 => 3,
    462 => 3,
    463 => 3,
    464 => 3,
    465 => 3,
    466 => 3,
    467 => 3,
    468 => 3,
    469 => 3,
    470 => 3,
    471 => 3,
    472 => 3,
    473 => 3,
    474 => 3,
    475 => 3,
    476 => 3,
    477 => 3,
    478 => 3,
    479 => 3,
    480 => 3,
    481 => 3,
    482 => 3,
    483 => 3,
    484 => 3,
    485 => 3,
    486 => 3,
    487 => 3,
    488 => 3,
    489 => 3,
    490 => 3,
    491 => 3,
    492 => 3,
    493 => 3,
    494 => 3,
    495 => 3,
    496 => 3,
    497 => 3,
    498 => 3,
    499 => 3,
    500 => 3,
    501 => 3,
    502 => 3,
    503 => 3,
    504 => 3,
    505 => 3,
    506 => 3,
    507 => 3,
    508 => 3,
    509 => 3,
    510 => 3,
    511 => 3,
    512 => 3,
    513 => 3,
    514 => 3,
    515 => 3,
    516 => 3,
    517 => 3,
    518 => 3,
    519 => 3,
    520 => 3,
    521 => 3,
    522 => 3,
    523 => 3,
    524 => 3,
    525 => 3,
    526 => 3,
    527 => 3,
    528 => 3,
    529 => 3,
    530 => 3,
    531 => 3,
    532 => 3,
    533 => 3,
    534 => 3,
    535 => 3,
    536 => 3,
    537 => 3,
    538 => 3,
    539 => 3,
    540 => 3,
    541 => 3,
    542 => 3,
    543 => 3,
    544 => 3,
    545 => 3,
    546 => 3,
    547 => 3,
    548 => 3,
    549 => 3,
    550 => 3,
    551 => 3,
    552 => 3,
    553 => 3,
    554 => 3,
    555 => 3,
    556 => 3,
    557 => 3,
    558 => 3,
    559 => 3,
    560 => 3,
    561 => 3,
    562 => 3,
    563 => 3,
    564 => 3,
    565 => 3,
    566 => 3,
    567 => 3,
    568 => 3,
    569 => 3,
    570 => 3,
    571 => 3,
    572 => 3,
    573 => 3,
    574 => 3,
    575 => 3,
    576 => 3,
    577 => 3,
    578 => 3,
    579 => 3,
    580 => 4,
    581 => 4,
    582 => 4,
    583 => 4,
    584 => 4,
    585 => 4,
    586 => 4,
    587 => 4,
    588 => 4,
    589 => 4,
    590 => 4,
    591 => 4,
    592 => 4,
    593 => 4,
    594 => 4,
    595 => 4,
    596 => 4,
    597 => 4,
    598 => 4,
    599 => 4,
    600 => 4,
    601 => 4,
    602 => 4,
    603 => 4,
    604 => 4,
    605 => 4,
    606 => 4,
    607 => 4,
    608 => 4,
    609 => 4,
    610 => 4,
    611 => 4,
    612 => 4,
    613 => 4,
    614 => 4,
    615 => 4,
    616 => 4,
    617 => 4,
    618 => 4,
    619 => 4,
    620 => 4,
    621 => 4,
    622 => 4,
    623 => 4,
    624 => 4,
    625 => 4,
    626 => 4,
    627 => 4,
    628 => 4,
    629 => 4,
    630 => 4,
    631 => 4,
    632 => 4,
    633 => 4,
    634 => 4,
    635 => 4,
    636 => 4,
    637 => 4,
    638 => 4,
    639 => 4,
    640 => 4,
    641 => 4,
    642 => 4,
    643 => 4,
    644 => 4,
    645 => 4,
    646 => 4,
    647 => 4,
    648 => 4,
    649 => 4,
    650 => 4,
    651 => 4,
    652 => 4,
    653 => 4,
    654 => 4,
    655 => 4,
    656 => 4,
    657 => 4,
    658 => 4,
    659 => 4,
    660 => 4,
    661 => 4,
    662 => 4,
    663 => 4,
    664 => 4,
    665 => 4,
    666 => 4,
    667 => 4,
    668 => 4,
    669 => 4,
    670 => 4,
    671 => 4,
    672 => 4,
    673 => 4,
    674 => 4,
    675 => 4,
    676 => 4,
    677 => 4,
    678 => 4,
    679 => 4,
    680 => 4,
    681 => 4,
    682 => 4,
    683 => 4,
    684 => 4,
    685 => 4,
    686 => 4,
    687 => 4,
    688 => 4,
    689 => 4,
    690 => 4,
    691 => 4,
    692 => 4,
    693 => 4,
    694 => 4,
    695 => 4,
    696 => 4,
    697 => 4,
    698 => 4,
    699 => 4,
    700 => 4,
    701 => 4,
    702 => 4,
    703 => 4,
    704 => 4,
    705 => 4,
    706 => 4,
    707 => 4,
    708 => 4,
    709 => 4,
    710 => 4,
    711 => 4,
    712 => 4,
    713 => 4,
    714 => 4,
    715 => 4,
    716 => 4,
    717 => 4,
    718 => 4,
    719 => 4,
    720 => 4,
    721 => 4,
    722 => 4,
    723 => 4,
    724 => 4,
    725 => 4,
    726 => 4,
    727 => 4,
    728 => 4,
    729 => 4,
    730 => 4,
    731 => 4,
    732 => 4,
    733 => 4,
    734 => 4,
    735 => 4,
    736 => 4,
    737 => 4,
    738 => 4,
    739 => 4,
    740 => 4,
    741 => 4,
    742 => 4,
    743 => 4,
    744 => 4,
    745 => 4,
    746 => 5,
    747 => 5,
    748 => 5,
    749 => 5,
    750 => 5,
    751 => 5,
    752 => 5,
    753 => 5,
    754 => 5,
    755 => 5,
    756 => 5,
    757 => 5,
    758 => 5,
    759 => 5,
    760 => 5,
    761 => 5,
    762 => 5,
    763 => 5,
    764 => 5,
    765 => 5,
    766 => 5,
    767 => 5,
    768 => 5,
    769 => 5,
    770 => 5,
    771 => 5,
    772 => 5,
    773 => 5,
    774 => 5,
    775 => 5,
    776 => 5,
    777 => 5,
    778 => 5,
    779 => 5,
    780 => 5,
    781 => 5,
    782 => 5,
    783 => 5,
    784 => 5,
    785 => 5,
    786 => 5,
    787 => 5,
    788 => 5,
    789 => 5,
    790 => 5,
    791 => 5,
    792 => 5,
    793 => 5,
    794 => 5,
    795 => 5,
    796 => 5,
    797 => 5,
    798 => 5,
    799 => 5,
    800 => 5,
    801 => 5,
    802 => 5,
    803 => 5,
    804 => 5,
    805 => 5,
    806 => 5,
    807 => 5,
    808 => 5,
    809 => 5,
    810 => 5,
    811 => 5,
    812 => 5,
    813 => 5,
    814 => 5,
    815 => 5,
    816 => 5,
    817 => 5,
    818 => 5,
    819 => 5,
    820 => 5,
    821 => 5,
    822 => 5,
    823 => 5,
    824 => 5,
    825 => 5,
    826 => 5,
    827 => 5,
    828 => 5,
    829 => 5,
    830 => 5,
    831 => 5,
    832 => 5,
    833 => 5,
    834 => 5,
    835 => 5,
    836 => 5,
    837 => 5,
    838 => 5,
    839 => 5,
    840 => 5,
    841 => 5,
    842 => 5,
    843 => 5,
    844 => 5,
    845 => 5,
    846 => 5,
    847 => 5,
    848 => 5,
    849 => 5,
    850 => 5,
    851 => 5,
    852 => 5,
    853 => 5,
    854 => 5,
    855 => 5,
    856 => 5,
    857 => 5,
    858 => 5,
    859 => 5,
    860 => 5,
    861 => 5,
    862 => 5,
    863 => 5,
    864 => 5,
    865 => 5,
    866 => 5,
    867 => 5,
    868 => 5,
    869 => 5,
    870 => 5,
    871 => 5,
    872 => 5,
    873 => 5,
    874 => 5,
    875 => 5,
    876 => 5,
    877 => 5,
    878 => 5,
    879 => 5,
    880 => 5,
    881 => 5,
    882 => 5,
    883 => 5,
    884 => 5,
    885 => 5,
    886 => 5,
    887 => 5,
    888 => 5,
    889 => 5,
    890 => 5,
    891 => 5,
    892 => 5,
    893 => 5,
    894 => 5,
    895 => 5,
    896 => 5,
    897 => 5,
    898 => 5,
    899 => 5,
    900 => 5,
    901 => 5,
    902 => 5,
    903 => 5,
    904 => 5,
    905 => 5,
    906 => 5,
    907 => 5,
    908 => 5,
    909 => 5,
    910 => 5,
    911 => 5,
    912 => 6,
    913 => 6,
    914 => 6,
    915 => 6,
    916 => 6,
    917 => 6,
    918 => 6,
    919 => 6,
    920 => 6,
    921 => 6,
    922 => 6,
    923 => 6,
    924 => 6,
    925 => 6,
    926 => 6,
    927 => 6,
    928 => 6,
    929 => 6,
    930 => 6,
    931 => 6,
    932 => 6,
    933 => 6,
    934 => 6,
    935 => 6,
    936 => 6,
    937 => 6,
    938 => 6,
    939 => 6,
    940 => 6,
    941 => 6,
    942 => 6,
    943 => 6,
    944 => 6,
    945 => 6,
    946 => 6,
    947 => 6,
    948 => 6,
    949 => 6,
    950 => 6,
    951 => 6,
    952 => 6,
    953 => 6,
    954 => 6,
    955 => 6,
    956 => 6,
    957 => 6,
    958 => 6,
    959 => 6,
    960 => 6,
    961 => 6,
    962 => 6,
    963 => 6,
    964 => 6,
    965 => 6,
    966 => 6,
    967 => 6,
    968 => 6,
    969 => 6,
    970 => 6,
    971 => 6,
    972 => 6,
    973 => 6,
    974 => 6,
    975 => 6,
    976 => 6,
    977 => 6,
    978 => 6,
    979 => 6,
    980 => 6,
    981 => 6,
    982 => 6,
    983 => 6,
    984 => 6,
    985 => 6,
    986 => 6,
    987 => 6,
    988 => 6,
    989 => 6,
    990 => 6,
    991 => 6,
    992 => 6,
    993 => 6,
    994 => 6,
    995 => 6,
    996 => 6,
    997 => 6,
    998 => 6,
    999 => 6,
    1000 => 6,
    1001 => 6,
    1002 => 6,
    1003 => 6,
    1004 => 6,
    1005 => 6,
    1006 => 6,
    1007 => 6,
    1008 => 6,
    1009 => 6,
    1010 => 6,
    1011 => 6,
    1012 => 6,
    1013 => 6,
    1014 => 6,
    1015 => 6,
    1016 => 6,
    1017 => 6,
    1018 => 6,
    1019 => 6,
    1020 => 6,
    1021 => 6,
    1022 => 6,
    1023 => 6,
    1024 => 6,
    1025 => 6,
    1026 => 6,
    1027 => 6,
    1028 => 6,
    1029 => 6,
    1030 => 6,
    1031 => 6,
    1032 => 6,
    1033 => 6,
    1034 => 6,
    1035 => 6,
    1036 => 6,
    1037 => 6,
    1038 => 6,
    1039 => 6,
    1040 => 6,
    1041 => 6,
    1042 => 6,
    1043 => 6,
    1044 => 6,
    1045 => 6,
    1046 => 6,
    1047 => 6,
    1048 => 6,
    1049 => 6,
    1050 => 6,
    1051 => 6,
    1052 => 6,
    1053 => 6,
    1054 => 6,
    1055 => 6,
    1056 => 6,
    1057 => 6,
    1058 => 6,
    1059 => 6,
    1060 => 6,
    1061 => 6,
    1062 => 6,
    1063 => 6,
    1064 => 6,
    1065 => 6,
    1066 => 6,
    1067 => 6,
    1068 => 6,
    1069 => 6,
    1070 => 6,
    1071 => 6,
    1072 => 6,
    1073 => 6,
    1074 => 6,
    1075 => 6,
    1076 => 6,
    1077 => 6,
    1078 => 6,
    1079 => 7,
    1080 => 7,
    1081 => 7,
    1082 => 7,
    1083 => 7,
    1084 => 7,
    1085 => 7,
    1086 => 7,
    1087 => 7,
    1088 => 7,
    1089 => 7,
    1090 => 7,
    1091 => 7,
    1092 => 7,
    1093 => 7,
    1094 => 7,
    1095 => 7,
    1096 => 7,
    1097 => 7,
    1098 => 7,
    1099 => 7,
    1100 => 7,
    1101 => 7,
    1102 => 7,
    1103 => 7,
    1104 => 7,
    1105 => 7,
    1106 => 7,
    1107 => 7,
    1108 => 7,
    1109 => 7,
    1110 => 7,
    1111 => 7,
    1112 => 7,
    1113 => 7,
    1114 => 7,
    1115 => 7,
    1116 => 7,
    1117 => 7,
    1118 => 7,
    1119 => 7,
    1120 => 7,
    1121 => 7,
    1122 => 7,
    1123 => 7,
    1124 => 7,
    1125 => 7,
    1126 => 7,
    1127 => 7,
    1128 => 7,
    1129 => 7,
    1130 => 7,
    1131 => 7,
    1132 => 7,
    1133 => 7,
    1134 => 7,
    1135 => 7,
    1136 => 7,
    1137 => 7,
    1138 => 7,
    1139 => 7,
    1140 => 7,
    1141 => 7,
    1142 => 7,
    1143 => 7,
    1144 => 7,
    1145 => 7,
    1146 => 7,
    1147 => 7,
    1148 => 7,
    1149 => 7,
    1150 => 7,
    1151 => 7,
    1152 => 7,
    1153 => 7,
    1154 => 7,
    1155 => 7,
    1156 => 7,
    1157 => 7,
    1158 => 7,
    1159 => 7,
    1160 => 7,
    1161 => 7,
    1162 => 7,
    1163 => 7,
    1164 => 7,
    1165 => 7,
    1166 => 7,
    1167 => 7,
    1168 => 7,
    1169 => 7,
    1170 => 7,
    1171 => 7,
    1172 => 7,
    1173 => 7,
    1174 => 7,
    1175 => 7,
    1176 => 7,
    1177 => 7,
    1178 => 7,
    1179 => 7,
    1180 => 7,
    1181 => 7,
    1182 => 7,
    1183 => 7,
    1184 => 7,
    1185 => 7,
    1186 => 7,
    1187 => 7,
    1188 => 7,
    1189 => 7,
    1190 => 7,
    1191 => 7,
    1192 => 7,
    1193 => 7,
    1194 => 7,
    1195 => 7,
    1196 => 7,
    1197 => 7,
    1198 => 7,
    1199 => 7,
    1200 => 7,
    1201 => 7,
    1202 => 7,
    1203 => 7,
    1204 => 7,
    1205 => 7,
    1206 => 7,
    1207 => 7,
    1208 => 7,
    1209 => 7,
    1210 => 7,
    1211 => 7,
    1212 => 7,
    1213 => 7,
    1214 => 7,
    1215 => 7,
    1216 => 7,
    1217 => 7,
    1218 => 7,
    1219 => 7,
    1220 => 7,
    1221 => 7,
    1222 => 7,
    1223 => 7,
    1224 => 7,
    1225 => 7,
    1226 => 7,
    1227 => 7,
    1228 => 7,
    1229 => 7,
    1230 => 7,
    1231 => 7,
    1232 => 7,
    1233 => 7,
    1234 => 7,
    1235 => 7,
    1236 => 7,
    1237 => 7,
    1238 => 7,
    1239 => 7,
    1240 => 7,
    1241 => 7,
    1242 => 7,
    1243 => 7,
    1244 => 7,
    1245 => 8,
    1246 => 8,
    1247 => 8,
    1248 => 8,
    1249 => 8,
    1250 => 8,
    1251 => 8,
    1252 => 8,
    1253 => 8,
    1254 => 8,
    1255 => 8,
    1256 => 8,
    1257 => 8,
    1258 => 8,
    1259 => 8,
    1260 => 8,
    1261 => 8,
    1262 => 8,
    1263 => 8,
    1264 => 8,
    1265 => 8,
    1266 => 8,
    1267 => 8,
    1268 => 8,
    1269 => 8,
    1270 => 8,
    1271 => 8,
    1272 => 8,
    1273 => 8,
    1274 => 8,
    1275 => 8,
    1276 => 8,
    1277 => 8,
    1278 => 8,
    1279 => 8,
    1280 => 8,
    1281 => 8,
    1282 => 8,
    1283 => 8,
    1284 => 8,
    1285 => 8,
    1286 => 8,
    1287 => 8,
    1288 => 8,
    1289 => 8,
    1290 => 8,
    1291 => 8,
    1292 => 8,
    1293 => 8,
    1294 => 8,
    1295 => 8,
    1296 => 8,
    1297 => 8,
    1298 => 8,
    1299 => 8,
    1300 => 8,
    1301 => 8,
    1302 => 8,
    1303 => 8,
    1304 => 8,
    1305 => 8,
    1306 => 8,
    1307 => 8,
    1308 => 8,
    1309 => 8,
    1310 => 8,
    1311 => 8,
    1312 => 8,
    1313 => 8,
    1314 => 8,
    1315 => 8,
    1316 => 8,
    1317 => 8,
    1318 => 8,
    1319 => 8,
    1320 => 8,
    1321 => 8,
    1322 => 8,
    1323 => 8,
    1324 => 8,
    1325 => 8,
    1326 => 8,
    1327 => 8,
    1328 => 8,
    1329 => 8,
    1330 => 8,
    1331 => 8,
    1332 => 8,
    1333 => 8,
    1334 => 8,
    1335 => 8,
    1336 => 8,
    1337 => 8,
    1338 => 8,
    1339 => 8,
    1340 => 8,
    1341 => 8,
    1342 => 8,
    1343 => 8,
    1344 => 8,
    1345 => 8,
    1346 => 8,
    1347 => 8,
    1348 => 8,
    1349 => 8,
    1350 => 8,
    1351 => 8,
    1352 => 8,
    1353 => 8,
    1354 => 8,
    1355 => 8,
    1356 => 8,
    1357 => 8,
    1358 => 8,
    1359 => 8,
    1360 => 8,
    1361 => 8,
    1362 => 8,
    1363 => 8,
    1364 => 8,
    1365 => 8,
    1366 => 8,
    1367 => 8,
    1368 => 8,
    1369 => 8,
    1370 => 8,
    1371 => 8,
    1372 => 8,
    1373 => 8,
    1374 => 8,
    1375 => 8,
    1376 => 8,
    1377 => 8,
    1378 => 8,
    1379 => 8,
    1380 => 8,
    1381 => 8,
    1382 => 8,
    1383 => 8,
    1384 => 8,
    1385 => 8,
    1386 => 8,
    1387 => 8,
    1388 => 8,
    1389 => 8,
    1390 => 8,
    1391 => 8,
    1392 => 8,
    1393 => 8,
    1394 => 8,
    1395 => 8,
    1396 => 8,
    1397 => 8,
    1398 => 8,
    1399 => 8,
    1400 => 8,
    1401 => 8,
    1402 => 8,
    1403 => 8,
    1404 => 8,
    1405 => 8,
    1406 => 8,
    1407 => 8,
    1408 => 8,
    1409 => 8,
    1410 => 8,
    1411 => 8,
    1412 => 9,
    1413 => 9,
    1414 => 9,
    1415 => 9,
    1416 => 9,
    1417 => 9,
    1418 => 9,
    1419 => 9,
    1420 => 9,
    1421 => 9,
    1422 => 9,
    1423 => 9,
    1424 => 9,
    1425 => 9,
    1426 => 9,
    1427 => 9,
    1428 => 9,
    1429 => 9,
    1430 => 9,
    1431 => 9,
    1432 => 9,
    1433 => 9,
    1434 => 9,
    1435 => 9,
    1436 => 9,
    1437 => 9,
    1438 => 9,
    1439 => 9,
    1440 => 9,
    1441 => 9,
    1442 => 9,
    1443 => 9,
    1444 => 9,
    1445 => 9,
    1446 => 9,
    1447 => 9,
    1448 => 9,
    1449 => 9,
    1450 => 9,
    1451 => 9,
    1452 => 9,
    1453 => 9,
    1454 => 9,
    1455 => 9,
    1456 => 9,
    1457 => 9,
    1458 => 9,
    1459 => 9,
    1460 => 9,
    1461 => 9,
    1462 => 9,
    1463 => 9,
    1464 => 9,
    1465 => 9,
    1466 => 9,
    1467 => 9,
    1468 => 9,
    1469 => 9,
    1470 => 9,
    1471 => 9,
    1472 => 9,
    1473 => 9,
    1474 => 9,
    1475 => 9,
    1476 => 9,
    1477 => 9,
    1478 => 9,
    1479 => 9,
    1480 => 9,
    1481 => 9,
    1482 => 9,
    1483 => 9,
    1484 => 9,
    1485 => 9,
    1486 => 9,
    1487 => 9,
    1488 => 9,
    1489 => 9,
    1490 => 9,
    1491 => 9,
    1492 => 9,
    1493 => 9,
    1494 => 9,
    1495 => 9,
    1496 => 9,
    1497 => 9,
    1498 => 9,
    1499 => 9,
    1500 => 9,
    1501 => 9,
    1502 => 9,
    1503 => 9,
    1504 => 9,
    1505 => 9,
    1506 => 9,
    1507 => 9,
    1508 => 9,
    1509 => 9,
    1510 => 9,
    1511 => 9,
    1512 => 9,
    1513 => 9,
    1514 => 9,
    1515 => 9,
    1516 => 9,
    1517 => 9,
    1518 => 9,
    1519 => 9,
    1520 => 9,
    1521 => 9,
    1522 => 9,
    1523 => 9,
    1524 => 9,
    1525 => 9,
    1526 => 9,
    1527 => 9,
    1528 => 9,
    1529 => 9,
    1530 => 9,
    1531 => 9,
    1532 => 9,
    1533 => 9,
    1534 => 9,
    1535 => 9,
    1536 => 9,
    1537 => 9,
    1538 => 9,
    1539 => 9,
    1540 => 9,
    1541 => 9,
    1542 => 9,
    1543 => 9,
    1544 => 9,
    1545 => 9,
    1546 => 9,
    1547 => 9,
    1548 => 9,
    1549 => 9,
    1550 => 9,
    1551 => 9,
    1552 => 9,
    1553 => 9,
    1554 => 9,
    1555 => 9,
    1556 => 9,
    1557 => 9,
    1558 => 9,
    1559 => 9,
    1560 => 9,
    1561 => 9,
    1562 => 9,
    1563 => 9,
    1564 => 9,
    1565 => 9,
    1566 => 9,
    1567 => 9,
    1568 => 9,
    1569 => 9,
    1570 => 9,
    1571 => 9,
    1572 => 9,
    1573 => 9,
    1574 => 9,
    1575 => 9,
    1576 => 9,
    1577 => 9,
    1578 => 9,
    1579 => 10,
    1580 => 10,
    1581 => 10,
    1582 => 10,
    1583 => 10,
    1584 => 10,
    1585 => 10,
    1586 => 10,
    1587 => 10,
    1588 => 10,
    1589 => 10,
    1590 => 10,
    1591 => 10,
    1592 => 10,
    1593 => 10,
    1594 => 10,
    1595 => 10,
    1596 => 10,
    1597 => 10,
    1598 => 10,
    1599 => 10,
    1600 => 10,
    1601 => 10,
    1602 => 10,
    1603 => 10,
    1604 => 10,
    1605 => 10,
    1606 => 10,
    1607 => 10,
    1608 => 10,
    1609 => 10,
    1610 => 10,
    1611 => 10,
    1612 => 10,
    1613 => 10,
    1614 => 10,
    1615 => 10,
    1616 => 10,
    1617 => 10,
    1618 => 10,
    1619 => 10,
    1620 => 10,
    1621 => 10,
    1622 => 10,
    1623 => 10,
    1624 => 10,
    1625 => 10,
    1626 => 10,
    1627 => 10,
    1628 => 10,
    1629 => 10,
    1630 => 10,
    1631 => 10,
    1632 => 10,
    1633 => 10,
    1634 => 10,
    1635 => 10,
    1636 => 10,
    1637 => 10,
    1638 => 10,
    1639 => 10,
    1640 => 10,
    1641 => 10,
    1642 => 10,
    1643 => 10,
    1644 => 10,
    1645 => 10,
    1646 => 10,
    1647 => 10,
    1648 => 10,
    1649 => 10,
    1650 => 10,
    1651 => 10,
    1652 => 10,
    1653 => 10,
    1654 => 10,
    1655 => 10,
    1656 => 10,
    1657 => 10,
    1658 => 10,
    1659 => 10,
    1660 => 10,
    1661 => 10,
    1662 => 10,
    1663 => 10,
    1664 => 10,
    1665 => 10,
    1666 => 10,
    1667 => 10,
    1668 => 10,
    1669 => 10,
    1670 => 10,
    1671 => 10,
    1672 => 10,
    1673 => 10,
    1674 => 10,
    1675 => 10,
    1676 => 10,
    1677 => 10,
    1678 => 10,
    1679 => 10,
    1680 => 10,
    1681 => 10,
    1682 => 10,
    1683 => 10,
    1684 => 10,
    1685 => 10,
    1686 => 10,
    1687 => 10,
    1688 => 10,
    1689 => 10,
    1690 => 10,
    1691 => 10,
    1692 => 10,
    1693 => 10,
    1694 => 10,
    1695 => 10,
    1696 => 10,
    1697 => 10,
    1698 => 10,
    1699 => 10,
    1700 => 10,
    1701 => 10,
    1702 => 10,
    1703 => 10,
    1704 => 10,
    1705 => 10,
    1706 => 10,
    1707 => 10,
    1708 => 10,
    1709 => 10,
    1710 => 10,
    1711 => 10,
    1712 => 10,
    1713 => 10,
    1714 => 10,
    1715 => 10,
    1716 => 10,
    1717 => 10,
    1718 => 10,
    1719 => 10,
    1720 => 10,
    1721 => 10,
    1722 => 10,
    1723 => 10,
    1724 => 10,
    1725 => 10,
    1726 => 10,
    1727 => 10,
    1728 => 10,
    1729 => 10,
    1730 => 10,
    1731 => 10,
    1732 => 10,
    1733 => 10,
    1734 => 10,
    1735 => 10,
    1736 => 10,
    1737 => 10,
    1738 => 10,
    1739 => 10,
    1740 => 10,
    1741 => 10,
    1742 => 10,
    1743 => 10,
    1744 => 10,
    1745 => 10,
    1746 => 10,
    1747 => 11,
    1748 => 11,
    1749 => 11,
    1750 => 11,
    1751 => 11,
    1752 => 11,
    1753 => 11,
    1754 => 11,
    1755 => 11,
    1756 => 11,
    1757 => 11,
    1758 => 11,
    1759 => 11,
    1760 => 11,
    1761 => 11,
    1762 => 11,
    1763 => 11,
    1764 => 11,
    1765 => 11,
    1766 => 11,
    1767 => 11,
    1768 => 11,
    1769 => 11,
    1770 => 11,
    1771 => 11,
    1772 => 11,
    1773 => 11,
    1774 => 11,
    1775 => 11,
    1776 => 11,
    1777 => 11,
    1778 => 11,
    1779 => 11,
    1780 => 11,
    1781 => 11,
    1782 => 11,
    1783 => 11,
    1784 => 11,
    1785 => 11,
    1786 => 11,
    1787 => 11,
    1788 => 11,
    1789 => 11,
    1790 => 11,
    1791 => 11,
    1792 => 11,
    1793 => 11,
    1794 => 11,
    1795 => 11,
    1796 => 11,
    1797 => 11,
    1798 => 11,
    1799 => 11,
    1800 => 11,
    1801 => 11,
    1802 => 11,
    1803 => 11,
    1804 => 11,
    1805 => 11,
    1806 => 11,
    1807 => 11,
    1808 => 11,
    1809 => 11,
    1810 => 11,
    1811 => 11,
    1812 => 11,
    1813 => 11,
    1814 => 11,
    1815 => 11,
    1816 => 11,
    1817 => 11,
    1818 => 11,
    1819 => 11,
    1820 => 11,
    1821 => 11,
    1822 => 11,
    1823 => 11,
    1824 => 11,
    1825 => 11,
    1826 => 11,
    1827 => 11,
    1828 => 11,
    1829 => 11,
    1830 => 11,
    1831 => 11,
    1832 => 11,
    1833 => 11,
    1834 => 11,
    1835 => 11,
    1836 => 11,
    1837 => 11,
    1838 => 11,
    1839 => 11,
    1840 => 11,
    1841 => 11,
    1842 => 11,
    1843 => 11,
    1844 => 11,
    1845 => 11,
    1846 => 11,
    1847 => 11,
    1848 => 11,
    1849 => 11,
    1850 => 11,
    1851 => 11,
    1852 => 11,
    1853 => 11,
    1854 => 11,
    1855 => 11,
    1856 => 11,
    1857 => 11,
    1858 => 11,
    1859 => 11,
    1860 => 11,
    1861 => 11,
    1862 => 11,
    1863 => 11,
    1864 => 11,
    1865 => 11,
    1866 => 11,
    1867 => 11,
    1868 => 11,
    1869 => 11,
    1870 => 11,
    1871 => 11,
    1872 => 11,
    1873 => 11,
    1874 => 11,
    1875 => 11,
    1876 => 11,
    1877 => 11,
    1878 => 11,
    1879 => 11,
    1880 => 11,
    1881 => 11,
    1882 => 11,
    1883 => 11,
    1884 => 11,
    1885 => 11,
    1886 => 11,
    1887 => 11,
    1888 => 11,
    1889 => 11,
    1890 => 11,
    1891 => 11,
    1892 => 11,
    1893 => 11,
    1894 => 11,
    1895 => 11,
    1896 => 11,
    1897 => 11,
    1898 => 11,
    1899 => 11,
    1900 => 11,
    1901 => 11,
    1902 => 11,
    1903 => 11,
    1904 => 11,
    1905 => 11,
    1906 => 11,
    1907 => 11,
    1908 => 11,
    1909 => 11,
    1910 => 11,
    1911 => 11,
    1912 => 11,
    1913 => 11,
    1914 => 11,
    1915 => 12,
    1916 => 12,
    1917 => 12,
    1918 => 12,
    1919 => 12,
    1920 => 12,
    1921 => 12,
    1922 => 12,
    1923 => 12,
    1924 => 12,
    1925 => 12,
    1926 => 12,
    1927 => 12,
    1928 => 12,
    1929 => 12,
    1930 => 12,
    1931 => 12,
    1932 => 12,
    1933 => 12,
    1934 => 12,
    1935 => 12,
    1936 => 12,
    1937 => 12,
    1938 => 12,
    1939 => 12,
    1940 => 12,
    1941 => 12,
    1942 => 12,
    1943 => 12,
    1944 => 12,
    1945 => 12,
    1946 => 12,
    1947 => 12,
    1948 => 12,
    1949 => 12,
    1950 => 12,
    1951 => 12,
    1952 => 12,
    1953 => 12,
    1954 => 12,
    1955 => 12,
    1956 => 12,
    1957 => 12,
    1958 => 12,
    1959 => 12,
    1960 => 12,
    1961 => 12,
    1962 => 12,
    1963 => 12,
    1964 => 12,
    1965 => 12,
    1966 => 12,
    1967 => 12,
    1968 => 12,
    1969 => 12,
    1970 => 12,
    1971 => 12,
    1972 => 12,
    1973 => 12,
    1974 => 12,
    1975 => 12,
    1976 => 12,
    1977 => 12,
    1978 => 12,
    1979 => 12,
    1980 => 12,
    1981 => 12,
    1982 => 12,
    1983 => 12,
    1984 => 12,
    1985 => 12,
    1986 => 12,
    1987 => 12,
    1988 => 12,
    1989 => 12,
    1990 => 12,
    1991 => 12,
    1992 => 12,
    1993 => 12,
    1994 => 12,
    1995 => 12,
    1996 => 12,
    1997 => 12,
    1998 => 12,
    1999 => 12,
    2000 => 12,
    2001 => 12,
    2002 => 12,
    2003 => 12,
    2004 => 12,
    2005 => 12,
    2006 => 12,
    2007 => 12,
    2008 => 12,
    2009 => 12,
    2010 => 12,
    2011 => 12,
    2012 => 12,
    2013 => 12,
    2014 => 12,
    2015 => 12,
    2016 => 12,
    2017 => 12,
    2018 => 12,
    2019 => 12,
    2020 => 12,
    2021 => 12,
    2022 => 12,
    2023 => 12,
    2024 => 12,
    2025 => 12,
    2026 => 12,
    2027 => 12,
    2028 => 12,
    2029 => 12,
    2030 => 12,
    2031 => 12,
    2032 => 12,
    2033 => 12,
    2034 => 12,
    2035 => 12,
    2036 => 12,
    2037 => 12,
    2038 => 12,
    2039 => 12,
    2040 => 12,
    2041 => 12,
    2042 => 12,
    2043 => 12,
    2044 => 12,
    2045 => 12,
    2046 => 12,
    2047 => 12,
    2048 => 12,
    2049 => 12,
    2050 => 12,
    2051 => 12,
    2052 => 12,
    2053 => 12,
    2054 => 12,
    2055 => 12,
    2056 => 12,
    2057 => 12,
    2058 => 12,
    2059 => 12,
    2060 => 12,
    2061 => 12,
    2062 => 12,
    2063 => 12,
    2064 => 12,
    2065 => 12,
    2066 => 12,
    2067 => 12,
    2068 => 12,
    2069 => 12,
    2070 => 12,
    2071 => 12,
    2072 => 12,
    2073 => 12,
    2074 => 12,
    2075 => 12,
    2076 => 12,
    2077 => 12,
    2078 => 12,
    2079 => 12,
    2080 => 12,
    2081 => 12,
    2082 => 12,
    2083 => 12,
    2084 => 13,
    2085 => 13,
    2086 => 13,
    2087 => 13,
    2088 => 13,
    2089 => 13,
    2090 => 13,
    2091 => 13,
    2092 => 13,
    2093 => 13,
    2094 => 13,
    2095 => 13,
    2096 => 13,
    2097 => 13,
    2098 => 13,
    2099 => 13,
    2100 => 13,
    2101 => 13,
    2102 => 13,
    2103 => 13,
    2104 => 13,
    2105 => 13,
    2106 => 13,
    2107 => 13,
    2108 => 13,
    2109 => 13,
    2110 => 13,
    2111 => 13,
    2112 => 13,
    2113 => 13,
    2114 => 13,
    2115 => 13,
    2116 => 13,
    2117 => 13,
    2118 => 13,
    2119 => 13,
    2120 => 13,
    2121 => 13,
    2122 => 13,
    2123 => 13,
    2124 => 13,
    2125 => 13,
    2126 => 13,
    2127 => 13,
    2128 => 13,
    2129 => 13,
    2130 => 13,
    2131 => 13,
    2132 => 13,
    2133 => 13,
    2134 => 13,
    2135 => 13,
    2136 => 13,
    2137 => 13,
    2138 => 13,
    2139 => 13,
    2140 => 13,
    2141 => 13,
    2142 => 13,
    2143 => 13,
    2144 => 13,
    2145 => 13,
    2146 => 13,
    2147 => 13,
    2148 => 13,
    2149 => 13,
    2150 => 13,
    2151 => 13,
    2152 => 13,
    2153 => 13,
    2154 => 13,
    2155 => 13,
    2156 => 13,
    2157 => 13,
    2158 => 13,
    2159 => 13,
    2160 => 13,
    2161 => 13,
    2162 => 13,
    2163 => 13,
    2164 => 13,
    2165 => 13,
    2166 => 13,
    2167 => 13,
    2168 => 13,
    2169 => 13,
    2170 => 13,
    2171 => 13,
    2172 => 13,
    2173 => 13,
    2174 => 13,
    2175 => 13,
    2176 => 13,
    2177 => 13,
    2178 => 13,
    2179 => 13,
    2180 => 13,
    2181 => 13,
    2182 => 13,
    2183 => 13,
    2184 => 13,
    2185 => 13,
    2186 => 13,
    2187 => 13,
    2188 => 13,
    2189 => 13,
    2190 => 13,
    2191 => 13,
    2192 => 13,
    2193 => 13,
    2194 => 13,
    2195 => 13,
    2196 => 13,
    2197 => 13,
    2198 => 13,
    2199 => 13,
    2200 => 13,
    2201 => 13,
    2202 => 13,
    2203 => 13,
    2204 => 13,
    2205 => 13,
    2206 => 13,
    2207 => 13,
    2208 => 13,
    2209 => 13,
    2210 => 13,
    2211 => 13,
    2212 => 13,
    2213 => 13,
    2214 => 13,
    2215 => 13,
    2216 => 13,
    2217 => 13,
    2218 => 13,
    2219 => 13,
    2220 => 13,
    2221 => 13,
    2222 => 13,
    2223 => 13,
    2224 => 13,
    2225 => 13,
    2226 => 13,
    2227 => 13,
    2228 => 13,
    2229 => 13,
    2230 => 13,
    2231 => 13,
    2232 => 13,
    2233 => 13,
    2234 => 13,
    2235 => 13,
    2236 => 13,
    2237 => 13,
    2238 => 13,
    2239 => 13,
    2240 => 13,
    2241 => 13,
    2242 => 13,
    2243 => 13,
    2244 => 13,
    2245 => 13,
    2246 => 13,
    2247 => 13,
    2248 => 13,
    2249 => 13,
    2250 => 13,
    2251 => 13,
    2252 => 13,
    2253 => 14,
    2254 => 14,
    2255 => 14,
    2256 => 14,
    2257 => 14,
    2258 => 14,
    2259 => 14,
    2260 => 14,
    2261 => 14,
    2262 => 14,
    2263 => 14,
    2264 => 14,
    2265 => 14,
    2266 => 14,
    2267 => 14,
    2268 => 14,
    2269 => 14,
    2270 => 14,
    2271 => 14,
    2272 => 14,
    2273 => 14,
    2274 => 14,
    2275 => 14,
    2276 => 14,
    2277 => 14,
    2278 => 14,
    2279 => 14,
    2280 => 14,
    2281 => 14,
    2282 => 14,
    2283 => 14,
    2284 => 14,
    2285 => 14,
    2286 => 14,
    2287 => 14,
    2288 => 14,
    2289 => 14,
    2290 => 14,
    2291 => 14,
    2292 => 14,
    2293 => 14,
    2294 => 14,
    2295 => 14,
    2296 => 14,
    2297 => 14,
    2298 => 14,
    2299 => 14,
    2300 => 14,
    2301 => 14,
    2302 => 14,
    2303 => 14,
    2304 => 14,
    2305 => 14,
    2306 => 14,
    2307 => 14,
    2308 => 14,
    2309 => 14,
    2310 => 14,
    2311 => 14,
    2312 => 14,
    2313 => 14,
    2314 => 14,
    2315 => 14,
    2316 => 14,
    2317 => 14,
    2318 => 14,
    2319 => 14,
    2320 => 14,
    2321 => 14,
    2322 => 14,
    2323 => 14,
    2324 => 14,
    2325 => 14,
    2326 => 14,
    2327 => 14,
    2328 => 14,
    2329 => 14,
    2330 => 14,
    2331 => 14,
    2332 => 14,
    2333 => 14,
    2334 => 14,
    2335 => 14,
    2336 => 14,
    2337 => 14,
    2338 => 14,
    2339 => 14,
    2340 => 14,
    2341 => 14,
    2342 => 14,
    2343 => 14,
    2344 => 14,
    2345 => 14,
    2346 => 14,
    2347 => 14,
    2348 => 14,
    2349 => 14,
    2350 => 14,
    2351 => 14,
    2352 => 14,
    2353 => 14,
    2354 => 14,
    2355 => 14,
    2356 => 14,
    2357 => 14,
    2358 => 14,
    2359 => 14,
    2360 => 14,
    2361 => 14,
    2362 => 14,
    2363 => 14,
    2364 => 14,
    2365 => 14,
    2366 => 14,
    2367 => 14,
    2368 => 14,
    2369 => 14,
    2370 => 14,
    2371 => 14,
    2372 => 14,
    2373 => 14,
    2374 => 14,
    2375 => 14,
    2376 => 14,
    2377 => 14,
    2378 => 14,
    2379 => 14,
    2380 => 14,
    2381 => 14,
    2382 => 14,
    2383 => 14,
    2384 => 14,
    2385 => 14,
    2386 => 14,
    2387 => 14,
    2388 => 14,
    2389 => 14,
    2390 => 14,
    2391 => 14,
    2392 => 14,
    2393 => 14,
    2394 => 14,
    2395 => 14,
    2396 => 14,
    2397 => 14,
    2398 => 14,
    2399 => 14,
    2400 => 14,
    2401 => 14,
    2402 => 14,
    2403 => 14,
    2404 => 14,
    2405 => 14,
    2406 => 14,
    2407 => 14,
    2408 => 14,
    2409 => 14,
    2410 => 14,
    2411 => 14,
    2412 => 14,
    2413 => 14,
    2414 => 14,
    2415 => 14,
    2416 => 14,
    2417 => 14,
    2418 => 14,
    2419 => 14,
    2420 => 14,
    2421 => 14,
    2422 => 14,
    2423 => 15,
    2424 => 15,
    2425 => 15,
    2426 => 15,
    2427 => 15,
    2428 => 15,
    2429 => 15,
    2430 => 15,
    2431 => 15,
    2432 => 15,
    2433 => 15,
    2434 => 15,
    2435 => 15,
    2436 => 15,
    2437 => 15,
    2438 => 15,
    2439 => 15,
    2440 => 15,
    2441 => 15,
    2442 => 15,
    2443 => 15,
    2444 => 15,
    2445 => 15,
    2446 => 15,
    2447 => 15,
    2448 => 15,
    2449 => 15,
    2450 => 15,
    2451 => 15,
    2452 => 15,
    2453 => 15,
    2454 => 15,
    2455 => 15,
    2456 => 15,
    2457 => 15,
    2458 => 15,
    2459 => 15,
    2460 => 15,
    2461 => 15,
    2462 => 15,
    2463 => 15,
    2464 => 15,
    2465 => 15,
    2466 => 15,
    2467 => 15,
    2468 => 15,
    2469 => 15,
    2470 => 15,
    2471 => 15,
    2472 => 15,
    2473 => 15,
    2474 => 15,
    2475 => 15,
    2476 => 15,
    2477 => 15,
    2478 => 15,
    2479 => 15,
    2480 => 15,
    2481 => 15,
    2482 => 15,
    2483 => 15,
    2484 => 15,
    2485 => 15,
    2486 => 15,
    2487 => 15,
    2488 => 15,
    2489 => 15,
    2490 => 15,
    2491 => 15,
    2492 => 15,
    2493 => 15,
    2494 => 15,
    2495 => 15,
    2496 => 15,
    2497 => 15,
    2498 => 15,
    2499 => 15,
    2500 => 15,
    2501 => 15,
    2502 => 15,
    2503 => 15,
    2504 => 15,
    2505 => 15,
    2506 => 15,
    2507 => 15,
    2508 => 15,
    2509 => 15,
    2510 => 15,
    2511 => 15,
    2512 => 15,
    2513 => 15,
    2514 => 15,
    2515 => 15,
    2516 => 15,
    2517 => 15,
    2518 => 15,
    2519 => 15,
    2520 => 15,
    2521 => 15,
    2522 => 15,
    2523 => 15,
    2524 => 15,
    2525 => 15,
    2526 => 15,
    2527 => 15,
    2528 => 15,
    2529 => 15,
    2530 => 15,
    2531 => 15,
    2532 => 15,
    2533 => 15,
    2534 => 15,
    2535 => 15,
    2536 => 15,
    2537 => 15,
    2538 => 15,
    2539 => 15,
    2540 => 15,
    2541 => 15,
    2542 => 15,
    2543 => 15,
    2544 => 15,
    2545 => 15,
    2546 => 15,
    2547 => 15,
    2548 => 15,
    2549 => 15,
    2550 => 15,
    2551 => 15,
    2552 => 15,
    2553 => 15,
    2554 => 15,
    2555 => 15,
    2556 => 15,
    2557 => 15,
    2558 => 15,
    2559 => 15,
    2560 => 15,
    2561 => 15,
    2562 => 15,
    2563 => 15,
    2564 => 15,
    2565 => 15,
    2566 => 15,
    2567 => 15,
    2568 => 15,
    2569 => 15,
    2570 => 15,
    2571 => 15,
    2572 => 15,
    2573 => 15,
    2574 => 15,
    2575 => 15,
    2576 => 15,
    2577 => 15,
    2578 => 15,
    2579 => 15,
    2580 => 15,
    2581 => 15,
    2582 => 15,
    2583 => 15,
    2584 => 15,
    2585 => 15,
    2586 => 15,
    2587 => 15,
    2588 => 15,
    2589 => 15,
    2590 => 15,
    2591 => 15,
    2592 => 15,
    2593 => 16,
    2594 => 16,
    2595 => 16,
    2596 => 16,
    2597 => 16,
    2598 => 16,
    2599 => 16,
    2600 => 16,
    2601 => 16,
    2602 => 16,
    2603 => 16,
    2604 => 16,
    2605 => 16,
    2606 => 16,
    2607 => 16,
    2608 => 16,
    2609 => 16,
    2610 => 16,
    2611 => 16,
    2612 => 16,
    2613 => 16,
    2614 => 16,
    2615 => 16,
    2616 => 16,
    2617 => 16,
    2618 => 16,
    2619 => 16,
    2620 => 16,
    2621 => 16,
    2622 => 16,
    2623 => 16,
    2624 => 16,
    2625 => 16,
    2626 => 16,
    2627 => 16,
    2628 => 16,
    2629 => 16,
    2630 => 16,
    2631 => 16,
    2632 => 16,
    2633 => 16,
    2634 => 16,
    2635 => 16,
    2636 => 16,
    2637 => 16,
    2638 => 16,
    2639 => 16,
    2640 => 16,
    2641 => 16,
    2642 => 16,
    2643 => 16,
    2644 => 16,
    2645 => 16,
    2646 => 16,
    2647 => 16,
    2648 => 16,
    2649 => 16,
    2650 => 16,
    2651 => 16,
    2652 => 16,
    2653 => 16,
    2654 => 16,
    2655 => 16,
    2656 => 16,
    2657 => 16,
    2658 => 16,
    2659 => 16,
    2660 => 16,
    2661 => 16,
    2662 => 16,
    2663 => 16,
    2664 => 16,
    2665 => 16,
    2666 => 16,
    2667 => 16,
    2668 => 16,
    2669 => 16,
    2670 => 16,
    2671 => 16,
    2672 => 16,
    2673 => 16,
    2674 => 16,
    2675 => 16,
    2676 => 16,
    2677 => 16,
    2678 => 16,
    2679 => 16,
    2680 => 16,
    2681 => 16,
    2682 => 16,
    2683 => 16,
    2684 => 16,
    2685 => 16,
    2686 => 16,
    2687 => 16,
    2688 => 16,
    2689 => 16,
    2690 => 16,
    2691 => 16,
    2692 => 16,
    2693 => 16,
    2694 => 16,
    2695 => 16,
    2696 => 16,
    2697 => 16,
    2698 => 16,
    2699 => 16,
    2700 => 16,
    2701 => 16,
    2702 => 16,
    2703 => 16,
    2704 => 16,
    2705 => 16,
    2706 => 16,
    2707 => 16,
    2708 => 16,
    2709 => 16,
    2710 => 16,
    2711 => 16,
    2712 => 16,
    2713 => 16,
    2714 => 16,
    2715 => 16,
    2716 => 16,
    2717 => 16,
    2718 => 16,
    2719 => 16,
    2720 => 16,
    2721 => 16,
    2722 => 16,
    2723 => 16,
    2724 => 16,
    2725 => 16,
    2726 => 16,
    2727 => 16,
    2728 => 16,
    2729 => 16,
    2730 => 16,
    2731 => 16,
    2732 => 16,
    2733 => 16,
    2734 => 16,
    2735 => 16,
    2736 => 16,
    2737 => 16,
    2738 => 16,
    2739 => 16,
    2740 => 16,
    2741 => 16,
    2742 => 16,
    2743 => 16,
    2744 => 16,
    2745 => 16,
    2746 => 16,
    2747 => 16,
    2748 => 16,
    2749 => 16,
    2750 => 16,
    2751 => 16,
    2752 => 16,
    2753 => 16,
    2754 => 16,
    2755 => 16,
    2756 => 16,
    2757 => 16,
    2758 => 16,
    2759 => 16,
    2760 => 16,
    2761 => 16,
    2762 => 16,
    2763 => 16,
    2764 => 16,
    2765 => 17,
    2766 => 17,
    2767 => 17,
    2768 => 17,
    2769 => 17,
    2770 => 17,
    2771 => 17,
    2772 => 17,
    2773 => 17,
    2774 => 17,
    2775 => 17,
    2776 => 17,
    2777 => 17,
    2778 => 17,
    2779 => 17,
    2780 => 17,
    2781 => 17,
    2782 => 17,
    2783 => 17,
    2784 => 17,
    2785 => 17,
    2786 => 17,
    2787 => 17,
    2788 => 17,
    2789 => 17,
    2790 => 17,
    2791 => 17,
    2792 => 17,
    2793 => 17,
    2794 => 17,
    2795 => 17,
    2796 => 17,
    2797 => 17,
    2798 => 17,
    2799 => 17,
    2800 => 17,
    2801 => 17,
    2802 => 17,
    2803 => 17,
    2804 => 17,
    2805 => 17,
    2806 => 17,
    2807 => 17,
    2808 => 17,
    2809 => 17,
    2810 => 17,
    2811 => 17,
    2812 => 17,
    2813 => 17,
    2814 => 17,
    2815 => 17,
    2816 => 17,
    2817 => 17,
    2818 => 17,
    2819 => 17,
    2820 => 17,
    2821 => 17,
    2822 => 17,
    2823 => 17,
    2824 => 17,
    2825 => 17,
    2826 => 17,
    2827 => 17,
    2828 => 17,
    2829 => 17,
    2830 => 17,
    2831 => 17,
    2832 => 17,
    2833 => 17,
    2834 => 17,
    2835 => 17,
    2836 => 17,
    2837 => 17,
    2838 => 17,
    2839 => 17,
    2840 => 17,
    2841 => 17,
    2842 => 17,
    2843 => 17,
    2844 => 17,
    2845 => 17,
    2846 => 17,
    2847 => 17,
    2848 => 17,
    2849 => 17,
    2850 => 17,
    2851 => 17,
    2852 => 17,
    2853 => 17,
    2854 => 17,
    2855 => 17,
    2856 => 17,
    2857 => 17,
    2858 => 17,
    2859 => 17,
    2860 => 17,
    2861 => 17,
    2862 => 17,
    2863 => 17,
    2864 => 17,
    2865 => 17,
    2866 => 17,
    2867 => 17,
    2868 => 17,
    2869 => 17,
    2870 => 17,
    2871 => 17,
    2872 => 17,
    2873 => 17,
    2874 => 17,
    2875 => 17,
    2876 => 17,
    2877 => 17,
    2878 => 17,
    2879 => 17,
    2880 => 17,
    2881 => 17,
    2882 => 17,
    2883 => 17,
    2884 => 17,
    2885 => 17,
    2886 => 17,
    2887 => 17,
    2888 => 17,
    2889 => 17,
    2890 => 17,
    2891 => 17,
    2892 => 17,
    2893 => 17,
    2894 => 17,
    2895 => 17,
    2896 => 17,
    2897 => 17,
    2898 => 17,
    2899 => 17,
    2900 => 17,
    2901 => 17,
    2902 => 17,
    2903 => 17,
    2904 => 17,
    2905 => 17,
    2906 => 17,
    2907 => 17,
    2908 => 17,
    2909 => 17,
    2910 => 17,
    2911 => 17,
    2912 => 17,
    2913 => 17,
    2914 => 17,
    2915 => 17,
    2916 => 17,
    2917 => 17,
    2918 => 17,
    2919 => 17,
    2920 => 17,
    2921 => 17,
    2922 => 17,
    2923 => 17,
    2924 => 17,
    2925 => 17,
    2926 => 17,
    2927 => 17,
    2928 => 17,
    2929 => 17,
    2930 => 17,
    2931 => 17,
    2932 => 17,
    2933 => 17,
    2934 => 17,
    2935 => 17,
    2936 => 18,
    2937 => 18,
    2938 => 18,
    2939 => 18,
    2940 => 18,
    2941 => 18,
    2942 => 18,
    2943 => 18,
    2944 => 18,
    2945 => 18,
    2946 => 18,
    2947 => 18,
    2948 => 18,
    2949 => 18,
    2950 => 18,
    2951 => 18,
    2952 => 18,
    2953 => 18,
    2954 => 18,
    2955 => 18,
    2956 => 18,
    2957 => 18,
    2958 => 18,
    2959 => 18,
    2960 => 18,
    2961 => 18,
    2962 => 18,
    2963 => 18,
    2964 => 18,
    2965 => 18,
    2966 => 18,
    2967 => 18,
    2968 => 18,
    2969 => 18,
    2970 => 18,
    2971 => 18,
    2972 => 18,
    2973 => 18,
    2974 => 18,
    2975 => 18,
    2976 => 18,
    2977 => 18,
    2978 => 18,
    2979 => 18,
    2980 => 18,
    2981 => 18,
    2982 => 18,
    2983 => 18,
    2984 => 18,
    2985 => 18,
    2986 => 18,
    2987 => 18,
    2988 => 18,
    2989 => 18,
    2990 => 18,
    2991 => 18,
    2992 => 18,
    2993 => 18,
    2994 => 18,
    2995 => 18,
    2996 => 18,
    2997 => 18,
    2998 => 18,
    2999 => 18,
    3000 => 18,
    3001 => 18,
    3002 => 18,
    3003 => 18,
    3004 => 18,
    3005 => 18,
    3006 => 18,
    3007 => 18,
    3008 => 18,
    3009 => 18,
    3010 => 18,
    3011 => 18,
    3012 => 18,
    3013 => 18,
    3014 => 18,
    3015 => 18,
    3016 => 18,
    3017 => 18,
    3018 => 18,
    3019 => 18,
    3020 => 18,
    3021 => 18,
    3022 => 18,
    3023 => 18,
    3024 => 18,
    3025 => 18,
    3026 => 18,
    3027 => 18,
    3028 => 18,
    3029 => 18,
    3030 => 18,
    3031 => 18,
    3032 => 18,
    3033 => 18,
    3034 => 18,
    3035 => 18,
    3036 => 18,
    3037 => 18,
    3038 => 18,
    3039 => 18,
    3040 => 18,
    3041 => 18,
    3042 => 18,
    3043 => 18,
    3044 => 18,
    3045 => 18,
    3046 => 18,
    3047 => 18,
    3048 => 18,
    3049 => 18,
    3050 => 18,
    3051 => 18,
    3052 => 18,
    3053 => 18,
    3054 => 18,
    3055 => 18,
    3056 => 18,
    3057 => 18,
    3058 => 18,
    3059 => 18,
    3060 => 18,
    3061 => 18,
    3062 => 18,
    3063 => 18,
    3064 => 18,
    3065 => 18,
    3066 => 18,
    3067 => 18,
    3068 => 18,
    3069 => 18,
    3070 => 18,
    3071 => 18,
    3072 => 18,
    3073 => 18,
    3074 => 18,
    3075 => 18,
    3076 => 18,
    3077 => 18,
    3078 => 18,
    3079 => 18,
    3080 => 18,
    3081 => 18,
    3082 => 18,
    3083 => 18,
    3084 => 18,
    3085 => 18,
    3086 => 18,
    3087 => 18,
    3088 => 18,
    3089 => 18,
    3090 => 18,
    3091 => 18,
    3092 => 18,
    3093 => 18,
    3094 => 18,
    3095 => 18,
    3096 => 18,
    3097 => 18,
    3098 => 18,
    3099 => 18,
    3100 => 18,
    3101 => 18,
    3102 => 18,
    3103 => 18,
    3104 => 18,
    3105 => 18,
    3106 => 18,
    3107 => 18,
    3108 => 18,
    3109 => 19,
    3110 => 19,
    3111 => 19,
    3112 => 19,
    3113 => 19,
    3114 => 19,
    3115 => 19,
    3116 => 19,
    3117 => 19,
    3118 => 19,
    3119 => 19,
    3120 => 19,
    3121 => 19,
    3122 => 19,
    3123 => 19,
    3124 => 19,
    3125 => 19,
    3126 => 19,
    3127 => 19,
    3128 => 19,
    3129 => 19,
    3130 => 19,
    3131 => 19,
    3132 => 19,
    3133 => 19,
    3134 => 19,
    3135 => 19,
    3136 => 19,
    3137 => 19,
    3138 => 19,
    3139 => 19,
    3140 => 19,
    3141 => 19,
    3142 => 19,
    3143 => 19,
    3144 => 19,
    3145 => 19,
    3146 => 19,
    3147 => 19,
    3148 => 19,
    3149 => 19,
    3150 => 19,
    3151 => 19,
    3152 => 19,
    3153 => 19,
    3154 => 19,
    3155 => 19,
    3156 => 19,
    3157 => 19,
    3158 => 19,
    3159 => 19,
    3160 => 19,
    3161 => 19,
    3162 => 19,
    3163 => 19,
    3164 => 19,
    3165 => 19,
    3166 => 19,
    3167 => 19,
    3168 => 19,
    3169 => 19,
    3170 => 19,
    3171 => 19,
    3172 => 19,
    3173 => 19,
    3174 => 19,
    3175 => 19,
    3176 => 19,
    3177 => 19,
    3178 => 19,
    3179 => 19,
    3180 => 19,
    3181 => 19,
    3182 => 19,
    3183 => 19,
    3184 => 19,
    3185 => 19,
    3186 => 19,
    3187 => 19,
    3188 => 19,
    3189 => 19,
    3190 => 19,
    3191 => 19,
    3192 => 19,
    3193 => 19,
    3194 => 19,
    3195 => 19,
    3196 => 19,
    3197 => 19,
    3198 => 19,
    3199 => 19,
    3200 => 19,
    3201 => 19,
    3202 => 19,
    3203 => 19,
    3204 => 19,
    3205 => 19,
    3206 => 19,
    3207 => 19,
    3208 => 19,
    3209 => 19,
    3210 => 19,
    3211 => 19,
    3212 => 19,
    3213 => 19,
    3214 => 19,
    3215 => 19,
    3216 => 19,
    3217 => 19,
    3218 => 19,
    3219 => 19,
    3220 => 19,
    3221 => 19,
    3222 => 19,
    3223 => 19,
    3224 => 19,
    3225 => 19,
    3226 => 19,
    3227 => 19,
    3228 => 19,
    3229 => 19,
    3230 => 19,
    3231 => 19,
    3232 => 19,
    3233 => 19,
    3234 => 19,
    3235 => 19,
    3236 => 19,
    3237 => 19,
    3238 => 19,
    3239 => 19,
    3240 => 19,
    3241 => 19,
    3242 => 19,
    3243 => 19,
    3244 => 19,
    3245 => 19,
    3246 => 19,
    3247 => 19,
    3248 => 19,
    3249 => 19,
    3250 => 19,
    3251 => 19,
    3252 => 19,
    3253 => 19,
    3254 => 19,
    3255 => 19,
    3256 => 19,
    3257 => 19,
    3258 => 19,
    3259 => 19,
    3260 => 19,
    3261 => 19,
    3262 => 19,
    3263 => 19,
    3264 => 19,
    3265 => 19,
    3266 => 19,
    3267 => 19,
    3268 => 19,
    3269 => 19,
    3270 => 19,
    3271 => 19,
    3272 => 19,
    3273 => 19,
    3274 => 19,
    3275 => 19,
    3276 => 19,
    3277 => 19,
    3278 => 19,
    3279 => 19,
    3280 => 19,
    3281 => 19,
    3282 => 19,
    3283 => 20,
    3284 => 20,
    3285 => 20,
    3286 => 20,
    3287 => 20,
    3288 => 20,
    3289 => 20,
    3290 => 20,
    3291 => 20,
    3292 => 20,
    3293 => 20,
    3294 => 20,
    3295 => 20,
    3296 => 20,
    3297 => 20,
    3298 => 20,
    3299 => 20,
    3300 => 20,
    3301 => 20,
    3302 => 20,
    3303 => 20,
    3304 => 20,
    3305 => 20,
    3306 => 20,
    3307 => 20,
    3308 => 20,
    3309 => 20,
    3310 => 20,
    3311 => 20,
    3312 => 20,
    3313 => 20,
    3314 => 20,
    3315 => 20,
    3316 => 20,
    3317 => 20,
    3318 => 20,
    3319 => 20,
    3320 => 20,
    3321 => 20,
    3322 => 20,
    3323 => 20,
    3324 => 20,
    3325 => 20,
    3326 => 20,
    3327 => 20,
    3328 => 20,
    3329 => 20,
    3330 => 20,
    3331 => 20,
    3332 => 20,
    3333 => 20,
    3334 => 20,
    3335 => 20,
    3336 => 20,
    3337 => 20,
    3338 => 20,
    3339 => 20,
    3340 => 20,
    3341 => 20,
    3342 => 20,
    3343 => 20,
    3344 => 20,
    3345 => 20,
    3346 => 20,
    3347 => 20,
    3348 => 20,
    3349 => 20,
    3350 => 20,
    3351 => 20,
    3352 => 20,
    3353 => 20,
    3354 => 20,
    3355 => 20,
    3356 => 20,
    3357 => 20,
    3358 => 20,
    3359 => 20,
    3360 => 20,
    3361 => 20,
    3362 => 20,
    3363 => 20,
    3364 => 20,
    3365 => 20,
    3366 => 20,
    3367 => 20,
    3368 => 20,
    3369 => 20,
    3370 => 20,
    3371 => 20,
    3372 => 20,
    3373 => 20,
    3374 => 20,
    3375 => 20,
    3376 => 20,
    3377 => 20,
    3378 => 20,
    3379 => 20,
    3380 => 20,
    3381 => 20,
    3382 => 20,
    3383 => 20,
    3384 => 20,
    3385 => 20,
    3386 => 20,
    3387 => 20,
    3388 => 20,
    3389 => 20,
    3390 => 20,
    3391 => 20,
    3392 => 20,
    3393 => 20,
    3394 => 20,
    3395 => 20,
    3396 => 20,
    3397 => 20,
    3398 => 20,
    3399 => 20,
    3400 => 20,
    3401 => 20,
    3402 => 20,
    3403 => 20,
    3404 => 20,
    3405 => 20,
    3406 => 20,
    3407 => 20,
    3408 => 20,
    3409 => 20,
    3410 => 20,
    3411 => 20,
    3412 => 20,
    3413 => 20,
    3414 => 20,
    3415 => 20,
    3416 => 20,
    3417 => 20,
    3418 => 20,
    3419 => 20,
    3420 => 20,
    3421 => 20,
    3422 => 20,
    3423 => 20,
    3424 => 20,
    3425 => 20,
    3426 => 20,
    3427 => 20,
    3428 => 20,
    3429 => 20,
    3430 => 20,
    3431 => 20,
    3432 => 20,
    3433 => 20,
    3434 => 20,
    3435 => 20,
    3436 => 20,
    3437 => 20,
    3438 => 20,
    3439 => 20,
    3440 => 20,
    3441 => 20,
    3442 => 20,
    3443 => 20,
    3444 => 20,
    3445 => 20,
    3446 => 20,
    3447 => 20,
    3448 => 20,
    3449 => 20,
    3450 => 20,
    3451 => 20,
    3452 => 20,
    3453 => 20,
    3454 => 20,
    3455 => 20,
    3456 => 20,
    3457 => 21,
    3458 => 21,
    3459 => 21,
    3460 => 21,
    3461 => 21,
    3462 => 21,
    3463 => 21,
    3464 => 21,
    3465 => 21,
    3466 => 21,
    3467 => 21,
    3468 => 21,
    3469 => 21,
    3470 => 21,
    3471 => 21,
    3472 => 21,
    3473 => 21,
    3474 => 21,
    3475 => 21,
    3476 => 21,
    3477 => 21,
    3478 => 21,
    3479 => 21,
    3480 => 21,
    3481 => 21,
    3482 => 21,
    3483 => 21,
    3484 => 21,
    3485 => 21,
    3486 => 21,
    3487 => 21,
    3488 => 21,
    3489 => 21,
    3490 => 21,
    3491 => 21,
    3492 => 21,
    3493 => 21,
    3494 => 21,
    3495 => 21,
    3496 => 21,
    3497 => 21,
    3498 => 21,
    3499 => 21,
    3500 => 21,
    3501 => 21,
    3502 => 21,
    3503 => 21,
    3504 => 21,
    3505 => 21,
    3506 => 21,
    3507 => 21,
    3508 => 21,
    3509 => 21,
    3510 => 21,
    3511 => 21,
    3512 => 21,
    3513 => 21,
    3514 => 21,
    3515 => 21,
    3516 => 21,
    3517 => 21,
    3518 => 21,
    3519 => 21,
    3520 => 21,
    3521 => 21,
    3522 => 21,
    3523 => 21,
    3524 => 21,
    3525 => 21,
    3526 => 21,
    3527 => 21,
    3528 => 21,
    3529 => 21,
    3530 => 21,
    3531 => 21,
    3532 => 21,
    3533 => 21,
    3534 => 21,
    3535 => 21,
    3536 => 21,
    3537 => 21,
    3538 => 21,
    3539 => 21,
    3540 => 21,
    3541 => 21,
    3542 => 21,
    3543 => 21,
    3544 => 21,
    3545 => 21,
    3546 => 21,
    3547 => 21,
    3548 => 21,
    3549 => 21,
    3550 => 21,
    3551 => 21,
    3552 => 21,
    3553 => 21,
    3554 => 21,
    3555 => 21,
    3556 => 21,
    3557 => 21,
    3558 => 21,
    3559 => 21,
    3560 => 21,
    3561 => 21,
    3562 => 21,
    3563 => 21,
    3564 => 21,
    3565 => 21,
    3566 => 21,
    3567 => 21,
    3568 => 21,
    3569 => 21,
    3570 => 21,
    3571 => 21,
    3572 => 21,
    3573 => 21,
    3574 => 21,
    3575 => 21,
    3576 => 21,
    3577 => 21,
    3578 => 21,
    3579 => 21,
    3580 => 21,
    3581 => 21,
    3582 => 21,
    3583 => 21,
    3584 => 21,
    3585 => 21,
    3586 => 21,
    3587 => 21,
    3588 => 21,
    3589 => 21,
    3590 => 21,
    3591 => 21,
    3592 => 21,
    3593 => 21,
    3594 => 21,
    3595 => 21,
    3596 => 21,
    3597 => 21,
    3598 => 21,
    3599 => 21,
    3600 => 21,
    3601 => 21,
    3602 => 21,
    3603 => 21,
    3604 => 21,
    3605 => 21,
    3606 => 21,
    3607 => 21,
    3608 => 21,
    3609 => 21,
    3610 => 21,
    3611 => 21,
    3612 => 21,
    3613 => 21,
    3614 => 21,
    3615 => 21,
    3616 => 21,
    3617 => 21,
    3618 => 21,
    3619 => 21,
    3620 => 21,
    3621 => 21,
    3622 => 21,
    3623 => 21,
    3624 => 21,
    3625 => 21,
    3626 => 21,
    3627 => 21,
    3628 => 21,
    3629 => 21,
    3630 => 21,
    3631 => 21,
    3632 => 21,
    3633 => 22,
    3634 => 22,
    3635 => 22,
    3636 => 22,
    3637 => 22,
    3638 => 22,
    3639 => 22,
    3640 => 22,
    3641 => 22,
    3642 => 22,
    3643 => 22,
    3644 => 22,
    3645 => 22,
    3646 => 22,
    3647 => 22,
    3648 => 22,
    3649 => 22,
    3650 => 22,
    3651 => 22,
    3652 => 22,
    3653 => 22,
    3654 => 22,
    3655 => 22,
    3656 => 22,
    3657 => 22,
    3658 => 22,
    3659 => 22,
    3660 => 22,
    3661 => 22,
    3662 => 22,
    3663 => 22,
    3664 => 22,
    3665 => 22,
    3666 => 22,
    3667 => 22,
    3668 => 22,
    3669 => 22,
    3670 => 22,
    3671 => 22,
    3672 => 22,
    3673 => 22,
    3674 => 22,
    3675 => 22,
    3676 => 22,
    3677 => 22,
    3678 => 22,
    3679 => 22,
    3680 => 22,
    3681 => 22,
    3682 => 22,
    3683 => 22,
    3684 => 22,
    3685 => 22,
    3686 => 22,
    3687 => 22,
    3688 => 22,
    3689 => 22,
    3690 => 22,
    3691 => 22,
    3692 => 22,
    3693 => 22,
    3694 => 22,
    3695 => 22,
    3696 => 22,
    3697 => 22,
    3698 => 22,
    3699 => 22,
    3700 => 22,
    3701 => 22,
    3702 => 22,
    3703 => 22,
    3704 => 22,
    3705 => 22,
    3706 => 22,
    3707 => 22,
    3708 => 22,
    3709 => 22,
    3710 => 22,
    3711 => 22,
    3712 => 22,
    3713 => 22,
    3714 => 22,
    3715 => 22,
    3716 => 22,
    3717 => 22,
    3718 => 22,
    3719 => 22,
    3720 => 22,
    3721 => 22,
    3722 => 22,
    3723 => 22,
    3724 => 22,
    3725 => 22,
    3726 => 22,
    3727 => 22,
    3728 => 22,
    3729 => 22,
    3730 => 22,
    3731 => 22,
    3732 => 22,
    3733 => 22,
    3734 => 22,
    3735 => 22,
    3736 => 22,
    3737 => 22,
    3738 => 22,
    3739 => 22,
    3740 => 22,
    3741 => 22,
    3742 => 22,
    3743 => 22,
    3744 => 22,
    3745 => 22,
    3746 => 22,
    3747 => 22,
    3748 => 22,
    3749 => 22,
    3750 => 22,
    3751 => 22,
    3752 => 22,
    3753 => 22,
    3754 => 22,
    3755 => 22,
    3756 => 22,
    3757 => 22,
    3758 => 22,
    3759 => 22,
    3760 => 22,
    3761 => 22,
    3762 => 22,
    3763 => 22,
    3764 => 22,
    3765 => 22,
    3766 => 22,
    3767 => 22,
    3768 => 22,
    3769 => 22,
    3770 => 22,
    3771 => 22,
    3772 => 22,
    3773 => 22,
    3774 => 22,
    3775 => 22,
    3776 => 22,
    3777 => 22,
    3778 => 22,
    3779 => 22,
    3780 => 22,
    3781 => 22,
    3782 => 22,
    3783 => 22,
    3784 => 22,
    3785 => 22,
    3786 => 22,
    3787 => 22,
    3788 => 22,
    3789 => 22,
    3790 => 22,
    3791 => 22,
    3792 => 22,
    3793 => 22,
    3794 => 22,
    3795 => 22,
    3796 => 22,
    3797 => 22,
    3798 => 22,
    3799 => 22,
    3800 => 22,
    3801 => 22,
    3802 => 22,
    3803 => 22,
    3804 => 22,
    3805 => 22,
    3806 => 22,
    3807 => 22,
    3808 => 22,
    3809 => 22,
    3810 => 23,
    3811 => 23,
    3812 => 23,
    3813 => 23,
    3814 => 23,
    3815 => 23,
    3816 => 23,
    3817 => 23,
    3818 => 23,
    3819 => 23,
    3820 => 23,
    3821 => 23,
    3822 => 23,
    3823 => 23,
    3824 => 23,
    3825 => 23,
    3826 => 23,
    3827 => 23,
    3828 => 23,
    3829 => 23,
    3830 => 23,
    3831 => 23,
    3832 => 23,
    3833 => 23,
    3834 => 23,
    3835 => 23,
    3836 => 23,
    3837 => 23,
    3838 => 23,
    3839 => 23,
    3840 => 23,
    3841 => 23,
    3842 => 23,
    3843 => 23,
    3844 => 23,
    3845 => 23,
    3846 => 23,
    3847 => 23,
    3848 => 23,
    3849 => 23,
    3850 => 23,
    3851 => 23,
    3852 => 23,
    3853 => 23,
    3854 => 23,
    3855 => 23,
    3856 => 23,
    3857 => 23,
    3858 => 23,
    3859 => 23,
    3860 => 23,
    3861 => 23,
    3862 => 23,
    3863 => 23,
    3864 => 23,
    3865 => 23,
    3866 => 23,
    3867 => 23,
    3868 => 23,
    3869 => 23,
    3870 => 23,
    3871 => 23,
    3872 => 23,
    3873 => 23,
    3874 => 23,
    3875 => 23,
    3876 => 23,
    3877 => 23,
    3878 => 23,
    3879 => 23,
    3880 => 23,
    3881 => 23,
    3882 => 23,
    3883 => 23,
    3884 => 23,
    3885 => 23,
    3886 => 23,
    3887 => 23,
    3888 => 23,
    3889 => 23,
    3890 => 23,
    3891 => 23,
    3892 => 23,
    3893 => 23,
    3894 => 23,
    3895 => 23,
    3896 => 23,
    3897 => 23,
    3898 => 23,
    3899 => 23,
    3900 => 23,
    3901 => 23,
    3902 => 23,
    3903 => 23,
    3904 => 23,
    3905 => 23,
    3906 => 23,
    3907 => 23,
    3908 => 23,
    3909 => 23,
    3910 => 23,
    3911 => 23,
    3912 => 23,
    3913 => 23,
    3914 => 23,
    3915 => 23,
    3916 => 23,
    3917 => 23,
    3918 => 23,
    3919 => 23,
    3920 => 23,
    3921 => 23,
    3922 => 23,
    3923 => 23,
    3924 => 23,
    3925 => 23,
    3926 => 23,
    3927 => 23,
    3928 => 23,
    3929 => 23,
    3930 => 23,
    3931 => 23,
    3932 => 23,
    3933 => 23,
    3934 => 23,
    3935 => 23,
    3936 => 23,
    3937 => 23,
    3938 => 23,
    3939 => 23,
    3940 => 23,
    3941 => 23,
    3942 => 23,
    3943 => 23,
    3944 => 23,
    3945 => 23,
    3946 => 23,
    3947 => 23,
    3948 => 23,
    3949 => 23,
    3950 => 23,
    3951 => 23,
    3952 => 23,
    3953 => 23,
    3954 => 23,
    3955 => 23,
    3956 => 23,
    3957 => 23,
    3958 => 23,
    3959 => 23,
    3960 => 23,
    3961 => 23,
    3962 => 23,
    3963 => 23,
    3964 => 23,
    3965 => 23,
    3966 => 23,
    3967 => 23,
    3968 => 23,
    3969 => 23,
    3970 => 23,
    3971 => 23,
    3972 => 23,
    3973 => 23,
    3974 => 23,
    3975 => 23,
    3976 => 23,
    3977 => 23,
    3978 => 23,
    3979 => 23,
    3980 => 23,
    3981 => 23,
    3982 => 23,
    3983 => 23,
    3984 => 23,
    3985 => 23,
    3986 => 23,
    3987 => 23,
    3988 => 24,
    3989 => 24,
    3990 => 24,
    3991 => 24,
    3992 => 24,
    3993 => 24,
    3994 => 24,
    3995 => 24,
    3996 => 24,
    3997 => 24,
    3998 => 24,
    3999 => 24,
    4000 => 24,
    4001 => 24,
    4002 => 24,
    4003 => 24,
    4004 => 24,
    4005 => 24,
    4006 => 24,
    4007 => 24,
    4008 => 24,
    4009 => 24,
    4010 => 24,
    4011 => 24,
    4012 => 24,
    4013 => 24,
    4014 => 24,
    4015 => 24,
    4016 => 24,
    4017 => 24,
    4018 => 24,
    4019 => 24,
    4020 => 24,
    4021 => 24,
    4022 => 24,
    4023 => 24,
    4024 => 24,
    4025 => 24,
    4026 => 24,
    4027 => 24,
    4028 => 24,
    4029 => 24,
    4030 => 24,
    4031 => 24,
    4032 => 24,
    4033 => 24,
    4034 => 24,
    4035 => 24,
    4036 => 24,
    4037 => 24,
    4038 => 24,
    4039 => 24,
    4040 => 24,
    4041 => 24,
    4042 => 24,
    4043 => 24,
    4044 => 24,
    4045 => 24,
    4046 => 24,
    4047 => 24,
    4048 => 24,
    4049 => 24,
    4050 => 24,
    4051 => 24,
    4052 => 24,
    4053 => 24,
    4054 => 24,
    4055 => 24,
    4056 => 24,
    4057 => 24,
    4058 => 24,
    4059 => 24,
    4060 => 24,
    4061 => 24,
    4062 => 24,
    4063 => 24,
    4064 => 24,
    4065 => 24,
    4066 => 24,
    4067 => 24,
    4068 => 24,
    4069 => 24,
    4070 => 24,
    4071 => 24,
    4072 => 24,
    4073 => 24,
    4074 => 24,
    4075 => 24,
    4076 => 24,
    4077 => 24,
    4078 => 24,
    4079 => 24,
    4080 => 24,
    4081 => 24,
    4082 => 24,
    4083 => 24,
    4084 => 24,
    4085 => 24,
    4086 => 24,
    4087 => 24,
    4088 => 24,
    4089 => 24,
    4090 => 24,
    4091 => 24,
    4092 => 24,
    4093 => 24,
    4094 => 24,
    4095 => 24,
    4096 => 24,
    4097 => 24,
    4098 => 24,
    4099 => 24,
    4100 => 24,
    4101 => 24,
    4102 => 24,
    4103 => 24,
    4104 => 24,
    4105 => 24,
    4106 => 24,
    4107 => 24,
    4108 => 24,
    4109 => 24,
    4110 => 24,
    4111 => 24,
    4112 => 24,
    4113 => 24,
    4114 => 24,
    4115 => 24,
    4116 => 24,
    4117 => 24,
    4118 => 24,
    4119 => 24,
    4120 => 24,
    4121 => 24,
    4122 => 24,
    4123 => 24,
    4124 => 24,
    4125 => 24,
    4126 => 24,
    4127 => 24,
    4128 => 24,
    4129 => 24,
    4130 => 24,
    4131 => 24,
    4132 => 24,
    4133 => 24,
    4134 => 24,
    4135 => 24,
    4136 => 24,
    4137 => 24,
    4138 => 24,
    4139 => 24,
    4140 => 24,
    4141 => 24,
    4142 => 24,
    4143 => 24,
    4144 => 24,
    4145 => 24,
    4146 => 24,
    4147 => 24,
    4148 => 24,
    4149 => 24,
    4150 => 24,
    4151 => 24,
    4152 => 24,
    4153 => 24,
    4154 => 24,
    4155 => 24,
    4156 => 24,
    4157 => 24,
    4158 => 24,
    4159 => 24,
    4160 => 24,
    4161 => 24,
    4162 => 24,
    4163 => 24,
    4164 => 24,
    4165 => 24,
    4166 => 24,
    4167 => 25,
    4168 => 25,
    4169 => 25,
    4170 => 25,
    4171 => 25,
    4172 => 25,
    4173 => 25,
    4174 => 25,
    4175 => 25,
    4176 => 25,
    4177 => 25,
    4178 => 25,
    4179 => 25,
    4180 => 25,
    4181 => 25,
    4182 => 25,
    4183 => 25,
    4184 => 25,
    4185 => 25,
    4186 => 25,
    4187 => 25,
    4188 => 25,
    4189 => 25,
    4190 => 25,
    4191 => 25,
    4192 => 25,
    4193 => 25,
    4194 => 25,
    4195 => 25,
    4196 => 25,
    4197 => 25,
    4198 => 25,
    4199 => 25,
    4200 => 25,
    4201 => 25,
    4202 => 25,
    4203 => 25,
    4204 => 25,
    4205 => 25,
    4206 => 25,
    4207 => 25,
    4208 => 25,
    4209 => 25,
    4210 => 25,
    4211 => 25,
    4212 => 25,
    4213 => 25,
    4214 => 25,
    4215 => 25,
    4216 => 25,
    4217 => 25,
    4218 => 25,
    4219 => 25,
    4220 => 25,
    4221 => 25,
    4222 => 25,
    4223 => 25,
    4224 => 25,
    4225 => 25,
    4226 => 25,
    4227 => 25,
    4228 => 25,
    4229 => 25,
    4230 => 25,
    4231 => 25,
    4232 => 25,
    4233 => 25,
    4234 => 25,
    4235 => 25,
    4236 => 25,
    4237 => 25,
    4238 => 25,
    4239 => 25,
    4240 => 25,
    4241 => 25,
    4242 => 25,
    4243 => 25,
    4244 => 25,
    4245 => 25,
    4246 => 25,
    4247 => 25,
    4248 => 25,
    4249 => 25,
    4250 => 25,
    4251 => 25,
    4252 => 25,
    4253 => 25,
    4254 => 25,
    4255 => 25,
    4256 => 25,
    4257 => 25,
    4258 => 25,
    4259 => 25,
    4260 => 25,
    4261 => 25,
    4262 => 25,
    4263 => 25,
    4264 => 25,
    4265 => 25,
    4266 => 25,
    4267 => 25,
    4268 => 25,
    4269 => 25,
    4270 => 25,
    4271 => 25,
    4272 => 25,
    4273 => 25,
    4274 => 25,
    4275 => 25,
    4276 => 25,
    4277 => 25,
    4278 => 25,
    4279 => 25,
    4280 => 25,
    4281 => 25,
    4282 => 25,
    4283 => 25,
    4284 => 25,
    4285 => 25,
    4286 => 25,
    4287 => 25,
    4288 => 25,
    4289 => 25,
    4290 => 25,
    4291 => 25,
    4292 => 25,
    4293 => 25,
    4294 => 25,
    4295 => 25,
    4296 => 25,
    4297 => 25,
    4298 => 25,
    4299 => 25,
    4300 => 25,
    4301 => 25,
    4302 => 25,
    4303 => 25,
    4304 => 25,
    4305 => 25,
    4306 => 25,
    4307 => 25,
    4308 => 25,
    4309 => 25,
    4310 => 25,
    4311 => 25,
    4312 => 25,
    4313 => 25,
    4314 => 25,
    4315 => 25,
    4316 => 25,
    4317 => 25,
    4318 => 25,
    4319 => 25,
    4320 => 25,
    4321 => 25,
    4322 => 25,
    4323 => 25,
    4324 => 25,
    4325 => 25,
    4326 => 25,
    4327 => 25,
    4328 => 25,
    4329 => 25,
    4330 => 25,
    4331 => 25,
    4332 => 25,
    4333 => 25,
    4334 => 25,
    4335 => 25,
    4336 => 25,
    4337 => 25,
    4338 => 25,
    4339 => 25,
    4340 => 25,
    4341 => 25,
    4342 => 25,
    4343 => 25,
    4344 => 25,
    4345 => 25,
    4346 => 25,
    4347 => 26,
    4348 => 26,
    4349 => 26,
    4350 => 26,
    4351 => 26,
    4352 => 26,
    4353 => 26,
    4354 => 26,
    4355 => 26,
    4356 => 26,
    4357 => 26,
    4358 => 26,
    4359 => 26,
    4360 => 26,
    4361 => 26,
    4362 => 26,
    4363 => 26,
    4364 => 26,
    4365 => 26,
    4366 => 26,
    4367 => 26,
    4368 => 26,
    4369 => 26,
    4370 => 26,
    4371 => 26,
    4372 => 26,
    4373 => 26,
    4374 => 26,
    4375 => 26,
    4376 => 26,
    4377 => 26,
    4378 => 26,
    4379 => 26,
    4380 => 26,
    4381 => 26,
    4382 => 26,
    4383 => 26,
    4384 => 26,
    4385 => 26,
    4386 => 26,
    4387 => 26,
    4388 => 26,
    4389 => 26,
    4390 => 26,
    4391 => 26,
    4392 => 26,
    4393 => 26,
    4394 => 26,
    4395 => 26,
    4396 => 26,
    4397 => 26,
    4398 => 26,
    4399 => 26,
    4400 => 26,
    4401 => 26,
    4402 => 26,
    4403 => 26,
    4404 => 26,
    4405 => 26,
    4406 => 26,
    4407 => 26,
    4408 => 26,
    4409 => 26,
    4410 => 26,
    4411 => 26,
    4412 => 26,
    4413 => 26,
    4414 => 26,
    4415 => 26,
    4416 => 26,
    4417 => 26,
    4418 => 26,
    4419 => 26,
    4420 => 26,
    4421 => 26,
    4422 => 26,
    4423 => 26,
    4424 => 26,
    4425 => 26,
    4426 => 26,
    4427 => 26,
    4428 => 26,
    4429 => 26,
    4430 => 26,
    4431 => 26,
    4432 => 26,
    4433 => 26,
    4434 => 26,
    4435 => 26,
    4436 => 26,
    4437 => 26,
    4438 => 26,
    4439 => 26,
    4440 => 26,
    4441 => 26,
    4442 => 26,
    4443 => 26,
    4444 => 26,
    4445 => 26,
    4446 => 26,
    4447 => 26,
    4448 => 26,
    4449 => 26,
    4450 => 26,
    4451 => 26,
    4452 => 26,
    4453 => 26,
    4454 => 26,
    4455 => 26,
    4456 => 26,
    4457 => 26,
    4458 => 26,
    4459 => 26,
    4460 => 26,
    4461 => 26,
    4462 => 26,
    4463 => 26,
    4464 => 26,
    4465 => 26,
    4466 => 26,
    4467 => 26,
    4468 => 26,
    4469 => 26,
    4470 => 26,
    4471 => 26,
    4472 => 26,
    4473 => 26,
    4474 => 26,
    4475 => 26,
    4476 => 26,
    4477 => 26,
    4478 => 26,
    4479 => 26,
    4480 => 26,
    4481 => 26,
    4482 => 26,
    4483 => 26,
    4484 => 26,
    4485 => 26,
    4486 => 26,
    4487 => 26,
    4488 => 26,
    4489 => 26,
    4490 => 26,
    4491 => 26,
    4492 => 26,
    4493 => 26,
    4494 => 26,
    4495 => 26,
    4496 => 26,
    4497 => 26,
    4498 => 26,
    4499 => 26,
    4500 => 26,
    4501 => 26,
    4502 => 26,
    4503 => 26,
    4504 => 26,
    4505 => 26,
    4506 => 26,
    4507 => 26,
    4508 => 26,
    4509 => 26,
    4510 => 26,
    4511 => 26,
    4512 => 26,
    4513 => 26,
    4514 => 26,
    4515 => 26,
    4516 => 26,
    4517 => 26,
    4518 => 26,
    4519 => 26,
    4520 => 26,
    4521 => 26,
    4522 => 26,
    4523 => 26,
    4524 => 26,
    4525 => 26,
    4526 => 26,
    4527 => 26,
    4528 => 26,
    4529 => 27,
    4530 => 27,
    4531 => 27,
    4532 => 27,
    4533 => 27,
    4534 => 27,
    4535 => 27,
    4536 => 27,
    4537 => 27,
    4538 => 27,
    4539 => 27,
    4540 => 27,
    4541 => 27,
    4542 => 27,
    4543 => 27,
    4544 => 27,
    4545 => 27,
    4546 => 27,
    4547 => 27,
    4548 => 27,
    4549 => 27,
    4550 => 27,
    4551 => 27,
    4552 => 27,
    4553 => 27,
    4554 => 27,
    4555 => 27,
    4556 => 27,
    4557 => 27,
    4558 => 27,
    4559 => 27,
    4560 => 27,
    4561 => 27,
    4562 => 27,
    4563 => 27,
    4564 => 27,
    4565 => 27,
    4566 => 27,
    4567 => 27,
    4568 => 27,
    4569 => 27,
    4570 => 27,
    4571 => 27,
    4572 => 27,
    4573 => 27,
    4574 => 27,
    4575 => 27,
    4576 => 27,
    4577 => 27,
    4578 => 27,
    4579 => 27,
    4580 => 27,
    4581 => 27,
    4582 => 27,
    4583 => 27,
    4584 => 27,
    4585 => 27,
    4586 => 27,
    4587 => 27,
    4588 => 27,
    4589 => 27,
    4590 => 27,
    4591 => 27,
    4592 => 27,
    4593 => 27,
    4594 => 27,
    4595 => 27,
    4596 => 27,
    4597 => 27,
    4598 => 27,
    4599 => 27,
    4600 => 27,
    4601 => 27,
    4602 => 27,
    4603 => 27,
    4604 => 27,
    4605 => 27,
    4606 => 27,
    4607 => 27,
    4608 => 27,
    4609 => 27,
    4610 => 27,
    4611 => 27,
    4612 => 27,
    4613 => 27,
    4614 => 27,
    4615 => 27,
    4616 => 27,
    4617 => 27,
    4618 => 27,
    4619 => 27,
    4620 => 27,
    4621 => 27,
    4622 => 27,
    4623 => 27,
    4624 => 27,
    4625 => 27,
    4626 => 27,
    4627 => 27,
    4628 => 27,
    4629 => 27,
    4630 => 27,
    4631 => 27,
    4632 => 27,
    4633 => 27,
    4634 => 27,
    4635 => 27,
    4636 => 27,
    4637 => 27,
    4638 => 27,
    4639 => 27,
    4640 => 27,
    4641 => 27,
    4642 => 27,
    4643 => 27,
    4644 => 27,
    4645 => 27,
    4646 => 27,
    4647 => 27,
    4648 => 27,
    4649 => 27,
    4650 => 27,
    4651 => 27,
    4652 => 27,
    4653 => 27,
    4654 => 27,
    4655 => 27,
    4656 => 27,
    4657 => 27,
    4658 => 27,
    4659 => 27,
    4660 => 27,
    4661 => 27,
    4662 => 27,
    4663 => 27,
    4664 => 27,
    4665 => 27,
    4666 => 27,
    4667 => 27,
    4668 => 27,
    4669 => 27,
    4670 => 27,
    4671 => 27,
    4672 => 27,
    4673 => 27,
    4674 => 27,
    4675 => 27,
    4676 => 27,
    4677 => 27,
    4678 => 27,
    4679 => 27,
    4680 => 27,
    4681 => 27,
    4682 => 27,
    4683 => 27,
    4684 => 27,
    4685 => 27,
    4686 => 27,
    4687 => 27,
    4688 => 27,
    4689 => 27,
    4690 => 27,
    4691 => 27,
    4692 => 27,
    4693 => 27,
    4694 => 27,
    4695 => 27,
    4696 => 27,
    4697 => 27,
    4698 => 27,
    4699 => 27,
    4700 => 27,
    4701 => 27,
    4702 => 27,
    4703 => 27,
    4704 => 27,
    4705 => 27,
    4706 => 27,
    4707 => 27,
    4708 => 27,
    4709 => 27,
    4710 => 27,
    4711 => 27,
    4712 => 28,
    4713 => 28,
    4714 => 28,
    4715 => 28,
    4716 => 28,
    4717 => 28,
    4718 => 28,
    4719 => 28,
    4720 => 28,
    4721 => 28,
    4722 => 28,
    4723 => 28,
    4724 => 28,
    4725 => 28,
    4726 => 28,
    4727 => 28,
    4728 => 28,
    4729 => 28,
    4730 => 28,
    4731 => 28,
    4732 => 28,
    4733 => 28,
    4734 => 28,
    4735 => 28,
    4736 => 28,
    4737 => 28,
    4738 => 28,
    4739 => 28,
    4740 => 28,
    4741 => 28,
    4742 => 28,
    4743 => 28,
    4744 => 28,
    4745 => 28,
    4746 => 28,
    4747 => 28,
    4748 => 28,
    4749 => 28,
    4750 => 28,
    4751 => 28,
    4752 => 28,
    4753 => 28,
    4754 => 28,
    4755 => 28,
    4756 => 28,
    4757 => 28,
    4758 => 28,
    4759 => 28,
    4760 => 28,
    4761 => 28,
    4762 => 28,
    4763 => 28,
    4764 => 28,
    4765 => 28,
    4766 => 28,
    4767 => 28,
    4768 => 28,
    4769 => 28,
    4770 => 28,
    4771 => 28,
    4772 => 28,
    4773 => 28,
    4774 => 28,
    4775 => 28,
    4776 => 28,
    4777 => 28,
    4778 => 28,
    4779 => 28,
    4780 => 28,
    4781 => 28,
    4782 => 28,
    4783 => 28,
    4784 => 28,
    4785 => 28,
    4786 => 28,
    4787 => 28,
    4788 => 28,
    4789 => 28,
    4790 => 28,
    4791 => 28,
    4792 => 28,
    4793 => 28,
    4794 => 28,
    4795 => 28,
    4796 => 28,
    4797 => 28,
    4798 => 28,
    4799 => 28,
    4800 => 28,
    4801 => 28,
    4802 => 28,
    4803 => 28,
    4804 => 28,
    4805 => 28,
    4806 => 28,
    4807 => 28,
    4808 => 28,
    4809 => 28,
    4810 => 28,
    4811 => 28,
    4812 => 28,
    4813 => 28,
    4814 => 28,
    4815 => 28,
    4816 => 28,
    4817 => 28,
    4818 => 28,
    4819 => 28,
    4820 => 28,
    4821 => 28,
    4822 => 28,
    4823 => 28,
    4824 => 28,
    4825 => 28,
    4826 => 28,
    4827 => 28,
    4828 => 28,
    4829 => 28,
    4830 => 28,
    4831 => 28,
    4832 => 28,
    4833 => 28,
    4834 => 28,
    4835 => 28,
    4836 => 28,
    4837 => 28,
    4838 => 28,
    4839 => 28,
    4840 => 28,
    4841 => 28,
    4842 => 28,
    4843 => 28,
    4844 => 28,
    4845 => 28,
    4846 => 28,
    4847 => 28,
    4848 => 28,
    4849 => 28,
    4850 => 28,
    4851 => 28,
    4852 => 28,
    4853 => 28,
    4854 => 28,
    4855 => 28,
    4856 => 28,
    4857 => 28,
    4858 => 28,
    4859 => 28,
    4860 => 28,
    4861 => 28,
    4862 => 28,
    4863 => 28,
    4864 => 28,
    4865 => 28,
    4866 => 28,
    4867 => 28,
    4868 => 28,
    4869 => 28,
    4870 => 28,
    4871 => 28,
    4872 => 28,
    4873 => 28,
    4874 => 28,
    4875 => 28,
    4876 => 28,
    4877 => 28,
    4878 => 28,
    4879 => 28,
    4880 => 28,
    4881 => 28,
    4882 => 28,
    4883 => 28,
    4884 => 28,
    4885 => 28,
    4886 => 28,
    4887 => 28,
    4888 => 28,
    4889 => 28,
    4890 => 28,
    4891 => 28,
    4892 => 28,
    4893 => 28,
    4894 => 28,
    4895 => 28,
    4896 => 28,
    4897 => 29,
    4898 => 29,
    4899 => 29,
    4900 => 29,
    4901 => 29,
    4902 => 29,
    4903 => 29,
    4904 => 29,
    4905 => 29,
    4906 => 29,
    4907 => 29,
    4908 => 29,
    4909 => 29,
    4910 => 29,
    4911 => 29,
    4912 => 29,
    4913 => 29,
    4914 => 29,
    4915 => 29,
    4916 => 29,
    4917 => 29,
    4918 => 29,
    4919 => 29,
    4920 => 29,
    4921 => 29,
    4922 => 29,
    4923 => 29,
    4924 => 29,
    4925 => 29,
    4926 => 29,
    4927 => 29,
    4928 => 29,
    4929 => 29,
    4930 => 29,
    4931 => 29,
    4932 => 29,
    4933 => 29,
    4934 => 29,
    4935 => 29,
    4936 => 29,
    4937 => 29,
    4938 => 29,
    4939 => 29,
    4940 => 29,
    4941 => 29,
    4942 => 29,
    4943 => 29,
    4944 => 29,
    4945 => 29,
    4946 => 29,
    4947 => 29,
    4948 => 29,
    4949 => 29,
    4950 => 29,
    4951 => 29,
    4952 => 29,
    4953 => 29,
    4954 => 29,
    4955 => 29,
    4956 => 29,
    4957 => 29,
    4958 => 29,
    4959 => 29,
    4960 => 29,
    4961 => 29,
    4962 => 29,
    4963 => 29,
    4964 => 29,
    4965 => 29,
    4966 => 29,
    4967 => 29,
    4968 => 29,
    4969 => 29,
    4970 => 29,
    4971 => 29,
    4972 => 29,
    4973 => 29,
    4974 => 29,
    4975 => 29,
    4976 => 29,
    4977 => 29,
    4978 => 29,
    4979 => 29,
    4980 => 29,
    4981 => 29,
    4982 => 29,
    4983 => 29,
    4984 => 29,
    4985 => 29,
    4986 => 29,
    4987 => 29,
    4988 => 29,
    4989 => 29,
    4990 => 29,
    4991 => 29,
    4992 => 29,
    4993 => 29,
    4994 => 29,
    4995 => 29,
    4996 => 29,
    4997 => 29,
    4998 => 29,
    4999 => 29,
    5000 => 29,
    5001 => 29,
    5002 => 29,
    5003 => 29,
    5004 => 29,
    5005 => 29,
    5006 => 29,
    5007 => 29,
    5008 => 29,
    5009 => 29,
    5010 => 29,
    5011 => 29,
    5012 => 29,
    5013 => 29,
    5014 => 29,
    5015 => 29,
    5016 => 29,
    5017 => 29,
    5018 => 29,
    5019 => 29,
    5020 => 29,
    5021 => 29,
    5022 => 29,
    5023 => 29,
    5024 => 29,
    5025 => 29,
    5026 => 29,
    5027 => 29,
    5028 => 29,
    5029 => 29,
    5030 => 29,
    5031 => 29,
    5032 => 29,
    5033 => 29,
    5034 => 29,
    5035 => 29,
    5036 => 29,
    5037 => 29,
    5038 => 29,
    5039 => 29,
    5040 => 29,
    5041 => 29,
    5042 => 29,
    5043 => 29,
    5044 => 29,
    5045 => 29,
    5046 => 29,
    5047 => 29,
    5048 => 29,
    5049 => 29,
    5050 => 29,
    5051 => 29,
    5052 => 29,
    5053 => 29,
    5054 => 29,
    5055 => 29,
    5056 => 29,
    5057 => 29,
    5058 => 29,
    5059 => 29,
    5060 => 29,
    5061 => 29,
    5062 => 29,
    5063 => 29,
    5064 => 29,
    5065 => 29,
    5066 => 29,
    5067 => 29,
    5068 => 29,
    5069 => 29,
    5070 => 29,
    5071 => 29,
    5072 => 29,
    5073 => 29,
    5074 => 29,
    5075 => 29,
    5076 => 29,
    5077 => 29,
    5078 => 29,
    5079 => 29,
    5080 => 29,
    5081 => 29,
    5082 => 29,
    5083 => 30,
    5084 => 30,
    5085 => 30,
    5086 => 30,
    5087 => 30,
    5088 => 30,
    5089 => 30,
    5090 => 30,
    5091 => 30,
    5092 => 30,
    5093 => 30,
    5094 => 30,
    5095 => 30,
    5096 => 30,
    5097 => 30,
    5098 => 30,
    5099 => 30,
    5100 => 30,
    5101 => 30,
    5102 => 30,
    5103 => 30,
    5104 => 30,
    5105 => 30,
    5106 => 30,
    5107 => 30,
    5108 => 30,
    5109 => 30,
    5110 => 30,
    5111 => 30,
    5112 => 30,
    5113 => 30,
    5114 => 30,
    5115 => 30,
    5116 => 30,
    5117 => 30,
    5118 => 30,
    5119 => 30,
    5120 => 30,
    5121 => 30,
    5122 => 30,
    5123 => 30,
    5124 => 30,
    5125 => 30,
    5126 => 30,
    5127 => 30,
    5128 => 30,
    5129 => 30,
    5130 => 30,
    5131 => 30,
    5132 => 30,
    5133 => 30,
    5134 => 30,
    5135 => 30,
    5136 => 30,
    5137 => 30,
    5138 => 30,
    5139 => 30,
    5140 => 30,
    5141 => 30,
    5142 => 30,
    5143 => 30,
    5144 => 30,
    5145 => 30,
    5146 => 30,
    5147 => 30,
    5148 => 30,
    5149 => 30,
    5150 => 30,
    5151 => 30,
    5152 => 30,
    5153 => 30,
    5154 => 30,
    5155 => 30,
    5156 => 30,
    5157 => 30,
    5158 => 30,
    5159 => 30,
    5160 => 30,
    5161 => 30,
    5162 => 30,
    5163 => 30,
    5164 => 30,
    5165 => 30,
    5166 => 30,
    5167 => 30,
    5168 => 30,
    5169 => 30,
    5170 => 30,
    5171 => 30,
    5172 => 30,
    5173 => 30,
    5174 => 30,
    5175 => 30,
    5176 => 30,
    5177 => 30,
    5178 => 30,
    5179 => 30,
    5180 => 30,
    5181 => 30,
    5182 => 30,
    5183 => 30,
    5184 => 30,
    5185 => 30,
    5186 => 30,
    5187 => 30,
    5188 => 30,
    5189 => 30,
    5190 => 30,
    5191 => 30,
    5192 => 30,
    5193 => 30,
    5194 => 30,
    5195 => 30,
    5196 => 30,
    5197 => 30,
    5198 => 30,
    5199 => 30,
    5200 => 30,
    5201 => 30,
    5202 => 30,
    5203 => 30,
    5204 => 30,
    5205 => 30,
    5206 => 30,
    5207 => 30,
    5208 => 30,
    5209 => 30,
    5210 => 30,
    5211 => 30,
    5212 => 30,
    5213 => 30,
    5214 => 30,
    5215 => 30,
    5216 => 30,
    5217 => 30,
    5218 => 30,
    5219 => 30,
    5220 => 30,
    5221 => 30,
    5222 => 30,
    5223 => 30,
    5224 => 30,
    5225 => 30,
    5226 => 30,
    5227 => 30,
    5228 => 30,
    5229 => 30,
    5230 => 30,
    5231 => 30,
    5232 => 30,
    5233 => 30,
    5234 => 30,
    5235 => 30,
    5236 => 30,
    5237 => 30,
    5238 => 30,
    5239 => 30,
    5240 => 30,
    5241 => 30,
    5242 => 30,
    5243 => 30,
    5244 => 30,
    5245 => 30,
    5246 => 30,
    5247 => 30,
    5248 => 30,
    5249 => 30,
    5250 => 30,
    5251 => 30,
    5252 => 30,
    5253 => 30,
    5254 => 30,
    5255 => 30,
    5256 => 30,
    5257 => 30,
    5258 => 30,
    5259 => 30,
    5260 => 30,
    5261 => 30,
    5262 => 30,
    5263 => 30,
    5264 => 30,
    5265 => 30,
    5266 => 30,
    5267 => 30,
    5268 => 30,
    5269 => 30,
    5270 => 30,
    5271 => 30,
    5272 => 31,
    5273 => 31,
    5274 => 31,
    5275 => 31,
    5276 => 31,
    5277 => 31,
    5278 => 31,
    5279 => 31,
    5280 => 31,
    5281 => 31,
    5282 => 31,
    5283 => 31,
    5284 => 31,
    5285 => 31,
    5286 => 31,
    5287 => 31,
    5288 => 31,
    5289 => 31,
    5290 => 31,
    5291 => 31,
    5292 => 31,
    5293 => 31,
    5294 => 31,
    5295 => 31,
    5296 => 31,
    5297 => 31,
    5298 => 31,
    5299 => 31,
    5300 => 31,
    5301 => 31,
    5302 => 31,
    5303 => 31,
    5304 => 31,
    5305 => 31,
    5306 => 31,
    5307 => 31,
    5308 => 31,
    5309 => 31,
    5310 => 31,
    5311 => 31,
    5312 => 31,
    5313 => 31,
    5314 => 31,
    5315 => 31,
    5316 => 31,
    5317 => 31,
    5318 => 31,
    5319 => 31,
    5320 => 31,
    5321 => 31,
    5322 => 31,
    5323 => 31,
    5324 => 31,
    5325 => 31,
    5326 => 31,
    5327 => 31,
    5328 => 31,
    5329 => 31,
    5330 => 31,
    5331 => 31,
    5332 => 31,
    5333 => 31,
    5334 => 31,
    5335 => 31,
    5336 => 31,
    5337 => 31,
    5338 => 31,
    5339 => 31,
    5340 => 31,
    5341 => 31,
    5342 => 31,
    5343 => 31,
    5344 => 31,
    5345 => 31,
    5346 => 31,
    5347 => 31,
    5348 => 31,
    5349 => 31,
    5350 => 31,
    5351 => 31,
    5352 => 31,
    5353 => 31,
    5354 => 31,
    5355 => 31,
    5356 => 31,
    5357 => 31,
    5358 => 31,
    5359 => 31,
    5360 => 31,
    5361 => 31,
    5362 => 31,
    5363 => 31,
    5364 => 31,
    5365 => 31,
    5366 => 31,
    5367 => 31,
    5368 => 31,
    5369 => 31,
    5370 => 31,
    5371 => 31,
    5372 => 31,
    5373 => 31,
    5374 => 31,
    5375 => 31,
    5376 => 31,
    5377 => 31,
    5378 => 31,
    5379 => 31,
    5380 => 31,
    5381 => 31,
    5382 => 31,
    5383 => 31,
    5384 => 31,
    5385 => 31,
    5386 => 31,
    5387 => 31,
    5388 => 31,
    5389 => 31,
    5390 => 31,
    5391 => 31,
    5392 => 31,
    5393 => 31,
    5394 => 31,
    5395 => 31,
    5396 => 31,
    5397 => 31,
    5398 => 31,
    5399 => 31,
    5400 => 31,
    5401 => 31,
    5402 => 31,
    5403 => 31,
    5404 => 31,
    5405 => 31,
    5406 => 31,
    5407 => 31,
    5408 => 31,
    5409 => 31,
    5410 => 31,
    5411 => 31,
    5412 => 31,
    5413 => 31,
    5414 => 31,
    5415 => 31,
    5416 => 31,
    5417 => 31,
    5418 => 31,
    5419 => 31,
    5420 => 31,
    5421 => 31,
    5422 => 31,
    5423 => 31,
    5424 => 31,
    5425 => 31,
    5426 => 31,
    5427 => 31,
    5428 => 31,
    5429 => 31,
    5430 => 31,
    5431 => 31,
    5432 => 31,
    5433 => 31,
    5434 => 31,
    5435 => 31,
    5436 => 31,
    5437 => 31,
    5438 => 31,
    5439 => 31,
    5440 => 31,
    5441 => 31,
    5442 => 31,
    5443 => 31,
    5444 => 31,
    5445 => 31,
    5446 => 31,
    5447 => 31,
    5448 => 31,
    5449 => 31,
    5450 => 31,
    5451 => 31,
    5452 => 31,
    5453 => 31,
    5454 => 31,
    5455 => 31,
    5456 => 31,
    5457 => 31,
    5458 => 31,
    5459 => 31,
    5460 => 31,
    5461 => 31,
    5462 => 32,
    5463 => 32,
    5464 => 32,
    5465 => 32,
    5466 => 32,
    5467 => 32,
    5468 => 32,
    5469 => 32,
    5470 => 32,
    5471 => 32,
    5472 => 32,
    5473 => 32,
    5474 => 32,
    5475 => 32,
    5476 => 32,
    5477 => 32,
    5478 => 32,
    5479 => 32,
    5480 => 32,
    5481 => 32,
    5482 => 32,
    5483 => 32,
    5484 => 32,
    5485 => 32,
    5486 => 32,
    5487 => 32,
    5488 => 32,
    5489 => 32,
    5490 => 32,
    5491 => 32,
    5492 => 32,
    5493 => 32,
    5494 => 32,
    5495 => 32,
    5496 => 32,
    5497 => 32,
    5498 => 32,
    5499 => 32,
    5500 => 32,
    5501 => 32,
    5502 => 32,
    5503 => 32,
    5504 => 32,
    5505 => 32,
    5506 => 32,
    5507 => 32,
    5508 => 32,
    5509 => 32,
    5510 => 32,
    5511 => 32,
    5512 => 32,
    5513 => 32,
    5514 => 32,
    5515 => 32,
    5516 => 32,
    5517 => 32,
    5518 => 32,
    5519 => 32,
    5520 => 32,
    5521 => 32,
    5522 => 32,
    5523 => 32,
    5524 => 32,
    5525 => 32,
    5526 => 32,
    5527 => 32,
    5528 => 32,
    5529 => 32,
    5530 => 32,
    5531 => 32,
    5532 => 32,
    5533 => 32,
    5534 => 32,
    5535 => 32,
    5536 => 32,
    5537 => 32,
    5538 => 32,
    5539 => 32,
    5540 => 32,
    5541 => 32,
    5542 => 32,
    5543 => 32,
    5544 => 32,
    5545 => 32,
    5546 => 32,
    5547 => 32,
    5548 => 32,
    5549 => 32,
    5550 => 32,
    5551 => 32,
    5552 => 32,
    5553 => 32,
    5554 => 32,
    5555 => 32,
    5556 => 32,
    5557 => 32,
    5558 => 32,
    5559 => 32,
    5560 => 32,
    5561 => 32,
    5562 => 32,
    5563 => 32,
    5564 => 32,
    5565 => 32,
    5566 => 32,
    5567 => 32,
    5568 => 32,
    5569 => 32,
    5570 => 32,
    5571 => 32,
    5572 => 32,
    5573 => 32,
    5574 => 32,
    5575 => 32,
    5576 => 32,
    5577 => 32,
    5578 => 32,
    5579 => 32,
    5580 => 32,
    5581 => 32,
    5582 => 32,
    5583 => 32,
    5584 => 32,
    5585 => 32,
    5586 => 32,
    5587 => 32,
    5588 => 32,
    5589 => 32,
    5590 => 32,
    5591 => 32,
    5592 => 32,
    5593 => 32,
    5594 => 32,
    5595 => 32,
    5596 => 32,
    5597 => 32,
    5598 => 32,
    5599 => 32,
    5600 => 32,
    5601 => 32,
    5602 => 32,
    5603 => 32,
    5604 => 32,
    5605 => 32,
    5606 => 32,
    5607 => 32,
    5608 => 32,
    5609 => 32,
    5610 => 32,
    5611 => 32,
    5612 => 32,
    5613 => 32,
    5614 => 32,
    5615 => 32,
    5616 => 32,
    5617 => 32,
    5618 => 32,
    5619 => 32,
    5620 => 32,
    5621 => 32,
    5622 => 32,
    5623 => 32,
    5624 => 32,
    5625 => 32,
    5626 => 32,
    5627 => 32,
    5628 => 32,
    5629 => 32,
    5630 => 32,
    5631 => 32,
    5632 => 32,
    5633 => 32,
    5634 => 32,
    5635 => 32,
    5636 => 32,
    5637 => 32,
    5638 => 32,
    5639 => 32,
    5640 => 32,
    5641 => 32,
    5642 => 32,
    5643 => 32,
    5644 => 32,
    5645 => 32,
    5646 => 32,
    5647 => 32,
    5648 => 32,
    5649 => 32,
    5650 => 32,
    5651 => 32,
    5652 => 32,
    5653 => 32,
    5654 => 33,
    5655 => 33,
    5656 => 33,
    5657 => 33,
    5658 => 33,
    5659 => 33,
    5660 => 33,
    5661 => 33,
    5662 => 33,
    5663 => 33,
    5664 => 33,
    5665 => 33,
    5666 => 33,
    5667 => 33,
    5668 => 33,
    5669 => 33,
    5670 => 33,
    5671 => 33,
    5672 => 33,
    5673 => 33,
    5674 => 33,
    5675 => 33,
    5676 => 33,
    5677 => 33,
    5678 => 33,
    5679 => 33,
    5680 => 33,
    5681 => 33,
    5682 => 33,
    5683 => 33,
    5684 => 33,
    5685 => 33,
    5686 => 33,
    5687 => 33,
    5688 => 33,
    5689 => 33,
    5690 => 33,
    5691 => 33,
    5692 => 33,
    5693 => 33,
    5694 => 33,
    5695 => 33,
    5696 => 33,
    5697 => 33,
    5698 => 33,
    5699 => 33,
    5700 => 33,
    5701 => 33,
    5702 => 33,
    5703 => 33,
    5704 => 33,
    5705 => 33,
    5706 => 33,
    5707 => 33,
    5708 => 33,
    5709 => 33,
    5710 => 33,
    5711 => 33,
    5712 => 33,
    5713 => 33,
    5714 => 33,
    5715 => 33,
    5716 => 33,
    5717 => 33,
    5718 => 33,
    5719 => 33,
    5720 => 33,
    5721 => 33,
    5722 => 33,
    5723 => 33,
    5724 => 33,
    5725 => 33,
    5726 => 33,
    5727 => 33,
    5728 => 33,
    5729 => 33,
    5730 => 33,
    5731 => 33,
    5732 => 33,
    5733 => 33,
    5734 => 33,
    5735 => 33,
    5736 => 33,
    5737 => 33,
    5738 => 33,
    5739 => 33,
    5740 => 33,
    5741 => 33,
    5742 => 33,
    5743 => 33,
    5744 => 33,
    5745 => 33,
    5746 => 33,
    5747 => 33,
    5748 => 33,
    5749 => 33,
    5750 => 33,
    5751 => 33,
    5752 => 33,
    5753 => 33,
    5754 => 33,
    5755 => 33,
    5756 => 33,
    5757 => 33,
    5758 => 33,
    5759 => 33,
    5760 => 33,
    5761 => 33,
    5762 => 33,
    5763 => 33,
    5764 => 33,
    5765 => 33,
    5766 => 33,
    5767 => 33,
    5768 => 33,
    5769 => 33,
    5770 => 33,
    5771 => 33,
    5772 => 33,
    5773 => 33,
    5774 => 33,
    5775 => 33,
    5776 => 33,
    5777 => 33,
    5778 => 33,
    5779 => 33,
    5780 => 33,
    5781 => 33,
    5782 => 33,
    5783 => 33,
    5784 => 33,
    5785 => 33,
    5786 => 33,
    5787 => 33,
    5788 => 33,
    5789 => 33,
    5790 => 33,
    5791 => 33,
    5792 => 33,
    5793 => 33,
    5794 => 33,
    5795 => 33,
    5796 => 33,
    5797 => 33,
    5798 => 33,
    5799 => 33,
    5800 => 33,
    5801 => 33,
    5802 => 33,
    5803 => 33,
    5804 => 33,
    5805 => 33,
    5806 => 33,
    5807 => 33,
    5808 => 33,
    5809 => 33,
    5810 => 33,
    5811 => 33,
    5812 => 33,
    5813 => 33,
    5814 => 33,
    5815 => 33,
    5816 => 33,
    5817 => 33,
    5818 => 33,
    5819 => 33,
    5820 => 33,
    5821 => 33,
    5822 => 33,
    5823 => 33,
    5824 => 33,
    5825 => 33,
    5826 => 33,
    5827 => 33,
    5828 => 33,
    5829 => 33,
    5830 => 33,
    5831 => 33,
    5832 => 33,
    5833 => 33,
    5834 => 33,
    5835 => 33,
    5836 => 33,
    5837 => 33,
    5838 => 33,
    5839 => 33,
    5840 => 33,
    5841 => 33,
    5842 => 33,
    5843 => 33,
    5844 => 33,
    5845 => 33,
    5846 => 33,
    5847 => 33,
    5848 => 34,
    5849 => 34,
    5850 => 34,
    5851 => 34,
    5852 => 34,
    5853 => 34,
    5854 => 34,
    5855 => 34,
    5856 => 34,
    5857 => 34,
    5858 => 34,
    5859 => 34,
    5860 => 34,
    5861 => 34,
    5862 => 34,
    5863 => 34,
    5864 => 34,
    5865 => 34,
    5866 => 34,
    5867 => 34,
    5868 => 34,
    5869 => 34,
    5870 => 34,
    5871 => 34,
    5872 => 34,
    5873 => 34,
    5874 => 34,
    5875 => 34,
    5876 => 34,
    5877 => 34,
    5878 => 34,
    5879 => 34,
    5880 => 34,
    5881 => 34,
    5882 => 34,
    5883 => 34,
    5884 => 34,
    5885 => 34,
    5886 => 34,
    5887 => 34,
    5888 => 34,
    5889 => 34,
    5890 => 34,
    5891 => 34,
    5892 => 34,
    5893 => 34,
    5894 => 34,
    5895 => 34,
    5896 => 34,
    5897 => 34,
    5898 => 34,
    5899 => 34,
    5900 => 34,
    5901 => 34,
    5902 => 34,
    5903 => 34,
    5904 => 34,
    5905 => 34,
    5906 => 34,
    5907 => 34,
    5908 => 34,
    5909 => 34,
    5910 => 34,
    5911 => 34,
    5912 => 34,
    5913 => 34,
    5914 => 34,
    5915 => 34,
    5916 => 34,
    5917 => 34,
    5918 => 34,
    5919 => 34,
    5920 => 34,
    5921 => 34,
    5922 => 34,
    5923 => 34,
    5924 => 34,
    5925 => 34,
    5926 => 34,
    5927 => 34,
    5928 => 34,
    5929 => 34,
    5930 => 34,
    5931 => 34,
    5932 => 34,
    5933 => 34,
    5934 => 34,
    5935 => 34,
    5936 => 34,
    5937 => 34,
    5938 => 34,
    5939 => 34,
    5940 => 34,
    5941 => 34,
    5942 => 34,
    5943 => 34,
    5944 => 34,
    5945 => 34,
    5946 => 34,
    5947 => 34,
    5948 => 34,
    5949 => 34,
    5950 => 34,
    5951 => 34,
    5952 => 34,
    5953 => 34,
    5954 => 34,
    5955 => 34,
    5956 => 34,
    5957 => 34,
    5958 => 34,
    5959 => 34,
    5960 => 34,
    5961 => 34,
    5962 => 34,
    5963 => 34,
    5964 => 34,
    5965 => 34,
    5966 => 34,
    5967 => 34,
    5968 => 34,
    5969 => 34,
    5970 => 34,
    5971 => 34,
    5972 => 34,
    5973 => 34,
    5974 => 34,
    5975 => 34,
    5976 => 34,
    5977 => 34,
    5978 => 34,
    5979 => 34,
    5980 => 34,
    5981 => 34,
    5982 => 34,
    5983 => 34,
    5984 => 34,
    5985 => 34,
    5986 => 34,
    5987 => 34,
    5988 => 34,
    5989 => 34,
    5990 => 34,
    5991 => 34,
    5992 => 34,
    5993 => 34,
    5994 => 34,
    5995 => 34,
    5996 => 34,
    5997 => 34,
    5998 => 34,
    5999 => 34,
    6000 => 34,
    6001 => 34,
    6002 => 34,
    6003 => 34,
    6004 => 34,
    6005 => 34,
    6006 => 34,
    6007 => 34,
    6008 => 34,
    6009 => 34,
    6010 => 34,
    6011 => 34,
    6012 => 34,
    6013 => 34,
    6014 => 34,
    6015 => 34,
    6016 => 34,
    6017 => 34,
    6018 => 34,
    6019 => 34,
    6020 => 34,
    6021 => 34,
    6022 => 34,
    6023 => 34,
    6024 => 34,
    6025 => 34,
    6026 => 34,
    6027 => 34,
    6028 => 34,
    6029 => 34,
    6030 => 34,
    6031 => 34,
    6032 => 34,
    6033 => 34,
    6034 => 34,
    6035 => 34,
    6036 => 34,
    6037 => 34,
    6038 => 34,
    6039 => 34,
    6040 => 34,
    6041 => 34,
    6042 => 34,
    6043 => 34,
    6044 => 34,
    6045 => 35,
    6046 => 35,
    6047 => 35,
    6048 => 35,
    6049 => 35,
    6050 => 35,
    6051 => 35,
    6052 => 35,
    6053 => 35,
    6054 => 35,
    6055 => 35,
    6056 => 35,
    6057 => 35,
    6058 => 35,
    6059 => 35,
    6060 => 35,
    6061 => 35,
    6062 => 35,
    6063 => 35,
    6064 => 35,
    6065 => 35,
    6066 => 35,
    6067 => 35,
    6068 => 35,
    6069 => 35,
    6070 => 35,
    6071 => 35,
    6072 => 35,
    6073 => 35,
    6074 => 35,
    6075 => 35,
    6076 => 35,
    6077 => 35,
    6078 => 35,
    6079 => 35,
    6080 => 35,
    6081 => 35,
    6082 => 35,
    6083 => 35,
    6084 => 35,
    6085 => 35,
    6086 => 35,
    6087 => 35,
    6088 => 35,
    6089 => 35,
    6090 => 35,
    6091 => 35,
    6092 => 35,
    6093 => 35,
    6094 => 35,
    6095 => 35,
    6096 => 35,
    6097 => 35,
    6098 => 35,
    6099 => 35,
    6100 => 35,
    6101 => 35,
    6102 => 35,
    6103 => 35,
    6104 => 35,
    6105 => 35,
    6106 => 35,
    6107 => 35,
    6108 => 35,
    6109 => 35,
    6110 => 35,
    6111 => 35,
    6112 => 35,
    6113 => 35,
    6114 => 35,
    6115 => 35,
    6116 => 35,
    6117 => 35,
    6118 => 35,
    6119 => 35,
    6120 => 35,
    6121 => 35,
    6122 => 35,
    6123 => 35,
    6124 => 35,
    6125 => 35,
    6126 => 35,
    6127 => 35,
    6128 => 35,
    6129 => 35,
    6130 => 35,
    6131 => 35,
    6132 => 35,
    6133 => 35,
    6134 => 35,
    6135 => 35,
    6136 => 35,
    6137 => 35,
    6138 => 35,
    6139 => 35,
    6140 => 35,
    6141 => 35,
    6142 => 35,
    6143 => 35,
    6144 => 35,
    6145 => 35,
    6146 => 35,
    6147 => 35,
    6148 => 35,
    6149 => 35,
    6150 => 35,
    6151 => 35,
    6152 => 35,
    6153 => 35,
    6154 => 35,
    6155 => 35,
    6156 => 35,
    6157 => 35,
    6158 => 35,
    6159 => 35,
    6160 => 35,
    6161 => 35,
    6162 => 35,
    6163 => 35,
    6164 => 35,
    6165 => 35,
    6166 => 35,
    6167 => 35,
    6168 => 35,
    6169 => 35,
    6170 => 35,
    6171 => 35,
    6172 => 35,
    6173 => 35,
    6174 => 35,
    6175 => 35,
    6176 => 35,
    6177 => 35,
    6178 => 35,
    6179 => 35,
    6180 => 35,
    6181 => 35,
    6182 => 35,
    6183 => 35,
    6184 => 35,
    6185 => 35,
    6186 => 35,
    6187 => 35,
    6188 => 35,
    6189 => 35,
    6190 => 35,
    6191 => 35,
    6192 => 35,
    6193 => 35,
    6194 => 35,
    6195 => 35,
    6196 => 35,
    6197 => 35,
    6198 => 35,
    6199 => 35,
    6200 => 35,
    6201 => 35,
    6202 => 35,
    6203 => 35,
    6204 => 35,
    6205 => 35,
    6206 => 35,
    6207 => 35,
    6208 => 35,
    6209 => 35,
    6210 => 35,
    6211 => 35,
    6212 => 35,
    6213 => 35,
    6214 => 35,
    6215 => 35,
    6216 => 35,
    6217 => 35,
    6218 => 35,
    6219 => 35,
    6220 => 35,
    6221 => 35,
    6222 => 35,
    6223 => 35,
    6224 => 35,
    6225 => 35,
    6226 => 35,
    6227 => 35,
    6228 => 35,
    6229 => 35,
    6230 => 35,
    6231 => 35,
    6232 => 35,
    6233 => 35,
    6234 => 35,
    6235 => 35,
    6236 => 35,
    6237 => 35,
    6238 => 35,
    6239 => 35,
    6240 => 35,
    6241 => 35,
    6242 => 35,
    6243 => 35,
    6244 => 36,
    6245 => 36,
    6246 => 36,
    6247 => 36,
    6248 => 36,
    6249 => 36,
    6250 => 36,
    6251 => 36,
    6252 => 36,
    6253 => 36,
    6254 => 36,
    6255 => 36,
    6256 => 36,
    6257 => 36,
    6258 => 36,
    6259 => 36,
    6260 => 36,
    6261 => 36,
    6262 => 36,
    6263 => 36,
    6264 => 36,
    6265 => 36,
    6266 => 36,
    6267 => 36,
    6268 => 36,
    6269 => 36,
    6270 => 36,
    6271 => 36,
    6272 => 36,
    6273 => 36,
    6274 => 36,
    6275 => 36,
    6276 => 36,
    6277 => 36,
    6278 => 36,
    6279 => 36,
    6280 => 36,
    6281 => 36,
    6282 => 36,
    6283 => 36,
    6284 => 36,
    6285 => 36,
    6286 => 36,
    6287 => 36,
    6288 => 36,
    6289 => 36,
    6290 => 36,
    6291 => 36,
    6292 => 36,
    6293 => 36,
    6294 => 36,
    6295 => 36,
    6296 => 36,
    6297 => 36,
    6298 => 36,
    6299 => 36,
    6300 => 36,
    6301 => 36,
    6302 => 36,
    6303 => 36,
    6304 => 36,
    6305 => 36,
    6306 => 36,
    6307 => 36,
    6308 => 36,
    6309 => 36,
    6310 => 36,
    6311 => 36,
    6312 => 36,
    6313 => 36,
    6314 => 36,
    6315 => 36,
    6316 => 36,
    6317 => 36,
    6318 => 36,
    6319 => 36,
    6320 => 36,
    6321 => 36,
    6322 => 36,
    6323 => 36,
    6324 => 36,
    6325 => 36,
    6326 => 36,
    6327 => 36,
    6328 => 36,
    6329 => 36,
    6330 => 36,
    6331 => 36,
    6332 => 36,
    6333 => 36,
    6334 => 36,
    6335 => 36,
    6336 => 36,
    6337 => 36,
    6338 => 36,
    6339 => 36,
    6340 => 36,
    6341 => 36,
    6342 => 36,
    6343 => 36,
    6344 => 36,
    6345 => 36,
    6346 => 36,
    6347 => 36,
    6348 => 36,
    6349 => 36,
    6350 => 36,
    6351 => 36,
    6352 => 36,
    6353 => 36,
    6354 => 36,
    6355 => 36,
    6356 => 36,
    6357 => 36,
    6358 => 36,
    6359 => 36,
    6360 => 36,
    6361 => 36,
    6362 => 36,
    6363 => 36,
    6364 => 36,
    6365 => 36,
    6366 => 36,
    6367 => 36,
    6368 => 36,
    6369 => 36,
    6370 => 36,
    6371 => 36,
    6372 => 36,
    6373 => 36,
    6374 => 36,
    6375 => 36,
    6376 => 36,
    6377 => 36,
    6378 => 36,
    6379 => 36,
    6380 => 36,
    6381 => 36,
    6382 => 36,
    6383 => 36,
    6384 => 36,
    6385 => 36,
    6386 => 36,
    6387 => 36,
    6388 => 36,
    6389 => 36,
    6390 => 36,
    6391 => 36,
    6392 => 36,
    6393 => 36,
    6394 => 36,
    6395 => 36,
    6396 => 36,
    6397 => 36,
    6398 => 36,
    6399 => 36,
    6400 => 36,
    6401 => 36,
    6402 => 36,
    6403 => 36,
    6404 => 36,
    6405 => 36,
    6406 => 36,
    6407 => 36,
    6408 => 36,
    6409 => 36,
    6410 => 36,
    6411 => 36,
    6412 => 36,
    6413 => 36,
    6414 => 36,
    6415 => 36,
    6416 => 36,
    6417 => 36,
    6418 => 36,
    6419 => 36,
    6420 => 36,
    6421 => 36,
    6422 => 36,
    6423 => 36,
    6424 => 36,
    6425 => 36,
    6426 => 36,
    6427 => 36,
    6428 => 36,
    6429 => 36,
    6430 => 36,
    6431 => 36,
    6432 => 36,
    6433 => 36,
    6434 => 36,
    6435 => 36,
    6436 => 36,
    6437 => 36,
    6438 => 36,
    6439 => 36,
    6440 => 36,
    6441 => 36,
    6442 => 36,
    6443 => 36,
    6444 => 36,
    6445 => 36,
    6446 => 37,
    6447 => 37,
    6448 => 37,
    6449 => 37,
    6450 => 37,
    6451 => 37,
    6452 => 37,
    6453 => 37,
    6454 => 37,
    6455 => 37,
    6456 => 37,
    6457 => 37,
    6458 => 37,
    6459 => 37,
    6460 => 37,
    6461 => 37,
    6462 => 37,
    6463 => 37,
    6464 => 37,
    6465 => 37,
    6466 => 37,
    6467 => 37,
    6468 => 37,
    6469 => 37,
    6470 => 37,
    6471 => 37,
    6472 => 37,
    6473 => 37,
    6474 => 37,
    6475 => 37,
    6476 => 37,
    6477 => 37,
    6478 => 37,
    6479 => 37,
    6480 => 37,
    6481 => 37,
    6482 => 37,
    6483 => 37,
    6484 => 37,
    6485 => 37,
    6486 => 37,
    6487 => 37,
    6488 => 37,
    6489 => 37,
    6490 => 37,
    6491 => 37,
    6492 => 37,
    6493 => 37,
    6494 => 37,
    6495 => 37,
    6496 => 37,
    6497 => 37,
    6498 => 37,
    6499 => 37,
    6500 => 37,
    6501 => 37,
    6502 => 37,
    6503 => 37,
    6504 => 37,
    6505 => 37,
    6506 => 37,
    6507 => 37,
    6508 => 37,
    6509 => 37,
    6510 => 37,
    6511 => 37,
    6512 => 37,
    6513 => 37,
    6514 => 37,
    6515 => 37,
    6516 => 37,
    6517 => 37,
    6518 => 37,
    6519 => 37,
    6520 => 37,
    6521 => 37,
    6522 => 37,
    6523 => 37,
    6524 => 37,
    6525 => 37,
    6526 => 37,
    6527 => 37,
    6528 => 37,
    6529 => 37,
    6530 => 37,
    6531 => 37,
    6532 => 37,
    6533 => 37,
    6534 => 37,
    6535 => 37,
    6536 => 37,
    6537 => 37,
    6538 => 37,
    6539 => 37,
    6540 => 37,
    6541 => 37,
    6542 => 37,
    6543 => 37,
    6544 => 37,
    6545 => 37,
    6546 => 37,
    6547 => 37,
    6548 => 37,
    6549 => 37,
    6550 => 37,
    6551 => 37,
    6552 => 37,
    6553 => 37,
    6554 => 37,
    6555 => 37,
    6556 => 37,
    6557 => 37,
    6558 => 37,
    6559 => 37,
    6560 => 37,
    6561 => 37,
    6562 => 37,
    6563 => 37,
    6564 => 37,
    6565 => 37,
    6566 => 37,
    6567 => 37,
    6568 => 37,
    6569 => 37,
    6570 => 37,
    6571 => 37,
    6572 => 37,
    6573 => 37,
    6574 => 37,
    6575 => 37,
    6576 => 37,
    6577 => 37,
    6578 => 37,
    6579 => 37,
    6580 => 37,
    6581 => 37,
    6582 => 37,
    6583 => 37,
    6584 => 37,
    6585 => 37,
    6586 => 37,
    6587 => 37,
    6588 => 37,
    6589 => 37,
    6590 => 37,
    6591 => 37,
    6592 => 37,
    6593 => 37,
    6594 => 37,
    6595 => 37,
    6596 => 37,
    6597 => 37,
    6598 => 37,
    6599 => 37,
    6600 => 37,
    6601 => 37,
    6602 => 37,
    6603 => 37,
    6604 => 37,
    6605 => 37,
    6606 => 37,
    6607 => 37,
    6608 => 37,
    6609 => 37,
    6610 => 37,
    6611 => 37,
    6612 => 37,
    6613 => 37,
    6614 => 37,
    6615 => 37,
    6616 => 37,
    6617 => 37,
    6618 => 37,
    6619 => 37,
    6620 => 37,
    6621 => 37,
    6622 => 37,
    6623 => 37,
    6624 => 37,
    6625 => 37,
    6626 => 37,
    6627 => 37,
    6628 => 37,
    6629 => 37,
    6630 => 37,
    6631 => 37,
    6632 => 37,
    6633 => 37,
    6634 => 37,
    6635 => 37,
    6636 => 37,
    6637 => 37,
    6638 => 37,
    6639 => 37,
    6640 => 37,
    6641 => 37,
    6642 => 37,
    6643 => 37,
    6644 => 37,
    6645 => 37,
    6646 => 37,
    6647 => 37,
    6648 => 37,
    6649 => 37,
    6650 => 37,
    6651 => 38,
    6652 => 38,
    6653 => 38,
    6654 => 38,
    6655 => 38,
    6656 => 38,
    6657 => 38,
    6658 => 38,
    6659 => 38,
    6660 => 38,
    6661 => 38,
    6662 => 38,
    6663 => 38,
    6664 => 38,
    6665 => 38,
    6666 => 38,
    6667 => 38,
    6668 => 38,
    6669 => 38,
    6670 => 38,
    6671 => 38,
    6672 => 38,
    6673 => 38,
    6674 => 38,
    6675 => 38,
    6676 => 38,
    6677 => 38,
    6678 => 38,
    6679 => 38,
    6680 => 38,
    6681 => 38,
    6682 => 38,
    6683 => 38,
    6684 => 38,
    6685 => 38,
    6686 => 38,
    6687 => 38,
    6688 => 38,
    6689 => 38,
    6690 => 38,
    6691 => 38,
    6692 => 38,
    6693 => 38,
    6694 => 38,
    6695 => 38,
    6696 => 38,
    6697 => 38,
    6698 => 38,
    6699 => 38,
    6700 => 38,
    6701 => 38,
    6702 => 38,
    6703 => 38,
    6704 => 38,
    6705 => 38,
    6706 => 38,
    6707 => 38,
    6708 => 38,
    6709 => 38,
    6710 => 38,
    6711 => 38,
    6712 => 38,
    6713 => 38,
    6714 => 38,
    6715 => 38,
    6716 => 38,
    6717 => 38,
    6718 => 38,
    6719 => 38,
    6720 => 38,
    6721 => 38,
    6722 => 38,
    6723 => 38,
    6724 => 38,
    6725 => 38,
    6726 => 38,
    6727 => 38,
    6728 => 38,
    6729 => 38,
    6730 => 38,
    6731 => 38,
    6732 => 38,
    6733 => 38,
    6734 => 38,
    6735 => 38,
    6736 => 38,
    6737 => 38,
    6738 => 38,
    6739 => 38,
    6740 => 38,
    6741 => 38,
    6742 => 38,
    6743 => 38,
    6744 => 38,
    6745 => 38,
    6746 => 38,
    6747 => 38,
    6748 => 38,
    6749 => 38,
    6750 => 38,
    6751 => 38,
    6752 => 38,
    6753 => 38,
    6754 => 38,
    6755 => 38,
    6756 => 38,
    6757 => 38,
    6758 => 38,
    6759 => 38,
    6760 => 38,
    6761 => 38,
    6762 => 38,
    6763 => 38,
    6764 => 38,
    6765 => 38,
    6766 => 38,
    6767 => 38,
    6768 => 38,
    6769 => 38,
    6770 => 38,
    6771 => 38,
    6772 => 38,
    6773 => 38,
    6774 => 38,
    6775 => 38,
    6776 => 38,
    6777 => 38,
    6778 => 38,
    6779 => 38,
    6780 => 38,
    6781 => 38,
    6782 => 38,
    6783 => 38,
    6784 => 38,
    6785 => 38,
    6786 => 38,
    6787 => 38,
    6788 => 38,
    6789 => 38,
    6790 => 38,
    6791 => 38,
    6792 => 38,
    6793 => 38,
    6794 => 38,
    6795 => 38,
    6796 => 38,
    6797 => 38,
    6798 => 38,
    6799 => 38,
    6800 => 38,
    6801 => 38,
    6802 => 38,
    6803 => 38,
    6804 => 38,
    6805 => 38,
    6806 => 38,
    6807 => 38,
    6808 => 38,
    6809 => 38,
    6810 => 38,
    6811 => 38,
    6812 => 38,
    6813 => 38,
    6814 => 38,
    6815 => 38,
    6816 => 38,
    6817 => 38,
    6818 => 38,
    6819 => 38,
    6820 => 38,
    6821 => 38,
    6822 => 38,
    6823 => 38,
    6824 => 38,
    6825 => 38,
    6826 => 38,
    6827 => 38,
    6828 => 38,
    6829 => 38,
    6830 => 38,
    6831 => 38,
    6832 => 38,
    6833 => 38,
    6834 => 38,
    6835 => 38,
    6836 => 38,
    6837 => 38,
    6838 => 38,
    6839 => 38,
    6840 => 38,
    6841 => 38,
    6842 => 38,
    6843 => 38,
    6844 => 38,
    6845 => 38,
    6846 => 38,
    6847 => 38,
    6848 => 38,
    6849 => 38,
    6850 => 38,
    6851 => 38,
    6852 => 38,
    6853 => 38,
    6854 => 38,
    6855 => 38,
    6856 => 38,
    6857 => 38,
    6858 => 39,
    6859 => 39,
    6860 => 39,
    6861 => 39,
    6862 => 39,
    6863 => 39,
    6864 => 39,
    6865 => 39,
    6866 => 39,
    6867 => 39,
    6868 => 39,
    6869 => 39,
    6870 => 39,
    6871 => 39,
    6872 => 39,
    6873 => 39,
    6874 => 39,
    6875 => 39,
    6876 => 39,
    6877 => 39,
    6878 => 39,
    6879 => 39,
    6880 => 39,
    6881 => 39,
    6882 => 39,
    6883 => 39,
    6884 => 39,
    6885 => 39,
    6886 => 39,
    6887 => 39,
    6888 => 39,
    6889 => 39,
    6890 => 39,
    6891 => 39,
    6892 => 39,
    6893 => 39,
    6894 => 39,
    6895 => 39,
    6896 => 39,
    6897 => 39,
    6898 => 39,
    6899 => 39,
    6900 => 39,
    6901 => 39,
    6902 => 39,
    6903 => 39,
    6904 => 39,
    6905 => 39,
    6906 => 39,
    6907 => 39,
    6908 => 39,
    6909 => 39,
    6910 => 39,
    6911 => 39,
    6912 => 39,
    6913 => 39,
    6914 => 39,
    6915 => 39,
    6916 => 39,
    6917 => 39,
    6918 => 39,
    6919 => 39,
    6920 => 39,
    6921 => 39,
    6922 => 39,
    6923 => 39,
    6924 => 39,
    6925 => 39,
    6926 => 39,
    6927 => 39,
    6928 => 39,
    6929 => 39,
    6930 => 39,
    6931 => 39,
    6932 => 39,
    6933 => 39,
    6934 => 39,
    6935 => 39,
    6936 => 39,
    6937 => 39,
    6938 => 39,
    6939 => 39,
    6940 => 39,
    6941 => 39,
    6942 => 39,
    6943 => 39,
    6944 => 39,
    6945 => 39,
    6946 => 39,
    6947 => 39,
    6948 => 39,
    6949 => 39,
    6950 => 39,
    6951 => 39,
    6952 => 39,
    6953 => 39,
    6954 => 39,
    6955 => 39,
    6956 => 39,
    6957 => 39,
    6958 => 39,
    6959 => 39,
    6960 => 39,
    6961 => 39,
    6962 => 39,
    6963 => 39,
    6964 => 39,
    6965 => 39,
    6966 => 39,
    6967 => 39,
    6968 => 39,
    6969 => 39,
    6970 => 39,
    6971 => 39,
    6972 => 39,
    6973 => 39,
    6974 => 39,
    6975 => 39,
    6976 => 39,
    6977 => 39,
    6978 => 39,
    6979 => 39,
    6980 => 39,
    6981 => 39,
    6982 => 39,
    6983 => 39,
    6984 => 39,
    6985 => 39,
    6986 => 39,
    6987 => 39,
    6988 => 39,
    6989 => 39,
    6990 => 39,
    6991 => 39,
    6992 => 39,
    6993 => 39,
    6994 => 39,
    6995 => 39,
    6996 => 39,
    6997 => 39,
    6998 => 39,
    6999 => 39,
    7000 => 39,
    7001 => 39,
    7002 => 39,
    7003 => 39,
    7004 => 39,
    7005 => 39,
    7006 => 39,
    7007 => 39,
    7008 => 39,
    7009 => 39,
    7010 => 39,
    7011 => 39,
    7012 => 39,
    7013 => 39,
    7014 => 39,
    7015 => 39,
    7016 => 39,
    7017 => 39,
    7018 => 39,
    7019 => 39,
    7020 => 39,
    7021 => 39,
    7022 => 39,
    7023 => 39,
    7024 => 39,
    7025 => 39,
    7026 => 39,
    7027 => 39,
    7028 => 39,
    7029 => 39,
    7030 => 39,
    7031 => 39,
    7032 => 39,
    7033 => 39,
    7034 => 39,
    7035 => 39,
    7036 => 39,
    7037 => 39,
    7038 => 39,
    7039 => 39,
    7040 => 39,
    7041 => 39,
    7042 => 39,
    7043 => 39,
    7044 => 39,
    7045 => 39,
    7046 => 39,
    7047 => 39,
    7048 => 39,
    7049 => 39,
    7050 => 39,
    7051 => 39,
    7052 => 39,
    7053 => 39,
    7054 => 39,
    7055 => 39,
    7056 => 39,
    7057 => 39,
    7058 => 39,
    7059 => 39,
    7060 => 39,
    7061 => 39,
    7062 => 39,
    7063 => 39,
    7064 => 39,
    7065 => 39,
    7066 => 39,
    7067 => 39,
    7068 => 39,
    7069 => 40,
    7070 => 40,
    7071 => 40,
    7072 => 40,
    7073 => 40,
    7074 => 40,
    7075 => 40,
    7076 => 40,
    7077 => 40,
    7078 => 40,
    7079 => 40,
    7080 => 40,
    7081 => 40,
    7082 => 40,
    7083 => 40,
    7084 => 40,
    7085 => 40,
    7086 => 40,
    7087 => 40,
    7088 => 40,
    7089 => 40,
    7090 => 40,
    7091 => 40,
    7092 => 40,
    7093 => 40,
    7094 => 40,
    7095 => 40,
    7096 => 40,
    7097 => 40,
    7098 => 40,
    7099 => 40,
    7100 => 40,
    7101 => 40,
    7102 => 40,
    7103 => 40,
    7104 => 40,
    7105 => 40,
    7106 => 40,
    7107 => 40,
    7108 => 40,
    7109 => 40,
    7110 => 40,
    7111 => 40,
    7112 => 40,
    7113 => 40,
    7114 => 40,
    7115 => 40,
    7116 => 40,
    7117 => 40,
    7118 => 40,
    7119 => 40,
    7120 => 40,
    7121 => 40,
    7122 => 40,
    7123 => 40,
    7124 => 40,
    7125 => 40,
    7126 => 40,
    7127 => 40,
    7128 => 40,
    7129 => 40,
    7130 => 40,
    7131 => 40,
    7132 => 40,
    7133 => 40,
    7134 => 40,
    7135 => 40,
    7136 => 40,
    7137 => 40,
    7138 => 40,
    7139 => 40,
    7140 => 40,
    7141 => 40,
    7142 => 40,
    7143 => 40,
    7144 => 40,
    7145 => 40,
    7146 => 40,
    7147 => 40,
    7148 => 40,
    7149 => 40,
    7150 => 40,
    7151 => 40,
    7152 => 40,
    7153 => 40,
    7154 => 40,
    7155 => 40,
    7156 => 40,
    7157 => 40,
    7158 => 40,
    7159 => 40,
    7160 => 40,
    7161 => 40,
    7162 => 40,
    7163 => 40,
    7164 => 40,
    7165 => 40,
    7166 => 40,
    7167 => 40,
    7168 => 40,
    7169 => 40,
    7170 => 40,
    7171 => 40,
    7172 => 40,
    7173 => 40,
    7174 => 40,
    7175 => 40,
    7176 => 40,
    7177 => 40,
    7178 => 40,
    7179 => 40,
    7180 => 40,
    7181 => 40,
    7182 => 40,
    7183 => 40,
    7184 => 40,
    7185 => 40,
    7186 => 40,
    7187 => 40,
    7188 => 40,
    7189 => 40,
    7190 => 40,
    7191 => 40,
    7192 => 40,
    7193 => 40,
    7194 => 40,
    7195 => 40,
    7196 => 40,
    7197 => 40,
    7198 => 40,
    7199 => 40,
    7200 => 40,
    7201 => 40,
    7202 => 40,
    7203 => 40,
    7204 => 40,
    7205 => 40,
    7206 => 40,
    7207 => 40,
    7208 => 40,
    7209 => 40,
    7210 => 40,
    7211 => 40,
    7212 => 40,
    7213 => 40,
    7214 => 40,
    7215 => 40,
    7216 => 40,
    7217 => 40,
    7218 => 40,
    7219 => 40,
    7220 => 40,
    7221 => 40,
    7222 => 40,
    7223 => 40,
    7224 => 40,
    7225 => 40,
    7226 => 40,
    7227 => 40,
    7228 => 40,
    7229 => 40,
    7230 => 40,
    7231 => 40,
    7232 => 40,
    7233 => 40,
    7234 => 40,
    7235 => 40,
    7236 => 40,
    7237 => 40,
    7238 => 40,
    7239 => 40,
    7240 => 40,
    7241 => 40,
    7242 => 40,
    7243 => 40,
    7244 => 40,
    7245 => 40,
    7246 => 40,
    7247 => 40,
    7248 => 40,
    7249 => 40,
    7250 => 40,
    7251 => 40,
    7252 => 40,
    7253 => 40,
    7254 => 40,
    7255 => 40,
    7256 => 40,
    7257 => 40,
    7258 => 40,
    7259 => 40,
    7260 => 40,
    7261 => 40,
    7262 => 40,
    7263 => 40,
    7264 => 40,
    7265 => 40,
    7266 => 40,
    7267 => 40,
    7268 => 40,
    7269 => 40,
    7270 => 40,
    7271 => 40,
    7272 => 40,
    7273 => 40,
    7274 => 40,
    7275 => 40,
    7276 => 40,
    7277 => 40,
    7278 => 40,
    7279 => 40,
    7280 => 40,
    7281 => 40,
    7282 => 40,
    7283 => 41,
    7284 => 41,
    7285 => 41,
    7286 => 41,
    7287 => 41,
    7288 => 41,
    7289 => 41,
    7290 => 41,
    7291 => 41,
    7292 => 41,
    7293 => 41,
    7294 => 41,
    7295 => 41,
    7296 => 41,
    7297 => 41,
    7298 => 41,
    7299 => 41,
    7300 => 41,
    7301 => 41,
    7302 => 41,
    7303 => 41,
    7304 => 41,
    7305 => 41,
    7306 => 41,
    7307 => 41,
    7308 => 41,
    7309 => 41,
    7310 => 41,
    7311 => 41,
    7312 => 41,
    7313 => 41,
    7314 => 41,
    7315 => 41,
    7316 => 41,
    7317 => 41,
    7318 => 41,
    7319 => 41,
    7320 => 41,
    7321 => 41,
    7322 => 41,
    7323 => 41,
    7324 => 41,
    7325 => 41,
    7326 => 41,
    7327 => 41,
    7328 => 41,
    7329 => 41,
    7330 => 41,
    7331 => 41,
    7332 => 41,
    7333 => 41,
    7334 => 41,
    7335 => 41,
    7336 => 41,
    7337 => 41,
    7338 => 41,
    7339 => 41,
    7340 => 41,
    7341 => 41,
    7342 => 41,
    7343 => 41,
    7344 => 41,
    7345 => 41,
    7346 => 41,
    7347 => 41,
    7348 => 41,
    7349 => 41,
    7350 => 41,
    7351 => 41,
    7352 => 41,
    7353 => 41,
    7354 => 41,
    7355 => 41,
    7356 => 41,
    7357 => 41,
    7358 => 41,
    7359 => 41,
    7360 => 41,
    7361 => 41,
    7362 => 41,
    7363 => 41,
    7364 => 41,
    7365 => 41,
    7366 => 41,
    7367 => 41,
    7368 => 41,
    7369 => 41,
    7370 => 41,
    7371 => 41,
    7372 => 41,
    7373 => 41,
    7374 => 41,
    7375 => 41,
    7376 => 41,
    7377 => 41,
    7378 => 41,
    7379 => 41,
    7380 => 41,
    7381 => 41,
    7382 => 41,
    7383 => 41,
    7384 => 41,
    7385 => 41,
    7386 => 41,
    7387 => 41,
    7388 => 41,
    7389 => 41,
    7390 => 41,
    7391 => 41,
    7392 => 41,
    7393 => 41,
    7394 => 41,
    7395 => 41,
    7396 => 41,
    7397 => 41,
    7398 => 41,
    7399 => 41,
    7400 => 41,
    7401 => 41,
    7402 => 41,
    7403 => 41,
    7404 => 41,
    7405 => 41,
    7406 => 41,
    7407 => 41,
    7408 => 41,
    7409 => 41,
    7410 => 41,
    7411 => 41,
    7412 => 41,
    7413 => 41,
    7414 => 41,
    7415 => 41,
    7416 => 41,
    7417 => 41,
    7418 => 41,
    7419 => 41,
    7420 => 41,
    7421 => 41,
    7422 => 41,
    7423 => 41,
    7424 => 41,
    7425 => 41,
    7426 => 41,
    7427 => 41,
    7428 => 41,
    7429 => 41,
    7430 => 41,
    7431 => 41,
    7432 => 41,
    7433 => 41,
    7434 => 41,
    7435 => 41,
    7436 => 41,
    7437 => 41,
    7438 => 41,
    7439 => 41,
    7440 => 41,
    7441 => 41,
    7442 => 41,
    7443 => 41,
    7444 => 41,
    7445 => 41,
    7446 => 41,
    7447 => 41,
    7448 => 41,
    7449 => 41,
    7450 => 41,
    7451 => 41,
    7452 => 41,
    7453 => 41,
    7454 => 41,
    7455 => 41,
    7456 => 41,
    7457 => 41,
    7458 => 41,
    7459 => 41,
    7460 => 41,
    7461 => 41,
    7462 => 41,
    7463 => 41,
    7464 => 41,
    7465 => 41,
    7466 => 41,
    7467 => 41,
    7468 => 41,
    7469 => 41,
    7470 => 41,
    7471 => 41,
    7472 => 41,
    7473 => 41,
    7474 => 41,
    7475 => 41,
    7476 => 41,
    7477 => 41,
    7478 => 41,
    7479 => 41,
    7480 => 41,
    7481 => 41,
    7482 => 41,
    7483 => 41,
    7484 => 41,
    7485 => 41,
    7486 => 41,
    7487 => 41,
    7488 => 41,
    7489 => 41,
    7490 => 41,
    7491 => 41,
    7492 => 41,
    7493 => 41,
    7494 => 41,
    7495 => 41,
    7496 => 41,
    7497 => 41,
    7498 => 41,
    7499 => 41,
    7500 => 41,
    7501 => 42,
    7502 => 42,
    7503 => 42,
    7504 => 42,
    7505 => 42,
    7506 => 42,
    7507 => 42,
    7508 => 42,
    7509 => 42,
    7510 => 42,
    7511 => 42,
    7512 => 42,
    7513 => 42,
    7514 => 42,
    7515 => 42,
    7516 => 42,
    7517 => 42,
    7518 => 42,
    7519 => 42,
    7520 => 42,
    7521 => 42,
    7522 => 42,
    7523 => 42,
    7524 => 42,
    7525 => 42,
    7526 => 42,
    7527 => 42,
    7528 => 42,
    7529 => 42,
    7530 => 42,
    7531 => 42,
    7532 => 42,
    7533 => 42,
    7534 => 42,
    7535 => 42,
    7536 => 42,
    7537 => 42,
    7538 => 42,
    7539 => 42,
    7540 => 42,
    7541 => 42,
    7542 => 42,
    7543 => 42,
    7544 => 42,
    7545 => 42,
    7546 => 42,
    7547 => 42,
    7548 => 42,
    7549 => 42,
    7550 => 42,
    7551 => 42,
    7552 => 42,
    7553 => 42,
    7554 => 42,
    7555 => 42,
    7556 => 42,
    7557 => 42,
    7558 => 42,
    7559 => 42,
    7560 => 42,
    7561 => 42,
    7562 => 42,
    7563 => 42,
    7564 => 42,
    7565 => 42,
    7566 => 42,
    7567 => 42,
    7568 => 42,
    7569 => 42,
    7570 => 42,
    7571 => 42,
    7572 => 42,
    7573 => 42,
    7574 => 42,
    7575 => 42,
    7576 => 42,
    7577 => 42,
    7578 => 42,
    7579 => 42,
    7580 => 42,
    7581 => 42,
    7582 => 42,
    7583 => 42,
    7584 => 42,
    7585 => 42,
    7586 => 42,
    7587 => 42,
    7588 => 42,
    7589 => 42,
    7590 => 42,
    7591 => 42,
    7592 => 42,
    7593 => 42,
    7594 => 42,
    7595 => 42,
    7596 => 42,
    7597 => 42,
    7598 => 42,
    7599 => 42,
    7600 => 42,
    7601 => 42,
    7602 => 42,
    7603 => 42,
    7604 => 42,
    7605 => 42,
    7606 => 42,
    7607 => 42,
    7608 => 42,
    7609 => 42,
    7610 => 42,
    7611 => 42,
    7612 => 42,
    7613 => 42,
    7614 => 42,
    7615 => 42,
    7616 => 42,
    7617 => 42,
    7618 => 42,
    7619 => 42,
    7620 => 42,
    7621 => 42,
    7622 => 42,
    7623 => 42,
    7624 => 42,
    7625 => 42,
    7626 => 42,
    7627 => 42,
    7628 => 42,
    7629 => 42,
    7630 => 42,
    7631 => 42,
    7632 => 42,
    7633 => 42,
    7634 => 42,
    7635 => 42,
    7636 => 42,
    7637 => 42,
    7638 => 42,
    7639 => 42,
    7640 => 42,
    7641 => 42,
    7642 => 42,
    7643 => 42,
    7644 => 42,
    7645 => 42,
    7646 => 42,
    7647 => 42,
    7648 => 42,
    7649 => 42,
    7650 => 42,
    7651 => 42,
    7652 => 42,
    7653 => 42,
    7654 => 42,
    7655 => 42,
    7656 => 42,
    7657 => 42,
    7658 => 42,
    7659 => 42,
    7660 => 42,
    7661 => 42,
    7662 => 42,
    7663 => 42,
    7664 => 42,
    7665 => 42,
    7666 => 42,
    7667 => 42,
    7668 => 42,
    7669 => 42,
    7670 => 42,
    7671 => 42,
    7672 => 42,
    7673 => 42,
    7674 => 42,
    7675 => 42,
    7676 => 42,
    7677 => 42,
    7678 => 42,
    7679 => 42,
    7680 => 42,
    7681 => 42,
    7682 => 42,
    7683 => 42,
    7684 => 42,
    7685 => 42,
    7686 => 42,
    7687 => 42,
    7688 => 42,
    7689 => 42,
    7690 => 42,
    7691 => 42,
    7692 => 42,
    7693 => 42,
    7694 => 42,
    7695 => 42,
    7696 => 42,
    7697 => 42,
    7698 => 42,
    7699 => 42,
    7700 => 42,
    7701 => 42,
    7702 => 42,
    7703 => 42,
    7704 => 42,
    7705 => 42,
    7706 => 42,
    7707 => 42,
    7708 => 42,
    7709 => 42,
    7710 => 42,
    7711 => 42,
    7712 => 42,
    7713 => 42,
    7714 => 42,
    7715 => 42,
    7716 => 42,
    7717 => 42,
    7718 => 42,
    7719 => 42,
    7720 => 42,
    7721 => 42,
    7722 => 42,
    7723 => 43,
    7724 => 43,
    7725 => 43,
    7726 => 43,
    7727 => 43,
    7728 => 43,
    7729 => 43,
    7730 => 43,
    7731 => 43,
    7732 => 43,
    7733 => 43,
    7734 => 43,
    7735 => 43,
    7736 => 43,
    7737 => 43,
    7738 => 43,
    7739 => 43,
    7740 => 43,
    7741 => 43,
    7742 => 43,
    7743 => 43,
    7744 => 43,
    7745 => 43,
    7746 => 43,
    7747 => 43,
    7748 => 43,
    7749 => 43,
    7750 => 43,
    7751 => 43,
    7752 => 43,
    7753 => 43,
    7754 => 43,
    7755 => 43,
    7756 => 43,
    7757 => 43,
    7758 => 43,
    7759 => 43,
    7760 => 43,
    7761 => 43,
    7762 => 43,
    7763 => 43,
    7764 => 43,
    7765 => 43,
    7766 => 43,
    7767 => 43,
    7768 => 43,
    7769 => 43,
    7770 => 43,
    7771 => 43,
    7772 => 43,
    7773 => 43,
    7774 => 43,
    7775 => 43,
    7776 => 43,
    7777 => 43,
    7778 => 43,
    7779 => 43,
    7780 => 43,
    7781 => 43,
    7782 => 43,
    7783 => 43,
    7784 => 43,
    7785 => 43,
    7786 => 43,
    7787 => 43,
    7788 => 43,
    7789 => 43,
    7790 => 43,
    7791 => 43,
    7792 => 43,
    7793 => 43,
    7794 => 43,
    7795 => 43,
    7796 => 43,
    7797 => 43,
    7798 => 43,
    7799 => 43,
    7800 => 43,
    7801 => 43,
    7802 => 43,
    7803 => 43,
    7804 => 43,
    7805 => 43,
    7806 => 43,
    7807 => 43,
    7808 => 43,
    7809 => 43,
    7810 => 43,
    7811 => 43,
    7812 => 43,
    7813 => 43,
    7814 => 43,
    7815 => 43,
    7816 => 43,
    7817 => 43,
    7818 => 43,
    7819 => 43,
    7820 => 43,
    7821 => 43,
    7822 => 43,
    7823 => 43,
    7824 => 43,
    7825 => 43,
    7826 => 43,
    7827 => 43,
    7828 => 43,
    7829 => 43,
    7830 => 43,
    7831 => 43,
    7832 => 43,
    7833 => 43,
    7834 => 43,
    7835 => 43,
    7836 => 43,
    7837 => 43,
    7838 => 43,
    7839 => 43,
    7840 => 43,
    7841 => 43,
    7842 => 43,
    7843 => 43,
    7844 => 43,
    7845 => 43,
    7846 => 43,
    7847 => 43,
    7848 => 43,
    7849 => 43,
    7850 => 43,
    7851 => 43,
    7852 => 43,
    7853 => 43,
    7854 => 43,
    7855 => 43,
    7856 => 43,
    7857 => 43,
    7858 => 43,
    7859 => 43,
    7860 => 43,
    7861 => 43,
    7862 => 43,
    7863 => 43,
    7864 => 43,
    7865 => 43,
    7866 => 43,
    7867 => 43,
    7868 => 43,
    7869 => 43,
    7870 => 43,
    7871 => 43,
    7872 => 43,
    7873 => 43,
    7874 => 43,
    7875 => 43,
    7876 => 43,
    7877 => 43,
    7878 => 43,
    7879 => 43,
    7880 => 43,
    7881 => 43,
    7882 => 43,
    7883 => 43,
    7884 => 43,
    7885 => 43,
    7886 => 43,
    7887 => 43,
    7888 => 43,
    7889 => 43,
    7890 => 43,
    7891 => 43,
    7892 => 43,
    7893 => 43,
    7894 => 43,
    7895 => 43,
    7896 => 43,
    7897 => 43,
    7898 => 43,
    7899 => 43,
    7900 => 43,
    7901 => 43,
    7902 => 43,
    7903 => 43,
    7904 => 43,
    7905 => 43,
    7906 => 43,
    7907 => 43,
    7908 => 43,
    7909 => 43,
    7910 => 43,
    7911 => 43,
    7912 => 43,
    7913 => 43,
    7914 => 43,
    7915 => 43,
    7916 => 43,
    7917 => 43,
    7918 => 43,
    7919 => 43,
    7920 => 43,
    7921 => 43,
    7922 => 43,
    7923 => 43,
    7924 => 43,
    7925 => 43,
    7926 => 43,
    7927 => 43,
    7928 => 43,
    7929 => 43,
    7930 => 43,
    7931 => 43,
    7932 => 43,
    7933 => 43,
    7934 => 43,
    7935 => 43,
    7936 => 43,
    7937 => 43,
    7938 => 43,
    7939 => 43,
    7940 => 43,
    7941 => 43,
    7942 => 43,
    7943 => 43,
    7944 => 43,
    7945 => 43,
    7946 => 43,
    7947 => 43,
    7948 => 43,
    7949 => 43,
    7950 => 44,
    7951 => 44,
    7952 => 44,
    7953 => 44,
    7954 => 44,
    7955 => 44,
    7956 => 44,
    7957 => 44,
    7958 => 44,
    7959 => 44,
    7960 => 44,
    7961 => 44,
    7962 => 44,
    7963 => 44,
    7964 => 44,
    7965 => 44,
    7966 => 44,
    7967 => 44,
    7968 => 44,
    7969 => 44,
    7970 => 44,
    7971 => 44,
    7972 => 44,
    7973 => 44,
    7974 => 44,
    7975 => 44,
    7976 => 44,
    7977 => 44,
    7978 => 44,
    7979 => 44,
    7980 => 44,
    7981 => 44,
    7982 => 44,
    7983 => 44,
    7984 => 44,
    7985 => 44,
    7986 => 44,
    7987 => 44,
    7988 => 44,
    7989 => 44,
    7990 => 44,
    7991 => 44,
    7992 => 44,
    7993 => 44,
    7994 => 44,
    7995 => 44,
    7996 => 44,
    7997 => 44,
    7998 => 44,
    7999 => 44,
    8000 => 44,
    8001 => 44,
    8002 => 44,
    8003 => 44,
    8004 => 44,
    8005 => 44,
    8006 => 44,
    8007 => 44,
    8008 => 44,
    8009 => 44,
    8010 => 44,
    8011 => 44,
    8012 => 44,
    8013 => 44,
    8014 => 44,
    8015 => 44,
    8016 => 44,
    8017 => 44,
    8018 => 44,
    8019 => 44,
    8020 => 44,
    8021 => 44,
    8022 => 44,
    8023 => 44,
    8024 => 44,
    8025 => 44,
    8026 => 44,
    8027 => 44,
    8028 => 44,
    8029 => 44,
    8030 => 44,
    8031 => 44,
    8032 => 44,
    8033 => 44,
    8034 => 44,
    8035 => 44,
    8036 => 44,
    8037 => 44,
    8038 => 44,
    8039 => 44,
    8040 => 44,
    8041 => 44,
    8042 => 44,
    8043 => 44,
    8044 => 44,
    8045 => 44,
    8046 => 44,
    8047 => 44,
    8048 => 44,
    8049 => 44,
    8050 => 44,
    8051 => 44,
    8052 => 44,
    8053 => 44,
    8054 => 44,
    8055 => 44,
    8056 => 44,
    8057 => 44,
    8058 => 44,
    8059 => 44,
    8060 => 44,
    8061 => 44,
    8062 => 44,
    8063 => 44,
    8064 => 44,
    8065 => 44,
    8066 => 44,
    8067 => 44,
    8068 => 44,
    8069 => 44,
    8070 => 44,
    8071 => 44,
    8072 => 44,
    8073 => 44,
    8074 => 44,
    8075 => 44,
    8076 => 44,
    8077 => 44,
    8078 => 44,
    8079 => 44,
    8080 => 44,
    8081 => 44,
    8082 => 44,
    8083 => 44,
    8084 => 44,
    8085 => 44,
    8086 => 44,
    8087 => 44,
    8088 => 44,
    8089 => 44,
    8090 => 44,
    8091 => 44,
    8092 => 44,
    8093 => 44,
    8094 => 44,
    8095 => 44,
    8096 => 44,
    8097 => 44,
    8098 => 44,
    8099 => 44,
    8100 => 44,
    8101 => 44,
    8102 => 44,
    8103 => 44,
    8104 => 44,
    8105 => 44,
    8106 => 44,
    8107 => 44,
    8108 => 44,
    8109 => 44,
    8110 => 44,
    8111 => 44,
    8112 => 44,
    8113 => 44,
    8114 => 44,
    8115 => 44,
    8116 => 44,
    8117 => 44,
    8118 => 44,
    8119 => 44,
    8120 => 44,
    8121 => 44,
    8122 => 44,
    8123 => 44,
    8124 => 44,
    8125 => 44,
    8126 => 44,
    8127 => 44,
    8128 => 44,
    8129 => 44,
    8130 => 44,
    8131 => 44,
    8132 => 44,
    8133 => 44,
    8134 => 44,
    8135 => 44,
    8136 => 44,
    8137 => 44,
    8138 => 44,
    8139 => 44,
    8140 => 44,
    8141 => 44,
    8142 => 44,
    8143 => 44,
    8144 => 44,
    8145 => 44,
    8146 => 44,
    8147 => 44,
    8148 => 44,
    8149 => 44,
    8150 => 44,
    8151 => 44,
    8152 => 44,
    8153 => 44,
    8154 => 44,
    8155 => 44,
    8156 => 44,
    8157 => 44,
    8158 => 44,
    8159 => 44,
    8160 => 44,
    8161 => 44,
    8162 => 44,
    8163 => 44,
    8164 => 44,
    8165 => 44,
    8166 => 44,
    8167 => 44,
    8168 => 44,
    8169 => 44,
    8170 => 44,
    8171 => 44,
    8172 => 44,
    8173 => 44,
    8174 => 44,
    8175 => 44,
    8176 => 44,
    8177 => 44,
    8178 => 44,
    8179 => 44,
    8180 => 44,
    8181 => 45,
    8182 => 45,
    8183 => 45,
    8184 => 45,
    8185 => 45,
    8186 => 45,
    8187 => 45,
    8188 => 45,
    8189 => 45,
    8190 => 45,
    8191 => 45,
    8192 => 45,
    8193 => 45,
    8194 => 45,
    8195 => 45,
    8196 => 45,
    8197 => 45,
    8198 => 45,
    8199 => 45,
    8200 => 45,
    8201 => 45,
    8202 => 45,
    8203 => 45,
    8204 => 45,
    8205 => 45,
    8206 => 45,
    8207 => 45,
    8208 => 45,
    8209 => 45,
    8210 => 45,
    8211 => 45,
    8212 => 45,
    8213 => 45,
    8214 => 45,
    8215 => 45,
    8216 => 45,
    8217 => 45,
    8218 => 45,
    8219 => 45,
    8220 => 45,
    8221 => 45,
    8222 => 45,
    8223 => 45,
    8224 => 45,
    8225 => 45,
    8226 => 45,
    8227 => 45,
    8228 => 45,
    8229 => 45,
    8230 => 45,
    8231 => 45,
    8232 => 45,
    8233 => 45,
    8234 => 45,
    8235 => 45,
    8236 => 45,
    8237 => 45,
    8238 => 45,
    8239 => 45,
    8240 => 45,
    8241 => 45,
    8242 => 45,
    8243 => 45,
    8244 => 45,
    8245 => 45,
    8246 => 45,
    8247 => 45,
    8248 => 45,
    8249 => 45,
    8250 => 45,
    8251 => 45,
    8252 => 45,
    8253 => 45,
    8254 => 45,
    8255 => 45,
    8256 => 45,
    8257 => 45,
    8258 => 45,
    8259 => 45,
    8260 => 45,
    8261 => 45,
    8262 => 45,
    8263 => 45,
    8264 => 45,
    8265 => 45,
    8266 => 45,
    8267 => 45,
    8268 => 45,
    8269 => 45,
    8270 => 45,
    8271 => 45,
    8272 => 45,
    8273 => 45,
    8274 => 45,
    8275 => 45,
    8276 => 45,
    8277 => 45,
    8278 => 45,
    8279 => 45,
    8280 => 45,
    8281 => 45,
    8282 => 45,
    8283 => 45,
    8284 => 45,
    8285 => 45,
    8286 => 45,
    8287 => 45,
    8288 => 45,
    8289 => 45,
    8290 => 45,
    8291 => 45,
    8292 => 45,
    8293 => 45,
    8294 => 45,
    8295 => 45,
    8296 => 45,
    8297 => 45,
    8298 => 45,
    8299 => 45,
    8300 => 45,
    8301 => 45,
    8302 => 45,
    8303 => 45,
    8304 => 45,
    8305 => 45,
    8306 => 45,
    8307 => 45,
    8308 => 45,
    8309 => 45,
    8310 => 45,
    8311 => 45,
    8312 => 45,
    8313 => 45,
    8314 => 45,
    8315 => 45,
    8316 => 45,
    8317 => 45,
    8318 => 45,
    8319 => 45,
    8320 => 45,
    8321 => 45,
    8322 => 45,
    8323 => 45,
    8324 => 45,
    8325 => 45,
    8326 => 45,
    8327 => 45,
    8328 => 45,
    8329 => 45,
    8330 => 45,
    8331 => 45,
    8332 => 45,
    8333 => 45,
    8334 => 45,
    8335 => 45,
    8336 => 45,
    8337 => 45,
    8338 => 45,
    8339 => 45,
    8340 => 45,
    8341 => 45,
    8342 => 45,
    8343 => 45,
    8344 => 45,
    8345 => 45,
    8346 => 45,
    8347 => 45,
    8348 => 45,
    8349 => 45,
    8350 => 45,
    8351 => 45,
    8352 => 45,
    8353 => 45,
    8354 => 45,
    8355 => 45,
    8356 => 45,
    8357 => 45,
    8358 => 45,
    8359 => 45,
    8360 => 45,
    8361 => 45,
    8362 => 45,
    8363 => 45,
    8364 => 45,
    8365 => 45,
    8366 => 45,
    8367 => 45,
    8368 => 45,
    8369 => 45,
    8370 => 45,
    8371 => 45,
    8372 => 45,
    8373 => 45,
    8374 => 45,
    8375 => 45,
    8376 => 45,
    8377 => 45,
    8378 => 45,
    8379 => 45,
    8380 => 45,
    8381 => 45,
    8382 => 45,
    8383 => 45,
    8384 => 45,
    8385 => 45,
    8386 => 45,
    8387 => 45,
    8388 => 45,
    8389 => 45,
    8390 => 45,
    8391 => 45,
    8392 => 45,
    8393 => 45,
    8394 => 45,
    8395 => 45,
    8396 => 45,
    8397 => 45,
    8398 => 45,
    8399 => 45,
    8400 => 45,
    8401 => 45,
    8402 => 45,
    8403 => 45,
    8404 => 45,
    8405 => 45,
    8406 => 45,
    8407 => 45,
    8408 => 45,
    8409 => 45,
    8410 => 45,
    8411 => 45,
    8412 => 45,
    8413 => 45,
    8414 => 45,
    8415 => 45,
    8416 => 45,
    8417 => 45,
    8418 => 46,
    8419 => 46,
    8420 => 46,
    8421 => 46,
    8422 => 46,
    8423 => 46,
    8424 => 46,
    8425 => 46,
    8426 => 46,
    8427 => 46,
    8428 => 46,
    8429 => 46,
    8430 => 46,
    8431 => 46,
    8432 => 46,
    8433 => 46,
    8434 => 46,
    8435 => 46,
    8436 => 46,
    8437 => 46,
    8438 => 46,
    8439 => 46,
    8440 => 46,
    8441 => 46,
    8442 => 46,
    8443 => 46,
    8444 => 46,
    8445 => 46,
    8446 => 46,
    8447 => 46,
    8448 => 46,
    8449 => 46,
    8450 => 46,
    8451 => 46,
    8452 => 46,
    8453 => 46,
    8454 => 46,
    8455 => 46,
    8456 => 46,
    8457 => 46,
    8458 => 46,
    8459 => 46,
    8460 => 46,
    8461 => 46,
    8462 => 46,
    8463 => 46,
    8464 => 46,
    8465 => 46,
    8466 => 46,
    8467 => 46,
    8468 => 46,
    8469 => 46,
    8470 => 46,
    8471 => 46,
    8472 => 46,
    8473 => 46,
    8474 => 46,
    8475 => 46,
    8476 => 46,
    8477 => 46,
    8478 => 46,
    8479 => 46,
    8480 => 46,
    8481 => 46,
    8482 => 46,
    8483 => 46,
    8484 => 46,
    8485 => 46,
    8486 => 46,
    8487 => 46,
    8488 => 46,
    8489 => 46,
    8490 => 46,
    8491 => 46,
    8492 => 46,
    8493 => 46,
    8494 => 46,
    8495 => 46,
    8496 => 46,
    8497 => 46,
    8498 => 46,
    8499 => 46,
    8500 => 46,
    8501 => 46,
    8502 => 46,
    8503 => 46,
    8504 => 46,
    8505 => 46,
    8506 => 46,
    8507 => 46,
    8508 => 46,
    8509 => 46,
    8510 => 46,
    8511 => 46,
    8512 => 46,
    8513 => 46,
    8514 => 46,
    8515 => 46,
    8516 => 46,
    8517 => 46,
    8518 => 46,
    8519 => 46,
    8520 => 46,
    8521 => 46,
    8522 => 46,
    8523 => 46,
    8524 => 46,
    8525 => 46,
    8526 => 46,
    8527 => 46,
    8528 => 46,
    8529 => 46,
    8530 => 46,
    8531 => 46,
    8532 => 46,
    8533 => 46,
    8534 => 46,
    8535 => 46,
    8536 => 46,
    8537 => 46,
    8538 => 46,
    8539 => 46,
    8540 => 46,
    8541 => 46,
    8542 => 46,
    8543 => 46,
    8544 => 46,
    8545 => 46,
    8546 => 46,
    8547 => 46,
    8548 => 46,
    8549 => 46,
    8550 => 46,
    8551 => 46,
    8552 => 46,
    8553 => 46,
    8554 => 46,
    8555 => 46,
    8556 => 46,
    8557 => 46,
    8558 => 46,
    8559 => 46,
    8560 => 46,
    8561 => 46,
    8562 => 46,
    8563 => 46,
    8564 => 46,
    8565 => 46,
    8566 => 46,
    8567 => 46,
    8568 => 46,
    8569 => 46,
    8570 => 46,
    8571 => 46,
    8572 => 46,
    8573 => 46,
    8574 => 46,
    8575 => 46,
    8576 => 46,
    8577 => 46,
    8578 => 46,
    8579 => 46,
    8580 => 46,
    8581 => 46,
    8582 => 46,
    8583 => 46,
    8584 => 46,
    8585 => 46,
    8586 => 46,
    8587 => 46,
    8588 => 46,
    8589 => 46,
    8590 => 46,
    8591 => 46,
    8592 => 46,
    8593 => 46,
    8594 => 46,
    8595 => 46,
    8596 => 46,
    8597 => 46,
    8598 => 46,
    8599 => 46,
    8600 => 46,
    8601 => 46,
    8602 => 46,
    8603 => 46,
    8604 => 46,
    8605 => 46,
    8606 => 46,
    8607 => 46,
    8608 => 46,
    8609 => 46,
    8610 => 46,
    8611 => 46,
    8612 => 46,
    8613 => 46,
    8614 => 46,
    8615 => 46,
    8616 => 46,
    8617 => 46,
    8618 => 46,
    8619 => 46,
    8620 => 46,
    8621 => 46,
    8622 => 46,
    8623 => 46,
    8624 => 46,
    8625 => 46,
    8626 => 46,
    8627 => 46,
    8628 => 46,
    8629 => 46,
    8630 => 46,
    8631 => 46,
    8632 => 46,
    8633 => 46,
    8634 => 46,
    8635 => 46,
    8636 => 46,
    8637 => 46,
    8638 => 46,
    8639 => 46,
    8640 => 46,
    8641 => 46,
    8642 => 46,
    8643 => 46,
    8644 => 46,
    8645 => 46,
    8646 => 46,
    8647 => 46,
    8648 => 46,
    8649 => 46,
    8650 => 46,
    8651 => 46,
    8652 => 46,
    8653 => 46,
    8654 => 46,
    8655 => 46,
    8656 => 46,
    8657 => 46,
    8658 => 46,
    8659 => 46,
    8660 => 47,
    8661 => 47,
    8662 => 47,
    8663 => 47,
    8664 => 47,
    8665 => 47,
    8666 => 47,
    8667 => 47,
    8668 => 47,
    8669 => 47,
    8670 => 47,
    8671 => 47,
    8672 => 47,
    8673 => 47,
    8674 => 47,
    8675 => 47,
    8676 => 47,
    8677 => 47,
    8678 => 47,
    8679 => 47,
    8680 => 47,
    8681 => 47,
    8682 => 47,
    8683 => 47,
    8684 => 47,
    8685 => 47,
    8686 => 47,
    8687 => 47,
    8688 => 47,
    8689 => 47,
    8690 => 47,
    8691 => 47,
    8692 => 47,
    8693 => 47,
    8694 => 47,
    8695 => 47,
    8696 => 47,
    8697 => 47,
    8698 => 47,
    8699 => 47,
    8700 => 47,
    8701 => 47,
    8702 => 47,
    8703 => 47,
    8704 => 47,
    8705 => 47,
    8706 => 47,
    8707 => 47,
    8708 => 47,
    8709 => 47,
    8710 => 47,
    8711 => 47,
    8712 => 47,
    8713 => 47,
    8714 => 47,
    8715 => 47,
    8716 => 47,
    8717 => 47,
    8718 => 47,
    8719 => 47,
    8720 => 47,
    8721 => 47,
    8722 => 47,
    8723 => 47,
    8724 => 47,
    8725 => 47,
    8726 => 47,
    8727 => 47,
    8728 => 47,
    8729 => 47,
    8730 => 47,
    8731 => 47,
    8732 => 47,
    8733 => 47,
    8734 => 47,
    8735 => 47,
    8736 => 47,
    8737 => 47,
    8738 => 47,
    8739 => 47,
    8740 => 47,
    8741 => 47,
    8742 => 47,
    8743 => 47,
    8744 => 47,
    8745 => 47,
    8746 => 47,
    8747 => 47,
    8748 => 47,
    8749 => 47,
    8750 => 47,
    8751 => 47,
    8752 => 47,
    8753 => 47,
    8754 => 47,
    8755 => 47,
    8756 => 47,
    8757 => 47,
    8758 => 47,
    8759 => 47,
    8760 => 47,
    8761 => 47,
    8762 => 47,
    8763 => 47,
    8764 => 47,
    8765 => 47,
    8766 => 47,
    8767 => 47,
    8768 => 47,
    8769 => 47,
    8770 => 47,
    8771 => 47,
    8772 => 47,
    8773 => 47,
    8774 => 47,
    8775 => 47,
    8776 => 47,
    8777 => 47,
    8778 => 47,
    8779 => 47,
    8780 => 47,
    8781 => 47,
    8782 => 47,
    8783 => 47,
    8784 => 47,
    8785 => 47,
    8786 => 47,
    8787 => 47,
    8788 => 47,
    8789 => 47,
    8790 => 47,
    8791 => 47,
    8792 => 47,
    8793 => 47,
    8794 => 47,
    8795 => 47,
    8796 => 47,
    8797 => 47,
    8798 => 47,
    8799 => 47,
    8800 => 47,
    8801 => 47,
    8802 => 47,
    8803 => 47,
    8804 => 47,
    8805 => 47,
    8806 => 47,
    8807 => 47,
    8808 => 47,
    8809 => 47,
    8810 => 47,
    8811 => 47,
    8812 => 47,
    8813 => 47,
    8814 => 47,
    8815 => 47,
    8816 => 47,
    8817 => 47,
    8818 => 47,
    8819 => 47,
    8820 => 47,
    8821 => 47,
    8822 => 47,
    8823 => 47,
    8824 => 47,
    8825 => 47,
    8826 => 47,
    8827 => 47,
    8828 => 47,
    8829 => 47,
    8830 => 47,
    8831 => 47,
    8832 => 47,
    8833 => 47,
    8834 => 47,
    8835 => 47,
    8836 => 47,
    8837 => 47,
    8838 => 47,
    8839 => 47,
    8840 => 47,
    8841 => 47,
    8842 => 47,
    8843 => 47,
    8844 => 47,
    8845 => 47,
    8846 => 47,
    8847 => 47,
    8848 => 47,
    8849 => 47,
    8850 => 47,
    8851 => 47,
    8852 => 47,
    8853 => 47,
    8854 => 47,
    8855 => 47,
    8856 => 47,
    8857 => 47,
    8858 => 47,
    8859 => 47,
    8860 => 47,
    8861 => 47,
    8862 => 47,
    8863 => 47,
    8864 => 47,
    8865 => 47,
    8866 => 47,
    8867 => 47,
    8868 => 47,
    8869 => 47,
    8870 => 47,
    8871 => 47,
    8872 => 47,
    8873 => 47,
    8874 => 47,
    8875 => 47,
    8876 => 47,
    8877 => 47,
    8878 => 47,
    8879 => 47,
    8880 => 47,
    8881 => 47,
    8882 => 47,
    8883 => 47,
    8884 => 47,
    8885 => 47,
    8886 => 47,
    8887 => 47,
    8888 => 47,
    8889 => 47,
    8890 => 47,
    8891 => 47,
    8892 => 47,
    8893 => 47,
    8894 => 47,
    8895 => 47,
    8896 => 47,
    8897 => 47,
    8898 => 47,
    8899 => 47,
    8900 => 47,
    8901 => 47,
    8902 => 47,
    8903 => 47,
    8904 => 47,
    8905 => 47,
    8906 => 47,
    8907 => 47,
    8908 => 47,
    8909 => 48,
    8910 => 48,
    8911 => 48,
    8912 => 48,
    8913 => 48,
    8914 => 48,
    8915 => 48,
    8916 => 48,
    8917 => 48,
    8918 => 48,
    8919 => 48,
    8920 => 48,
    8921 => 48,
    8922 => 48,
    8923 => 48,
    8924 => 48,
    8925 => 48,
    8926 => 48,
    8927 => 48,
    8928 => 48,
    8929 => 48,
    8930 => 48,
    8931 => 48,
    8932 => 48,
    8933 => 48,
    8934 => 48,
    8935 => 48,
    8936 => 48,
    8937 => 48,
    8938 => 48,
    8939 => 48,
    8940 => 48,
    8941 => 48,
    8942 => 48,
    8943 => 48,
    8944 => 48,
    8945 => 48,
    8946 => 48,
    8947 => 48,
    8948 => 48,
    8949 => 48,
    8950 => 48,
    8951 => 48,
    8952 => 48,
    8953 => 48,
    8954 => 48,
    8955 => 48,
    8956 => 48,
    8957 => 48,
    8958 => 48,
    8959 => 48,
    8960 => 48,
    8961 => 48,
    8962 => 48,
    8963 => 48,
    8964 => 48,
    8965 => 48,
    8966 => 48,
    8967 => 48,
    8968 => 48,
    8969 => 48,
    8970 => 48,
    8971 => 48,
    8972 => 48,
    8973 => 48,
    8974 => 48,
    8975 => 48,
    8976 => 48,
    8977 => 48,
    8978 => 48,
    8979 => 48,
    8980 => 48,
    8981 => 48,
    8982 => 48,
    8983 => 48,
    8984 => 48,
    8985 => 48,
    8986 => 48,
    8987 => 48,
    8988 => 48,
    8989 => 48,
    8990 => 48,
    8991 => 48,
    8992 => 48,
    8993 => 48,
    8994 => 48,
    8995 => 48,
    8996 => 48,
    8997 => 48,
    8998 => 48,
    8999 => 48,
    9000 => 48,
    9001 => 48,
    9002 => 48,
    9003 => 48,
    9004 => 48,
    9005 => 48,
    9006 => 48,
    9007 => 48,
    9008 => 48,
    9009 => 48,
    9010 => 48,
    9011 => 48,
    9012 => 48,
    9013 => 48,
    9014 => 48,
    9015 => 48,
    9016 => 48,
    9017 => 48,
    9018 => 48,
    9019 => 48,
    9020 => 48,
    9021 => 48,
    9022 => 48,
    9023 => 48,
    9024 => 48,
    9025 => 48,
    9026 => 48,
    9027 => 48,
    9028 => 48,
    9029 => 48,
    9030 => 48,
    9031 => 48,
    9032 => 48,
    9033 => 48,
    9034 => 48,
    9035 => 48,
    9036 => 48,
    9037 => 48,
    9038 => 48,
    9039 => 48,
    9040 => 48,
    9041 => 48,
    9042 => 48,
    9043 => 48,
    9044 => 48,
    9045 => 48,
    9046 => 48,
    9047 => 48,
    9048 => 48,
    9049 => 48,
    9050 => 48,
    9051 => 48,
    9052 => 48,
    9053 => 48,
    9054 => 48,
    9055 => 48,
    9056 => 48,
    9057 => 48,
    9058 => 48,
    9059 => 48,
    9060 => 48,
    9061 => 48,
    9062 => 48,
    9063 => 48,
    9064 => 48,
    9065 => 48,
    9066 => 48,
    9067 => 48,
    9068 => 48,
    9069 => 48,
    9070 => 48,
    9071 => 48,
    9072 => 48,
    9073 => 48,
    9074 => 48,
    9075 => 48,
    9076 => 48,
    9077 => 48,
    9078 => 48,
    9079 => 48,
    9080 => 48,
    9081 => 48,
    9082 => 48,
    9083 => 48,
    9084 => 48,
    9085 => 48,
    9086 => 48,
    9087 => 48,
    9088 => 48,
    9089 => 48,
    9090 => 48,
    9091 => 48,
    9092 => 48,
    9093 => 48,
    9094 => 48,
    9095 => 48,
    9096 => 48,
    9097 => 48,
    9098 => 48,
    9099 => 48,
    9100 => 48,
    9101 => 48,
    9102 => 48,
    9103 => 48,
    9104 => 48,
    9105 => 48,
    9106 => 48,
    9107 => 48,
    9108 => 48,
    9109 => 48,
    9110 => 48,
    9111 => 48,
    9112 => 48,
    9113 => 48,
    9114 => 48,
    9115 => 48,
    9116 => 48,
    9117 => 48,
    9118 => 48,
    9119 => 48,
    9120 => 48,
    9121 => 48,
    9122 => 48,
    9123 => 48,
    9124 => 48,
    9125 => 48,
    9126 => 48,
    9127 => 48,
    9128 => 48,
    9129 => 48,
    9130 => 48,
    9131 => 48,
    9132 => 48,
    9133 => 48,
    9134 => 48,
    9135 => 48,
    9136 => 48,
    9137 => 48,
    9138 => 48,
    9139 => 48,
    9140 => 48,
    9141 => 48,
    9142 => 48,
    9143 => 48,
    9144 => 48,
    9145 => 48,
    9146 => 48,
    9147 => 48,
    9148 => 48,
    9149 => 48,
    9150 => 48,
    9151 => 48,
    9152 => 48,
    9153 => 48,
    9154 => 48,
    9155 => 48,
    9156 => 48,
    9157 => 48,
    9158 => 48,
    9159 => 48,
    9160 => 48,
    9161 => 48,
    9162 => 48,
    9163 => 48,
    9164 => 48,
    9165 => 49,
    9166 => 49,
    9167 => 49,
    9168 => 49,
    9169 => 49,
    9170 => 49,
    9171 => 49,
    9172 => 49,
    9173 => 49,
    9174 => 49,
    9175 => 49,
    9176 => 49,
    9177 => 49,
    9178 => 49,
    9179 => 49,
    9180 => 49,
    9181 => 49,
    9182 => 49,
    9183 => 49,
    9184 => 49,
    9185 => 49,
    9186 => 49,
    9187 => 49,
    9188 => 49,
    9189 => 49,
    9190 => 49,
    9191 => 49,
    9192 => 49,
    9193 => 49,
    9194 => 49,
    9195 => 49,
    9196 => 49,
    9197 => 49,
    9198 => 49,
    9199 => 49,
    9200 => 49,
    9201 => 49,
    9202 => 49,
    9203 => 49,
    9204 => 49,
    9205 => 49,
    9206 => 49,
    9207 => 49,
    9208 => 49,
    9209 => 49,
    9210 => 49,
    9211 => 49,
    9212 => 49,
    9213 => 49,
    9214 => 49,
    9215 => 49,
    9216 => 49,
    9217 => 49,
    9218 => 49,
    9219 => 49,
    9220 => 49,
    9221 => 49,
    9222 => 49,
    9223 => 49,
    9224 => 49,
    9225 => 49,
    9226 => 49,
    9227 => 49,
    9228 => 49,
    9229 => 49,
    9230 => 49,
    9231 => 49,
    9232 => 49,
    9233 => 49,
    9234 => 49,
    9235 => 49,
    9236 => 49,
    9237 => 49,
    9238 => 49,
    9239 => 49,
    9240 => 49,
    9241 => 49,
    9242 => 49,
    9243 => 49,
    9244 => 49,
    9245 => 49,
    9246 => 49,
    9247 => 49,
    9248 => 49,
    9249 => 49,
    9250 => 49,
    9251 => 49,
    9252 => 49,
    9253 => 49,
    9254 => 49,
    9255 => 49,
    9256 => 49,
    9257 => 49,
    9258 => 49,
    9259 => 49,
    9260 => 49,
    9261 => 49,
    9262 => 49,
    9263 => 49,
    9264 => 49,
    9265 => 49,
    9266 => 49,
    9267 => 49,
    9268 => 49,
    9269 => 49,
    9270 => 49,
    9271 => 49,
    9272 => 49,
    9273 => 49,
    9274 => 49,
    9275 => 49,
    9276 => 49,
    9277 => 49,
    9278 => 49,
    9279 => 49,
    9280 => 49,
    9281 => 49,
    9282 => 49,
    9283 => 49,
    9284 => 49,
    9285 => 49,
    9286 => 49,
    9287 => 49,
    9288 => 49,
    9289 => 49,
    9290 => 49,
    9291 => 49,
    9292 => 49,
    9293 => 49,
    9294 => 49,
    9295 => 49,
    9296 => 49,
    9297 => 49,
    9298 => 49,
    9299 => 49,
    9300 => 49,
    9301 => 49,
    9302 => 49,
    9303 => 49,
    9304 => 49,
    9305 => 49,
    9306 => 49,
    9307 => 49,
    9308 => 49,
    9309 => 49,
    9310 => 49,
    9311 => 49,
    9312 => 49,
    9313 => 49,
    9314 => 49,
    9315 => 49,
    9316 => 49,
    9317 => 49,
    9318 => 49,
    9319 => 49,
    9320 => 49,
    9321 => 49,
    9322 => 49,
    9323 => 49,
    9324 => 49,
    9325 => 49,
    9326 => 49,
    9327 => 49,
    9328 => 49,
    9329 => 49,
    9330 => 49,
    9331 => 49,
    9332 => 49,
    9333 => 49,
    9334 => 49,
    9335 => 49,
    9336 => 49,
    9337 => 49,
    9338 => 49,
    9339 => 49,
    9340 => 49,
    9341 => 49,
    9342 => 49,
    9343 => 49,
    9344 => 49,
    9345 => 49,
    9346 => 49,
    9347 => 49,
    9348 => 49,
    9349 => 49,
    9350 => 49,
    9351 => 49,
    9352 => 49,
    9353 => 49,
    9354 => 49,
    9355 => 49,
    9356 => 49,
    9357 => 49,
    9358 => 49,
    9359 => 49,
    9360 => 49,
    9361 => 49,
    9362 => 49,
    9363 => 49,
    9364 => 49,
    9365 => 49,
    9366 => 49,
    9367 => 49,
    9368 => 49,
    9369 => 49,
    9370 => 49,
    9371 => 49,
    9372 => 49,
    9373 => 49,
    9374 => 49,
    9375 => 49,
    9376 => 49,
    9377 => 49,
    9378 => 49,
    9379 => 49,
    9380 => 49,
    9381 => 49,
    9382 => 49,
    9383 => 49,
    9384 => 49,
    9385 => 49,
    9386 => 49,
    9387 => 49,
    9388 => 49,
    9389 => 49,
    9390 => 49,
    9391 => 49,
    9392 => 49,
    9393 => 49,
    9394 => 49,
    9395 => 49,
    9396 => 49,
    9397 => 49,
    9398 => 49,
    9399 => 49,
    9400 => 49,
    9401 => 49,
    9402 => 49,
    9403 => 49,
    9404 => 49,
    9405 => 49,
    9406 => 49,
    9407 => 49,
    9408 => 49,
    9409 => 49,
    9410 => 49,
    9411 => 49,
    9412 => 49,
    9413 => 49,
    9414 => 49,
    9415 => 49,
    9416 => 49,
    9417 => 49,
    9418 => 49,
    9419 => 49,
    9420 => 49,
    9421 => 49,
    9422 => 49,
    9423 => 49,
    9424 => 49,
    9425 => 49,
    9426 => 49,
    9427 => 49,
    9428 => 50,
    9429 => 50,
    9430 => 50,
    9431 => 50,
    9432 => 50,
    9433 => 50,
    9434 => 50,
    9435 => 50,
    9436 => 50,
    9437 => 50,
    9438 => 50,
    9439 => 50,
    9440 => 50,
    9441 => 50,
    9442 => 50,
    9443 => 50,
    9444 => 50,
    9445 => 50,
    9446 => 50,
    9447 => 50,
    9448 => 50,
    9449 => 50,
    9450 => 50,
    9451 => 50,
    9452 => 50,
    9453 => 50,
    9454 => 50,
    9455 => 50,
    9456 => 50,
    9457 => 50,
    9458 => 50,
    9459 => 50,
    9460 => 50,
    9461 => 50,
    9462 => 50,
    9463 => 50,
    9464 => 50,
    9465 => 50,
    9466 => 50,
    9467 => 50,
    9468 => 50,
    9469 => 50,
    9470 => 50,
    9471 => 50,
    9472 => 50,
    9473 => 50,
    9474 => 50,
    9475 => 50,
    9476 => 50,
    9477 => 50,
    9478 => 50,
    9479 => 50,
    9480 => 50,
    9481 => 50,
    9482 => 50,
    9483 => 50,
    9484 => 50,
    9485 => 50,
    9486 => 50,
    9487 => 50,
    9488 => 50,
    9489 => 50,
    9490 => 50,
    9491 => 50,
    9492 => 50,
    9493 => 50,
    9494 => 50,
    9495 => 50,
    9496 => 50,
    9497 => 50,
    9498 => 50,
    9499 => 50,
    9500 => 50,
    9501 => 50,
    9502 => 50,
    9503 => 50,
    9504 => 50,
    9505 => 50,
    9506 => 50,
    9507 => 50,
    9508 => 50,
    9509 => 50,
    9510 => 50,
    9511 => 50,
    9512 => 50,
    9513 => 50,
    9514 => 50,
    9515 => 50,
    9516 => 50,
    9517 => 50,
    9518 => 50,
    9519 => 50,
    9520 => 50,
    9521 => 50,
    9522 => 50,
    9523 => 50,
    9524 => 50,
    9525 => 50,
    9526 => 50,
    9527 => 50,
    9528 => 50,
    9529 => 50,
    9530 => 50,
    9531 => 50,
    9532 => 50,
    9533 => 50,
    9534 => 50,
    9535 => 50,
    9536 => 50,
    9537 => 50,
    9538 => 50,
    9539 => 50,
    9540 => 50,
    9541 => 50,
    9542 => 50,
    9543 => 50,
    9544 => 50,
    9545 => 50,
    9546 => 50,
    9547 => 50,
    9548 => 50,
    9549 => 50,
    9550 => 50,
    9551 => 50,
    9552 => 50,
    9553 => 50,
    9554 => 50,
    9555 => 50,
    9556 => 50,
    9557 => 50,
    9558 => 50,
    9559 => 50,
    9560 => 50,
    9561 => 50,
    9562 => 50,
    9563 => 50,
    9564 => 50,
    9565 => 50,
    9566 => 50,
    9567 => 50,
    9568 => 50,
    9569 => 50,
    9570 => 50,
    9571 => 50,
    9572 => 50,
    9573 => 50,
    9574 => 50,
    9575 => 50,
    9576 => 50,
    9577 => 50,
    9578 => 50,
    9579 => 50,
    9580 => 50,
    9581 => 50,
    9582 => 50,
    9583 => 50,
    9584 => 50,
    9585 => 50,
    9586 => 50,
    9587 => 50,
    9588 => 50,
    9589 => 50,
    9590 => 50,
    9591 => 50,
    9592 => 50,
    9593 => 50,
    9594 => 50,
    9595 => 50,
    9596 => 50,
    9597 => 50,
    9598 => 50,
    9599 => 50,
    9600 => 50,
    9601 => 50,
    9602 => 50,
    9603 => 50,
    9604 => 50,
    9605 => 50,
    9606 => 50,
    9607 => 50,
    9608 => 50,
    9609 => 50,
    9610 => 50,
    9611 => 50,
    9612 => 50,
    9613 => 50,
    9614 => 50,
    9615 => 50,
    9616 => 50,
    9617 => 50,
    9618 => 50,
    9619 => 50,
    9620 => 50,
    9621 => 50,
    9622 => 50,
    9623 => 50,
    9624 => 50,
    9625 => 50,
    9626 => 50,
    9627 => 50,
    9628 => 50,
    9629 => 50,
    9630 => 50,
    9631 => 50,
    9632 => 50,
    9633 => 50,
    9634 => 50,
    9635 => 50,
    9636 => 50,
    9637 => 50,
    9638 => 50,
    9639 => 50,
    9640 => 50,
    9641 => 50,
    9642 => 50,
    9643 => 50,
    9644 => 50,
    9645 => 50,
    9646 => 50,
    9647 => 50,
    9648 => 50,
    9649 => 50,
    9650 => 50,
    9651 => 50,
    9652 => 50,
    9653 => 50,
    9654 => 50,
    9655 => 50,
    9656 => 50,
    9657 => 50,
    9658 => 50,
    9659 => 50,
    9660 => 50,
    9661 => 50,
    9662 => 50,
    9663 => 50,
    9664 => 50,
    9665 => 50,
    9666 => 50,
    9667 => 50,
    9668 => 50,
    9669 => 50,
    9670 => 50,
    9671 => 50,
    9672 => 50,
    9673 => 50,
    9674 => 50,
    9675 => 50,
    9676 => 50,
    9677 => 50,
    9678 => 50,
    9679 => 50,
    9680 => 50,
    9681 => 50,
    9682 => 50,
    9683 => 50,
    9684 => 50,
    9685 => 50,
    9686 => 50,
    9687 => 50,
    9688 => 50,
    9689 => 50,
    9690 => 50,
    9691 => 50,
    9692 => 50,
    9693 => 50,
    9694 => 50,
    9695 => 50,
    9696 => 50,
    9697 => 50,
    9698 => 50,
    9699 => 50,
    9700 => 51,
    9701 => 51,
    9702 => 51,
    9703 => 51,
    9704 => 51,
    9705 => 51,
    9706 => 51,
    9707 => 51,
    9708 => 51,
    9709 => 51,
    9710 => 51,
    9711 => 51,
    9712 => 51,
    9713 => 51,
    9714 => 51,
    9715 => 51,
    9716 => 51,
    9717 => 51,
    9718 => 51,
    9719 => 51,
    9720 => 51,
    9721 => 51,
    9722 => 51,
    9723 => 51,
    9724 => 51,
    9725 => 51,
    9726 => 51,
    9727 => 51,
    9728 => 51,
    9729 => 51,
    9730 => 51,
    9731 => 51,
    9732 => 51,
    9733 => 51,
    9734 => 51,
    9735 => 51,
    9736 => 51,
    9737 => 51,
    9738 => 51,
    9739 => 51,
    9740 => 51,
    9741 => 51,
    9742 => 51,
    9743 => 51,
    9744 => 51,
    9745 => 51,
    9746 => 51,
    9747 => 51,
    9748 => 51,
    9749 => 51,
    9750 => 51,
    9751 => 51,
    9752 => 51,
    9753 => 51,
    9754 => 51,
    9755 => 51,
    9756 => 51,
    9757 => 51,
    9758 => 51,
    9759 => 51,
    9760 => 51,
    9761 => 51,
    9762 => 51,
    9763 => 51,
    9764 => 51,
    9765 => 51,
    9766 => 51,
    9767 => 51,
    9768 => 51,
    9769 => 51,
    9770 => 51,
    9771 => 51,
    9772 => 51,
    9773 => 51,
    9774 => 51,
    9775 => 51,
    9776 => 51,
    9777 => 51,
    9778 => 51,
    9779 => 51,
    9780 => 51,
    9781 => 51,
    9782 => 51,
    9783 => 51,
    9784 => 51,
    9785 => 51,
    9786 => 51,
    9787 => 51,
    9788 => 51,
    9789 => 51,
    9790 => 51,
    9791 => 51,
    9792 => 51,
    9793 => 51,
    9794 => 51,
    9795 => 51,
    9796 => 51,
    9797 => 51,
    9798 => 51,
    9799 => 51,
    9800 => 51,
    9801 => 51,
    9802 => 51,
    9803 => 51,
    9804 => 51,
    9805 => 51,
    9806 => 51,
    9807 => 51,
    9808 => 51,
    9809 => 51,
    9810 => 51,
    9811 => 51,
    9812 => 51,
    9813 => 51,
    9814 => 51,
    9815 => 51,
    9816 => 51,
    9817 => 51,
    9818 => 51,
    9819 => 51,
    9820 => 51,
    9821 => 51,
    9822 => 51,
    9823 => 51,
    9824 => 51,
    9825 => 51,
    9826 => 51,
    9827 => 51,
    9828 => 51,
    9829 => 51,
    9830 => 51,
    9831 => 51,
    9832 => 51,
    9833 => 51,
    9834 => 51,
    9835 => 51,
    9836 => 51,
    9837 => 51,
    9838 => 51,
    9839 => 51,
    9840 => 51,
    9841 => 51,
    9842 => 51,
    9843 => 51,
    9844 => 51,
    9845 => 51,
    9846 => 51,
    9847 => 51,
    9848 => 51,
    9849 => 51,
    9850 => 51,
    9851 => 51,
    9852 => 51,
    9853 => 51,
    9854 => 51,
    9855 => 51,
    9856 => 51,
    9857 => 51,
    9858 => 51,
    9859 => 51,
    9860 => 51,
    9861 => 51,
    9862 => 51,
    9863 => 51,
    9864 => 51,
    9865 => 51,
    9866 => 51,
    9867 => 51,
    9868 => 51,
    9869 => 51,
    9870 => 51,
    9871 => 51,
    9872 => 51,
    9873 => 51,
    9874 => 51,
    9875 => 51,
    9876 => 51,
    9877 => 51,
    9878 => 51,
    9879 => 51,
    9880 => 51,
    9881 => 51,
    9882 => 51,
    9883 => 51,
    9884 => 51,
    9885 => 51,
    9886 => 51,
    9887 => 51,
    9888 => 51,
    9889 => 51,
    9890 => 51,
    9891 => 51,
    9892 => 51,
    9893 => 51,
    9894 => 51,
    9895 => 51,
    9896 => 51,
    9897 => 51,
    9898 => 51,
    9899 => 51,
    9900 => 51,
    9901 => 51,
    9902 => 51,
    9903 => 51,
    9904 => 51,
    9905 => 51,
    9906 => 51,
    9907 => 51,
    9908 => 51,
    9909 => 51,
    9910 => 51,
    9911 => 51,
    9912 => 51,
    9913 => 51,
    9914 => 51,
    9915 => 51,
    9916 => 51,
    9917 => 51,
    9918 => 51,
    9919 => 51,
    9920 => 51,
    9921 => 51,
    9922 => 51,
    9923 => 51,
    9924 => 51,
    9925 => 51,
    9926 => 51,
    9927 => 51,
    9928 => 51,
    9929 => 51,
    9930 => 51,
    9931 => 51,
    9932 => 51,
    9933 => 51,
    9934 => 51,
    9935 => 51,
    9936 => 51,
    9937 => 51,
    9938 => 51,
    9939 => 51,
    9940 => 51,
    9941 => 51,
    9942 => 51,
    9943 => 51,
    9944 => 51,
    9945 => 51,
    9946 => 51,
    9947 => 51,
    9948 => 51,
    9949 => 51,
    9950 => 51,
    9951 => 51,
    9952 => 51,
    9953 => 51,
    9954 => 51,
    9955 => 51,
    9956 => 51,
    9957 => 51,
    9958 => 51,
    9959 => 51,
    9960 => 51,
    9961 => 51,
    9962 => 51,
    9963 => 51,
    9964 => 51,
    9965 => 51,
    9966 => 51,
    9967 => 51,
    9968 => 51,
    9969 => 51,
    9970 => 51,
    9971 => 51,
    9972 => 51,
    9973 => 51,
    9974 => 51,
    9975 => 51,
    9976 => 51,
    9977 => 51,
    9978 => 51,
    9979 => 51,
    9980 => 51,
    9981 => 51,
    9982 => 52,
    9983 => 52,
    9984 => 52,
    9985 => 52,
    9986 => 52,
    9987 => 52,
    9988 => 52,
    9989 => 52,
    9990 => 52,
    9991 => 52,
    9992 => 52,
    9993 => 52,
    9994 => 52,
    9995 => 52,
    9996 => 52,
    9997 => 52,
    9998 => 52,
    9999 => 52,
    10000 => 52,
    10001 => 52,
    10002 => 52,
    10003 => 52,
    10004 => 52,
    10005 => 52,
    10006 => 52,
    10007 => 52,
    10008 => 52,
    10009 => 52,
    10010 => 52,
    10011 => 52,
    10012 => 52,
    10013 => 52,
    10014 => 52,
    10015 => 52,
    10016 => 52,
    10017 => 52,
    10018 => 52,
    10019 => 52,
    10020 => 52,
    10021 => 52,
    10022 => 52,
    10023 => 52,
    10024 => 52,
    10025 => 52,
    10026 => 52,
    10027 => 52,
    10028 => 52,
    10029 => 52,
    10030 => 52,
    10031 => 52,
    10032 => 52,
    10033 => 52,
    10034 => 52,
    10035 => 52,
    10036 => 52,
    10037 => 52,
    10038 => 52,
    10039 => 52,
    10040 => 52,
    10041 => 52,
    10042 => 52,
    10043 => 52,
    10044 => 52,
    10045 => 52,
    10046 => 52,
    10047 => 52,
    10048 => 52,
    10049 => 52,
    10050 => 52,
    10051 => 52,
    10052 => 52,
    10053 => 52,
    10054 => 52,
    10055 => 52,
    10056 => 52,
    10057 => 52,
    10058 => 52,
    10059 => 52,
    10060 => 52,
    10061 => 52,
    10062 => 52,
    10063 => 52,
    10064 => 52,
    10065 => 52,
    10066 => 52,
    10067 => 52,
    10068 => 52,
    10069 => 52,
    10070 => 52,
    10071 => 52,
    10072 => 52,
    10073 => 52,
    10074 => 52,
    10075 => 52,
    10076 => 52,
    10077 => 52,
    10078 => 52,
    10079 => 52,
    10080 => 52,
    10081 => 52,
    10082 => 52,
    10083 => 52,
    10084 => 52,
    10085 => 52,
    10086 => 52,
    10087 => 52,
    10088 => 52,
    10089 => 52,
    10090 => 52,
    10091 => 52,
    10092 => 52,
    10093 => 52,
    10094 => 52,
    10095 => 52,
    10096 => 52,
    10097 => 52,
    10098 => 52,
    10099 => 52,
    10100 => 52,
    10101 => 52,
    10102 => 52,
    10103 => 52,
    10104 => 52,
    10105 => 52,
    10106 => 52,
    10107 => 52,
    10108 => 52,
    10109 => 52,
    10110 => 52,
    10111 => 52,
    10112 => 52,
    10113 => 52,
    10114 => 52,
    10115 => 52,
    10116 => 52,
    10117 => 52,
    10118 => 52,
    10119 => 52,
    10120 => 52,
    10121 => 52,
    10122 => 52,
    10123 => 52,
    10124 => 52,
    10125 => 52,
    10126 => 52,
    10127 => 52,
    10128 => 52,
    10129 => 52,
    10130 => 52,
    10131 => 52,
    10132 => 52,
    10133 => 52,
    10134 => 52,
    10135 => 52,
    10136 => 52,
    10137 => 52,
    10138 => 52,
    10139 => 52,
    10140 => 52,
    10141 => 52,
    10142 => 52,
    10143 => 52,
    10144 => 52,
    10145 => 52,
    10146 => 52,
    10147 => 52,
    10148 => 52,
    10149 => 52,
    10150 => 52,
    10151 => 52,
    10152 => 52,
    10153 => 52,
    10154 => 52,
    10155 => 52,
    10156 => 52,
    10157 => 52,
    10158 => 52,
    10159 => 52,
    10160 => 52,
    10161 => 52,
    10162 => 52,
    10163 => 52,
    10164 => 52,
    10165 => 52,
    10166 => 52,
    10167 => 52,
    10168 => 52,
    10169 => 52,
    10170 => 52,
    10171 => 52,
    10172 => 52,
    10173 => 52,
    10174 => 52,
    10175 => 52,
    10176 => 52,
    10177 => 52,
    10178 => 52,
    10179 => 52,
    10180 => 52,
    10181 => 52,
    10182 => 52,
    10183 => 52,
    10184 => 52,
    10185 => 52,
    10186 => 52,
    10187 => 52,
    10188 => 52,
    10189 => 52,
    10190 => 52,
    10191 => 52,
    10192 => 52,
    10193 => 52,
    10194 => 52,
    10195 => 52,
    10196 => 52,
    10197 => 52,
    10198 => 52,
    10199 => 52,
    10200 => 52,
    10201 => 52,
    10202 => 52,
    10203 => 52,
    10204 => 52,
    10205 => 52,
    10206 => 52,
    10207 => 52,
    10208 => 52,
    10209 => 52,
    10210 => 52,
    10211 => 52,
    10212 => 52,
    10213 => 52,
    10214 => 52,
    10215 => 52,
    10216 => 52,
    10217 => 52,
    10218 => 52,
    10219 => 52,
    10220 => 52,
    10221 => 52,
    10222 => 52,
    10223 => 52,
    10224 => 52,
    10225 => 52,
    10226 => 52,
    10227 => 52,
    10228 => 52,
    10229 => 52,
    10230 => 52,
    10231 => 52,
    10232 => 52,
    10233 => 52,
    10234 => 52,
    10235 => 52,
    10236 => 52,
    10237 => 52,
    10238 => 52,
    10239 => 52,
    10240 => 52,
    10241 => 52,
    10242 => 52,
    10243 => 52,
    10244 => 52,
    10245 => 52,
    10246 => 52,
    10247 => 52,
    10248 => 52,
    10249 => 52,
    10250 => 52,
    10251 => 52,
    10252 => 52,
    10253 => 52,
    10254 => 52,
    10255 => 52,
    10256 => 52,
    10257 => 52,
    10258 => 52,
    10259 => 52,
    10260 => 52,
    10261 => 52,
    10262 => 52,
    10263 => 52,
    10264 => 52,
    10265 => 52,
    10266 => 52,
    10267 => 52,
    10268 => 52,
    10269 => 52,
    10270 => 52,
    10271 => 52,
    10272 => 52,
    10273 => 52,
    10274 => 52,
    10275 => 52,
    10276 => 53,
    10277 => 53,
    10278 => 53,
    10279 => 53,
    10280 => 53,
    10281 => 53,
    10282 => 53,
    10283 => 53,
    10284 => 53,
    10285 => 53,
    10286 => 53,
    10287 => 53,
    10288 => 53,
    10289 => 53,
    10290 => 53,
    10291 => 53,
    10292 => 53,
    10293 => 53,
    10294 => 53,
    10295 => 53,
    10296 => 53,
    10297 => 53,
    10298 => 53,
    10299 => 53,
    10300 => 53,
    10301 => 53,
    10302 => 53,
    10303 => 53,
    10304 => 53,
    10305 => 53,
    10306 => 53,
    10307 => 53,
    10308 => 53,
    10309 => 53,
    10310 => 53,
    10311 => 53,
    10312 => 53,
    10313 => 53,
    10314 => 53,
    10315 => 53,
    10316 => 53,
    10317 => 53,
    10318 => 53,
    10319 => 53,
    10320 => 53,
    10321 => 53,
    10322 => 53,
    10323 => 53,
    10324 => 53,
    10325 => 53,
    10326 => 53,
    10327 => 53,
    10328 => 53,
    10329 => 53,
    10330 => 53,
    10331 => 53,
    10332 => 53,
    10333 => 53,
    10334 => 53,
    10335 => 53,
    10336 => 53,
    10337 => 53,
    10338 => 53,
    10339 => 53,
    10340 => 53,
    10341 => 53,
    10342 => 53,
    10343 => 53,
    10344 => 53,
    10345 => 53,
    10346 => 53,
    10347 => 53,
    10348 => 53,
    10349 => 53,
    10350 => 53,
    10351 => 53,
    10352 => 53,
    10353 => 53,
    10354 => 53,
    10355 => 53,
    10356 => 53,
    10357 => 53,
    10358 => 53,
    10359 => 53,
    10360 => 53,
    10361 => 53,
    10362 => 53,
    10363 => 53,
    10364 => 53,
    10365 => 53,
    10366 => 53,
    10367 => 53,
    10368 => 53,
    10369 => 53,
    10370 => 53,
    10371 => 53,
    10372 => 53,
    10373 => 53,
    10374 => 53,
    10375 => 53,
    10376 => 53,
    10377 => 53,
    10378 => 53,
    10379 => 53,
    10380 => 53,
    10381 => 53,
    10382 => 53,
    10383 => 53,
    10384 => 53,
    10385 => 53,
    10386 => 53,
    10387 => 53,
    10388 => 53,
    10389 => 53,
    10390 => 53,
    10391 => 53,
    10392 => 53,
    10393 => 53,
    10394 => 53,
    10395 => 53,
    10396 => 53,
    10397 => 53,
    10398 => 53,
    10399 => 53,
    10400 => 53,
    10401 => 53,
    10402 => 53,
    10403 => 53,
    10404 => 53,
    10405 => 53,
    10406 => 53,
    10407 => 53,
    10408 => 53,
    10409 => 53,
    10410 => 53,
    10411 => 53,
    10412 => 53,
    10413 => 53,
    10414 => 53,
    10415 => 53,
    10416 => 53,
    10417 => 53,
    10418 => 53,
    10419 => 53,
    10420 => 53,
    10421 => 53,
    10422 => 53,
    10423 => 53,
    10424 => 53,
    10425 => 53,
    10426 => 53,
    10427 => 53,
    10428 => 53,
    10429 => 53,
    10430 => 53,
    10431 => 53,
    10432 => 53,
    10433 => 53,
    10434 => 53,
    10435 => 53,
    10436 => 53,
    10437 => 53,
    10438 => 53,
    10439 => 53,
    10440 => 53,
    10441 => 53,
    10442 => 53,
    10443 => 53,
    10444 => 53,
    10445 => 53,
    10446 => 53,
    10447 => 53,
    10448 => 53,
    10449 => 53,
    10450 => 53,
    10451 => 53,
    10452 => 53,
    10453 => 53,
    10454 => 53,
    10455 => 53,
    10456 => 53,
    10457 => 53,
    10458 => 53,
    10459 => 53,
    10460 => 53,
    10461 => 53,
    10462 => 53,
    10463 => 53,
    10464 => 53,
    10465 => 53,
    10466 => 53,
    10467 => 53,
    10468 => 53,
    10469 => 53,
    10470 => 53,
    10471 => 53,
    10472 => 53,
    10473 => 53,
    10474 => 53,
    10475 => 53,
    10476 => 53,
    10477 => 53,
    10478 => 53,
    10479 => 53,
    10480 => 53,
    10481 => 53,
    10482 => 53,
    10483 => 53,
    10484 => 53,
    10485 => 53,
    10486 => 53,
    10487 => 53,
    10488 => 53,
    10489 => 53,
    10490 => 53,
    10491 => 53,
    10492 => 53,
    10493 => 53,
    10494 => 53,
    10495 => 53,
    10496 => 53,
    10497 => 53,
    10498 => 53,
    10499 => 53,
    10500 => 53,
    10501 => 53,
    10502 => 53,
    10503 => 53,
    10504 => 53,
    10505 => 53,
    10506 => 53,
    10507 => 53,
    10508 => 53,
    10509 => 53,
    10510 => 53,
    10511 => 53,
    10512 => 53,
    10513 => 53,
    10514 => 53,
    10515 => 53,
    10516 => 53,
    10517 => 53,
    10518 => 53,
    10519 => 53,
    10520 => 53,
    10521 => 53,
    10522 => 53,
    10523 => 53,
    10524 => 53,
    10525 => 53,
    10526 => 53,
    10527 => 53,
    10528 => 53,
    10529 => 53,
    10530 => 53,
    10531 => 53,
    10532 => 53,
    10533 => 53,
    10534 => 53,
    10535 => 53,
    10536 => 53,
    10537 => 53,
    10538 => 53,
    10539 => 53,
    10540 => 53,
    10541 => 53,
    10542 => 53,
    10543 => 53,
    10544 => 53,
    10545 => 53,
    10546 => 53,
    10547 => 53,
    10548 => 53,
    10549 => 53,
    10550 => 53,
    10551 => 53,
    10552 => 53,
    10553 => 53,
    10554 => 53,
    10555 => 53,
    10556 => 53,
    10557 => 53,
    10558 => 53,
    10559 => 53,
    10560 => 53,
    10561 => 53,
    10562 => 53,
    10563 => 53,
    10564 => 53,
    10565 => 53,
    10566 => 53,
    10567 => 53,
    10568 => 53,
    10569 => 53,
    10570 => 53,
    10571 => 53,
    10572 => 53,
    10573 => 53,
    10574 => 53,
    10575 => 53,
    10576 => 53,
    10577 => 53,
    10578 => 53,
    10579 => 53,
    10580 => 53,
    10581 => 53,
    10582 => 54,
    10583 => 54,
    10584 => 54,
    10585 => 54,
    10586 => 54,
    10587 => 54,
    10588 => 54,
    10589 => 54,
    10590 => 54,
    10591 => 54,
    10592 => 54,
    10593 => 54,
    10594 => 54,
    10595 => 54,
    10596 => 54,
    10597 => 54,
    10598 => 54,
    10599 => 54,
    10600 => 54,
    10601 => 54,
    10602 => 54,
    10603 => 54,
    10604 => 54,
    10605 => 54,
    10606 => 54,
    10607 => 54,
    10608 => 54,
    10609 => 54,
    10610 => 54,
    10611 => 54,
    10612 => 54,
    10613 => 54,
    10614 => 54,
    10615 => 54,
    10616 => 54,
    10617 => 54,
    10618 => 54,
    10619 => 54,
    10620 => 54,
    10621 => 54,
    10622 => 54,
    10623 => 54,
    10624 => 54,
    10625 => 54,
    10626 => 54,
    10627 => 54,
    10628 => 54,
    10629 => 54,
    10630 => 54,
    10631 => 54,
    10632 => 54,
    10633 => 54,
    10634 => 54,
    10635 => 54,
    10636 => 54,
    10637 => 54,
    10638 => 54,
    10639 => 54,
    10640 => 54,
    10641 => 54,
    10642 => 54,
    10643 => 54,
    10644 => 54,
    10645 => 54,
    10646 => 54,
    10647 => 54,
    10648 => 54,
    10649 => 54,
    10650 => 54,
    10651 => 54,
    10652 => 54,
    10653 => 54,
    10654 => 54,
    10655 => 54,
    10656 => 54,
    10657 => 54,
    10658 => 54,
    10659 => 54,
    10660 => 54,
    10661 => 54,
    10662 => 54,
    10663 => 54,
    10664 => 54,
    10665 => 54,
    10666 => 54,
    10667 => 54,
    10668 => 54,
    10669 => 54,
    10670 => 54,
    10671 => 54,
    10672 => 54,
    10673 => 54,
    10674 => 54,
    10675 => 54,
    10676 => 54,
    10677 => 54,
    10678 => 54,
    10679 => 54,
    10680 => 54,
    10681 => 54,
    10682 => 54,
    10683 => 54,
    10684 => 54,
    10685 => 54,
    10686 => 54,
    10687 => 54,
    10688 => 54,
    10689 => 54,
    10690 => 54,
    10691 => 54,
    10692 => 54,
    10693 => 54,
    10694 => 54,
    10695 => 54,
    10696 => 54,
    10697 => 54,
    10698 => 54,
    10699 => 54,
    10700 => 54,
    10701 => 54,
    10702 => 54,
    10703 => 54,
    10704 => 54,
    10705 => 54,
    10706 => 54,
    10707 => 54,
    10708 => 54,
    10709 => 54,
    10710 => 54,
    10711 => 54,
    10712 => 54,
    10713 => 54,
    10714 => 54,
    10715 => 54,
    10716 => 54,
    10717 => 54,
    10718 => 54,
    10719 => 54,
    10720 => 54,
    10721 => 54,
    10722 => 54,
    10723 => 54,
    10724 => 54,
    10725 => 54,
    10726 => 54,
    10727 => 54,
    10728 => 54,
    10729 => 54,
    10730 => 54,
    10731 => 54,
    10732 => 54,
    10733 => 54,
    10734 => 54,
    10735 => 54,
    10736 => 54,
    10737 => 54,
    10738 => 54,
    10739 => 54,
    10740 => 54,
    10741 => 54,
    10742 => 54,
    10743 => 54,
    10744 => 54,
    10745 => 54,
    10746 => 54,
    10747 => 54,
    10748 => 54,
    10749 => 54,
    10750 => 54,
    10751 => 54,
    10752 => 54,
    10753 => 54,
    10754 => 54,
    10755 => 54,
    10756 => 54,
    10757 => 54,
    10758 => 54,
    10759 => 54,
    10760 => 54,
    10761 => 54,
    10762 => 54,
    10763 => 54,
    10764 => 54,
    10765 => 54,
    10766 => 54,
    10767 => 54,
    10768 => 54,
    10769 => 54,
    10770 => 54,
    10771 => 54,
    10772 => 54,
    10773 => 54,
    10774 => 54,
    10775 => 54,
    10776 => 54,
    10777 => 54,
    10778 => 54,
    10779 => 54,
    10780 => 54,
    10781 => 54,
    10782 => 54,
    10783 => 54,
    10784 => 54,
    10785 => 54,
    10786 => 54,
    10787 => 54,
    10788 => 54,
    10789 => 54,
    10790 => 54,
    10791 => 54,
    10792 => 54,
    10793 => 54,
    10794 => 54,
    10795 => 54,
    10796 => 54,
    10797 => 54,
    10798 => 54,
    10799 => 54,
    10800 => 54,
    10801 => 54,
    10802 => 54,
    10803 => 54,
    10804 => 54,
    10805 => 54,
    10806 => 54,
    10807 => 54,
    10808 => 54,
    10809 => 54,
    10810 => 54,
    10811 => 54,
    10812 => 54,
    10813 => 54,
    10814 => 54,
    10815 => 54,
    10816 => 54,
    10817 => 54,
    10818 => 54,
    10819 => 54,
    10820 => 54,
    10821 => 54,
    10822 => 54,
    10823 => 54,
    10824 => 54,
    10825 => 54,
    10826 => 54,
    10827 => 54,
    10828 => 54,
    10829 => 54,
    10830 => 54,
    10831 => 54,
    10832 => 54,
    10833 => 54,
    10834 => 54,
    10835 => 54,
    10836 => 54,
    10837 => 54,
    10838 => 54,
    10839 => 54,
    10840 => 54,
    10841 => 54,
    10842 => 54,
    10843 => 54,
    10844 => 54,
    10845 => 54,
    10846 => 54,
    10847 => 54,
    10848 => 54,
    10849 => 54,
    10850 => 54,
    10851 => 54,
    10852 => 54,
    10853 => 54,
    10854 => 54,
    10855 => 54,
    10856 => 54,
    10857 => 54,
    10858 => 54,
    10859 => 54,
    10860 => 54,
    10861 => 54,
    10862 => 54,
    10863 => 54,
    10864 => 54,
    10865 => 54,
    10866 => 54,
    10867 => 54,
    10868 => 54,
    10869 => 54,
    10870 => 54,
    10871 => 54,
    10872 => 54,
    10873 => 54,
    10874 => 54,
    10875 => 54,
    10876 => 54,
    10877 => 54,
    10878 => 54,
    10879 => 54,
    10880 => 54,
    10881 => 54,
    10882 => 54,
    10883 => 54,
    10884 => 54,
    10885 => 54,
    10886 => 54,
    10887 => 54,
    10888 => 54,
    10889 => 54,
    10890 => 54,
    10891 => 54,
    10892 => 54,
    10893 => 54,
    10894 => 54,
    10895 => 54,
    10896 => 54,
    10897 => 54,
    10898 => 54,
    10899 => 54,
    10900 => 54,
    10901 => 54,
    10902 => 54,
    10903 => 55,
    10904 => 55,
    10905 => 55,
    10906 => 55,
    10907 => 55,
    10908 => 55,
    10909 => 55,
    10910 => 55,
    10911 => 55,
    10912 => 55,
    10913 => 55,
    10914 => 55,
    10915 => 55,
    10916 => 55,
    10917 => 55,
    10918 => 55,
    10919 => 55,
    10920 => 55,
    10921 => 55,
    10922 => 55,
    10923 => 55,
    10924 => 55,
    10925 => 55,
    10926 => 55,
    10927 => 55,
    10928 => 55,
    10929 => 55,
    10930 => 55,
    10931 => 55,
    10932 => 55,
    10933 => 55,
    10934 => 55,
    10935 => 55,
    10936 => 55,
    10937 => 55,
    10938 => 55,
    10939 => 55,
    10940 => 55,
    10941 => 55,
    10942 => 55,
    10943 => 55,
    10944 => 55,
    10945 => 55,
    10946 => 55,
    10947 => 55,
    10948 => 55,
    10949 => 55,
    10950 => 55,
    10951 => 55,
    10952 => 55,
    10953 => 55,
    10954 => 55,
    10955 => 55,
    10956 => 55,
    10957 => 55,
    10958 => 55,
    10959 => 55,
    10960 => 55,
    10961 => 55,
    10962 => 55,
    10963 => 55,
    10964 => 55,
    10965 => 55,
    10966 => 55,
    10967 => 55,
    10968 => 55,
    10969 => 55,
    10970 => 55,
    10971 => 55,
    10972 => 55,
    10973 => 55,
    10974 => 55,
    10975 => 55,
    10976 => 55,
    10977 => 55,
    10978 => 55,
    10979 => 55,
    10980 => 55,
    10981 => 55,
    10982 => 55,
    10983 => 55,
    10984 => 55,
    10985 => 55,
    10986 => 55,
    10987 => 55,
    10988 => 55,
    10989 => 55,
    10990 => 55,
    10991 => 55,
    10992 => 55,
    10993 => 55,
    10994 => 55,
    10995 => 55,
    10996 => 55,
    10997 => 55,
    10998 => 55,
    10999 => 55,
    11000 => 55,
    11001 => 55,
    11002 => 55,
    11003 => 55,
    11004 => 55,
    11005 => 55,
    11006 => 55,
    11007 => 55,
    11008 => 55,
    11009 => 55,
    11010 => 55,
    11011 => 55,
    11012 => 55,
    11013 => 55,
    11014 => 55,
    11015 => 55,
    11016 => 55,
    11017 => 55,
    11018 => 55,
    11019 => 55,
    11020 => 55,
    11021 => 55,
    11022 => 55,
    11023 => 55,
    11024 => 55,
    11025 => 55,
    11026 => 55,
    11027 => 55,
    11028 => 55,
    11029 => 55,
    11030 => 55,
    11031 => 55,
    11032 => 55,
    11033 => 55,
    11034 => 55,
    11035 => 55,
    11036 => 55,
    11037 => 55,
    11038 => 55,
    11039 => 55,
    11040 => 55,
    11041 => 55,
    11042 => 55,
    11043 => 55,
    11044 => 55,
    11045 => 55,
    11046 => 55,
    11047 => 55,
    11048 => 55,
    11049 => 55,
    11050 => 55,
    11051 => 55,
    11052 => 55,
    11053 => 55,
    11054 => 55,
    11055 => 55,
    11056 => 55,
    11057 => 55,
    11058 => 55,
    11059 => 55,
    11060 => 55,
    11061 => 55,
    11062 => 55,
    11063 => 55,
    11064 => 55,
    11065 => 55,
    11066 => 55,
    11067 => 55,
    11068 => 55,
    11069 => 55,
    11070 => 55,
    11071 => 55,
    11072 => 55,
    11073 => 55,
    11074 => 55,
    11075 => 55,
    11076 => 55,
    11077 => 55,
    11078 => 55,
    11079 => 55,
    11080 => 55,
    11081 => 55,
    11082 => 55,
    11083 => 55,
    11084 => 55,
    11085 => 55,
    11086 => 55,
    11087 => 55,
    11088 => 55,
    11089 => 55,
    11090 => 55,
    11091 => 55,
    11092 => 55,
    11093 => 55,
    11094 => 55,
    11095 => 55,
    11096 => 55,
    11097 => 55,
    11098 => 55,
    11099 => 55,
    11100 => 55,
    11101 => 55,
    11102 => 55,
    11103 => 55,
    11104 => 55,
    11105 => 55,
    11106 => 55,
    11107 => 55,
    11108 => 55,
    11109 => 55,
    11110 => 55,
    11111 => 55,
    11112 => 55,
    11113 => 55,
    11114 => 55,
    11115 => 55,
    11116 => 55,
    11117 => 55,
    11118 => 55,
    11119 => 55,
    11120 => 55,
    11121 => 55,
    11122 => 55,
    11123 => 55,
    11124 => 55,
    11125 => 55,
    11126 => 55,
    11127 => 55,
    11128 => 55,
    11129 => 55,
    11130 => 55,
    11131 => 55,
    11132 => 55,
    11133 => 55,
    11134 => 55,
    11135 => 55,
    11136 => 55,
    11137 => 55,
    11138 => 55,
    11139 => 55,
    11140 => 55,
    11141 => 55,
    11142 => 55,
    11143 => 55,
    11144 => 55,
    11145 => 55,
    11146 => 55,
    11147 => 55,
    11148 => 55,
    11149 => 55,
    11150 => 55,
    11151 => 55,
    11152 => 55,
    11153 => 55,
    11154 => 55,
    11155 => 55,
    11156 => 55,
    11157 => 55,
    11158 => 55,
    11159 => 55,
    11160 => 55,
    11161 => 55,
    11162 => 55,
    11163 => 55,
    11164 => 55,
    11165 => 55,
    11166 => 55,
    11167 => 55,
    11168 => 55,
    11169 => 55,
    11170 => 55,
    11171 => 55,
    11172 => 55,
    11173 => 55,
    11174 => 55,
    11175 => 55,
    11176 => 55,
    11177 => 55,
    11178 => 55,
    11179 => 55,
    11180 => 55,
    11181 => 55,
    11182 => 55,
    11183 => 55,
    11184 => 55,
    11185 => 55,
    11186 => 55,
    11187 => 55,
    11188 => 55,
    11189 => 55,
    11190 => 55,
    11191 => 55,
    11192 => 55,
    11193 => 55,
    11194 => 55,
    11195 => 55,
    11196 => 55,
    11197 => 55,
    11198 => 55,
    11199 => 55,
    11200 => 55,
    11201 => 55,
    11202 => 55,
    11203 => 55,
    11204 => 55,
    11205 => 55,
    11206 => 55,
    11207 => 55,
    11208 => 55,
    11209 => 55,
    11210 => 55,
    11211 => 55,
    11212 => 55,
    11213 => 55,
    11214 => 55,
    11215 => 55,
    11216 => 55,
    11217 => 55,
    11218 => 55,
    11219 => 55,
    11220 => 55,
    11221 => 55,
    11222 => 55,
    11223 => 55,
    11224 => 55,
    11225 => 55,
    11226 => 55,
    11227 => 55,
    11228 => 55,
    11229 => 55,
    11230 => 55,
    11231 => 55,
    11232 => 55,
    11233 => 55,
    11234 => 55,
    11235 => 55,
    11236 => 55,
    11237 => 55,
    11238 => 55,
    11239 => 55,
    11240 => 55,
    11241 => 55,
    11242 => 55,
    11243 => 56,
    11244 => 56,
    11245 => 56,
    11246 => 56,
    11247 => 56,
    11248 => 56,
    11249 => 56,
    11250 => 56,
    11251 => 56,
    11252 => 56,
    11253 => 56,
    11254 => 56,
    11255 => 56,
    11256 => 56,
    11257 => 56,
    11258 => 56,
    11259 => 56,
    11260 => 56,
    11261 => 56,
    11262 => 56,
    11263 => 56,
    11264 => 56,
    11265 => 56,
    11266 => 56,
    11267 => 56,
    11268 => 56,
    11269 => 56,
    11270 => 56,
    11271 => 56,
    11272 => 56,
    11273 => 56,
    11274 => 56,
    11275 => 56,
    11276 => 56,
    11277 => 56,
    11278 => 56,
    11279 => 56,
    11280 => 56,
    11281 => 56,
    11282 => 56,
    11283 => 56,
    11284 => 56,
    11285 => 56,
    11286 => 56,
    11287 => 56,
    11288 => 56,
    11289 => 56,
    11290 => 56,
    11291 => 56,
    11292 => 56,
    11293 => 56,
    11294 => 56,
    11295 => 56,
    11296 => 56,
    11297 => 56,
    11298 => 56,
    11299 => 56,
    11300 => 56,
    11301 => 56,
    11302 => 56,
    11303 => 56,
    11304 => 56,
    11305 => 56,
    11306 => 56,
    11307 => 56,
    11308 => 56,
    11309 => 56,
    11310 => 56,
    11311 => 56,
    11312 => 56,
    11313 => 56,
    11314 => 56,
    11315 => 56,
    11316 => 56,
    11317 => 56,
    11318 => 56,
    11319 => 56,
    11320 => 56,
    11321 => 56,
    11322 => 56,
    11323 => 56,
    11324 => 56,
    11325 => 56,
    11326 => 56,
    11327 => 56,
    11328 => 56,
    11329 => 56,
    11330 => 56,
    11331 => 56,
    11332 => 56,
    11333 => 56,
    11334 => 56,
    11335 => 56,
    11336 => 56,
    11337 => 56,
    11338 => 56,
    11339 => 56,
    11340 => 56,
    11341 => 56,
    11342 => 56,
    11343 => 56,
    11344 => 56,
    11345 => 56,
    11346 => 56,
    11347 => 56,
    11348 => 56,
    11349 => 56,
    11350 => 56,
    11351 => 56,
    11352 => 56,
    11353 => 56,
    11354 => 56,
    11355 => 56,
    11356 => 56,
    11357 => 56,
    11358 => 56,
    11359 => 56,
    11360 => 56,
    11361 => 56,
    11362 => 56,
    11363 => 56,
    11364 => 56,
    11365 => 56,
    11366 => 56,
    11367 => 56,
    11368 => 56,
    11369 => 56,
    11370 => 56,
    11371 => 56,
    11372 => 56,
    11373 => 56,
    11374 => 56,
    11375 => 56,
    11376 => 56,
    11377 => 56,
    11378 => 56,
    11379 => 56,
    11380 => 56,
    11381 => 56,
    11382 => 56,
    11383 => 56,
    11384 => 56,
    11385 => 56,
    11386 => 56,
    11387 => 56,
    11388 => 56,
    11389 => 56,
    11390 => 56,
    11391 => 56,
    11392 => 56,
    11393 => 56,
    11394 => 56,
    11395 => 56,
    11396 => 56,
    11397 => 56,
    11398 => 56,
    11399 => 56,
    11400 => 56,
    11401 => 56,
    11402 => 56,
    11403 => 56,
    11404 => 56,
    11405 => 56,
    11406 => 56,
    11407 => 56,
    11408 => 56,
    11409 => 56,
    11410 => 56,
    11411 => 56,
    11412 => 56,
    11413 => 56,
    11414 => 56,
    11415 => 56,
    11416 => 56,
    11417 => 56,
    11418 => 56,
    11419 => 56,
    11420 => 56,
    11421 => 56,
    11422 => 56,
    11423 => 56,
    11424 => 56,
    11425 => 56,
    11426 => 56,
    11427 => 56,
    11428 => 56,
    11429 => 56,
    11430 => 56,
    11431 => 56,
    11432 => 56,
    11433 => 56,
    11434 => 56,
    11435 => 56,
    11436 => 56,
    11437 => 56,
    11438 => 56,
    11439 => 56,
    11440 => 56,
    11441 => 56,
    11442 => 56,
    11443 => 56,
    11444 => 56,
    11445 => 56,
    11446 => 56,
    11447 => 56,
    11448 => 56,
    11449 => 56,
    11450 => 56,
    11451 => 56,
    11452 => 56,
    11453 => 56,
    11454 => 56,
    11455 => 56,
    11456 => 56,
    11457 => 56,
    11458 => 56,
    11459 => 56,
    11460 => 56,
    11461 => 56,
    11462 => 56,
    11463 => 56,
    11464 => 56,
    11465 => 56,
    11466 => 56,
    11467 => 56,
    11468 => 56,
    11469 => 56,
    11470 => 56,
    11471 => 56,
    11472 => 56,
    11473 => 56,
    11474 => 56,
    11475 => 56,
    11476 => 56,
    11477 => 56,
    11478 => 56,
    11479 => 56,
    11480 => 56,
    11481 => 56,
    11482 => 56,
    11483 => 56,
    11484 => 56,
    11485 => 56,
    11486 => 56,
    11487 => 56,
    11488 => 56,
    11489 => 56,
    11490 => 56,
    11491 => 56,
    11492 => 56,
    11493 => 56,
    11494 => 56,
    11495 => 56,
    11496 => 56,
    11497 => 56,
    11498 => 56,
    11499 => 56,
    11500 => 56,
    11501 => 56,
    11502 => 56,
    11503 => 56,
    11504 => 56,
    11505 => 56,
    11506 => 56,
    11507 => 56,
    11508 => 56,
    11509 => 56,
    11510 => 56,
    11511 => 56,
    11512 => 56,
    11513 => 56,
    11514 => 56,
    11515 => 56,
    11516 => 56,
    11517 => 56,
    11518 => 56,
    11519 => 56,
    11520 => 56,
    11521 => 56,
    11522 => 56,
    11523 => 56,
    11524 => 56,
    11525 => 56,
    11526 => 56,
    11527 => 56,
    11528 => 56,
    11529 => 56,
    11530 => 56,
    11531 => 56,
    11532 => 56,
    11533 => 56,
    11534 => 56,
    11535 => 56,
    11536 => 56,
    11537 => 56,
    11538 => 56,
    11539 => 56,
    11540 => 56,
    11541 => 56,
    11542 => 56,
    11543 => 56,
    11544 => 56,
    11545 => 56,
    11546 => 56,
    11547 => 56,
    11548 => 56,
    11549 => 56,
    11550 => 56,
    11551 => 56,
    11552 => 56,
    11553 => 56,
    11554 => 56,
    11555 => 56,
    11556 => 56,
    11557 => 56,
    11558 => 56,
    11559 => 56,
    11560 => 56,
    11561 => 56,
    11562 => 56,
    11563 => 56,
    11564 => 56,
    11565 => 56,
    11566 => 56,
    11567 => 56,
    11568 => 56,
    11569 => 56,
    11570 => 56,
    11571 => 56,
    11572 => 56,
    11573 => 56,
    11574 => 56,
    11575 => 56,
    11576 => 56,
    11577 => 56,
    11578 => 56,
    11579 => 56,
    11580 => 56,
    11581 => 56,
    11582 => 56,
    11583 => 56,
    11584 => 56,
    11585 => 56,
    11586 => 56,
    11587 => 56,
    11588 => 56,
    11589 => 56,
    11590 => 56,
    11591 => 56,
    11592 => 56,
    11593 => 56,
    11594 => 56,
    11595 => 56,
    11596 => 56,
    11597 => 56,
    11598 => 56,
    11599 => 56,
    11600 => 56,
    11601 => 56,
    11602 => 56,
    11603 => 56,
    11604 => 56,
    11605 => 57,
    11606 => 57,
    11607 => 57,
    11608 => 57,
    11609 => 57,
    11610 => 57,
    11611 => 57,
    11612 => 57,
    11613 => 57,
    11614 => 57,
    11615 => 57,
    11616 => 57,
    11617 => 57,
    11618 => 57,
    11619 => 57,
    11620 => 57,
    11621 => 57,
    11622 => 57,
    11623 => 57,
    11624 => 57,
    11625 => 57,
    11626 => 57,
    11627 => 57,
    11628 => 57,
    11629 => 57,
    11630 => 57,
    11631 => 57,
    11632 => 57,
    11633 => 57,
    11634 => 57,
    11635 => 57,
    11636 => 57,
    11637 => 57,
    11638 => 57,
    11639 => 57,
    11640 => 57,
    11641 => 57,
    11642 => 57,
    11643 => 57,
    11644 => 57,
    11645 => 57,
    11646 => 57,
    11647 => 57,
    11648 => 57,
    11649 => 57,
    11650 => 57,
    11651 => 57,
    11652 => 57,
    11653 => 57,
    11654 => 57,
    11655 => 57,
    11656 => 57,
    11657 => 57,
    11658 => 57,
    11659 => 57,
    11660 => 57,
    11661 => 57,
    11662 => 57,
    11663 => 57,
    11664 => 57,
    11665 => 57,
    11666 => 57,
    11667 => 57,
    11668 => 57,
    11669 => 57,
    11670 => 57,
    11671 => 57,
    11672 => 57,
    11673 => 57,
    11674 => 57,
    11675 => 57,
    11676 => 57,
    11677 => 57,
    11678 => 57,
    11679 => 57,
    11680 => 57,
    11681 => 57,
    11682 => 57,
    11683 => 57,
    11684 => 57,
    11685 => 57,
    11686 => 57,
    11687 => 57,
    11688 => 57,
    11689 => 57,
    11690 => 57,
    11691 => 57,
    11692 => 57,
    11693 => 57,
    11694 => 57,
    11695 => 57,
    11696 => 57,
    11697 => 57,
    11698 => 57,
    11699 => 57,
    11700 => 57,
    11701 => 57,
    11702 => 57,
    11703 => 57,
    11704 => 57,
    11705 => 57,
    11706 => 57,
    11707 => 57,
    11708 => 57,
    11709 => 57,
    11710 => 57,
    11711 => 57,
    11712 => 57,
    11713 => 57,
    11714 => 57,
    11715 => 57,
    11716 => 57,
    11717 => 57,
    11718 => 57,
    11719 => 57,
    11720 => 57,
    11721 => 57,
    11722 => 57,
    11723 => 57,
    11724 => 57,
    11725 => 57,
    11726 => 57,
    11727 => 57,
    11728 => 57,
    11729 => 57,
    11730 => 57,
    11731 => 57,
    11732 => 57,
    11733 => 57,
    11734 => 57,
    11735 => 57,
    11736 => 57,
    11737 => 57,
    11738 => 57,
    11739 => 57,
    11740 => 57,
    11741 => 57,
    11742 => 57,
    11743 => 57,
    11744 => 57,
    11745 => 57,
    11746 => 57,
    11747 => 57,
    11748 => 57,
    11749 => 57,
    11750 => 57,
    11751 => 57,
    11752 => 57,
    11753 => 57,
    11754 => 57,
    11755 => 57,
    11756 => 57,
    11757 => 57,
    11758 => 57,
    11759 => 57,
    11760 => 57,
    11761 => 57,
    11762 => 57,
    11763 => 57,
    11764 => 57,
    11765 => 57,
    11766 => 57,
    11767 => 57,
    11768 => 57,
    11769 => 57,
    11770 => 57,
    11771 => 57,
    11772 => 57,
    11773 => 57,
    11774 => 57,
    11775 => 57,
    11776 => 57,
    11777 => 57,
    11778 => 57,
    11779 => 57,
    11780 => 57,
    11781 => 57,
    11782 => 57,
    11783 => 57,
    11784 => 57,
    11785 => 57,
    11786 => 57,
    11787 => 57,
    11788 => 57,
    11789 => 57,
    11790 => 57,
    11791 => 57,
    11792 => 57,
    11793 => 57,
    11794 => 57,
    11795 => 57,
    11796 => 57,
    11797 => 57,
    11798 => 57,
    11799 => 57,
    11800 => 57,
    11801 => 57,
    11802 => 57,
    11803 => 57,
    11804 => 57,
    11805 => 57,
    11806 => 57,
    11807 => 57,
    11808 => 57,
    11809 => 57,
    11810 => 57,
    11811 => 57,
    11812 => 57,
    11813 => 57,
    11814 => 57,
    11815 => 57,
    11816 => 57,
    11817 => 57,
    11818 => 57,
    11819 => 57,
    11820 => 57,
    11821 => 57,
    11822 => 57,
    11823 => 57,
    11824 => 57,
    11825 => 57,
    11826 => 57,
    11827 => 57,
    11828 => 57,
    11829 => 57,
    11830 => 57,
    11831 => 57,
    11832 => 57,
    11833 => 57,
    11834 => 57,
    11835 => 57,
    11836 => 57,
    11837 => 57,
    11838 => 57,
    11839 => 57,
    11840 => 57,
    11841 => 57,
    11842 => 57,
    11843 => 57,
    11844 => 57,
    11845 => 57,
    11846 => 57,
    11847 => 57,
    11848 => 57,
    11849 => 57,
    11850 => 57,
    11851 => 57,
    11852 => 57,
    11853 => 57,
    11854 => 57,
    11855 => 57,
    11856 => 57,
    11857 => 57,
    11858 => 57,
    11859 => 57,
    11860 => 57,
    11861 => 57,
    11862 => 57,
    11863 => 57,
    11864 => 57,
    11865 => 57,
    11866 => 57,
    11867 => 57,
    11868 => 57,
    11869 => 57,
    11870 => 57,
    11871 => 57,
    11872 => 57,
    11873 => 57,
    11874 => 57,
    11875 => 57,
    11876 => 57,
    11877 => 57,
    11878 => 57,
    11879 => 57,
    11880 => 57,
    11881 => 57,
    11882 => 57,
    11883 => 57,
    11884 => 57,
    11885 => 57,
    11886 => 57,
    11887 => 57,
    11888 => 57,
    11889 => 57,
    11890 => 57,
    11891 => 57,
    11892 => 57,
    11893 => 57,
    11894 => 57,
    11895 => 57,
    11896 => 57,
    11897 => 57,
    11898 => 57,
    11899 => 57,
    11900 => 57,
    11901 => 57,
    11902 => 57,
    11903 => 57,
    11904 => 57,
    11905 => 57,
    11906 => 57,
    11907 => 57,
    11908 => 57,
    11909 => 57,
    11910 => 57,
    11911 => 57,
    11912 => 57,
    11913 => 57,
    11914 => 57,
    11915 => 57,
    11916 => 57,
    11917 => 57,
    11918 => 57,
    11919 => 57,
    11920 => 57,
    11921 => 57,
    11922 => 57,
    11923 => 57,
    11924 => 57,
    11925 => 57,
    11926 => 57,
    11927 => 57,
    11928 => 57,
    11929 => 57,
    11930 => 57,
    11931 => 57,
    11932 => 57,
    11933 => 57,
    11934 => 57,
    11935 => 57,
    11936 => 57,
    11937 => 57,
    11938 => 57,
    11939 => 57,
    11940 => 57,
    11941 => 57,
    11942 => 57,
    11943 => 57,
    11944 => 57,
    11945 => 57,
    11946 => 57,
    11947 => 57,
    11948 => 57,
    11949 => 57,
    11950 => 57,
    11951 => 57,
    11952 => 57,
    11953 => 57,
    11954 => 57,
    11955 => 57,
    11956 => 57,
    11957 => 57,
    11958 => 57,
    11959 => 57,
    11960 => 57,
    11961 => 57,
    11962 => 57,
    11963 => 57,
    11964 => 57,
    11965 => 57,
    11966 => 57,
    11967 => 57,
    11968 => 57,
    11969 => 57,
    11970 => 57,
    11971 => 57,
    11972 => 57,
    11973 => 57,
    11974 => 57,
    11975 => 57,
    11976 => 57,
    11977 => 57,
    11978 => 57,
    11979 => 57,
    11980 => 57,
    11981 => 57,
    11982 => 57,
    11983 => 57,
    11984 => 57,
    11985 => 57,
    11986 => 57,
    11987 => 57,
    11988 => 57,
    11989 => 57,
    11990 => 57,
    11991 => 57,
    11992 => 57,
    11993 => 57,
    11994 => 58,
    11995 => 58,
    11996 => 58,
    11997 => 58,
    11998 => 58,
    11999 => 58,
    12000 => 58,
    12001 => 58,
    12002 => 58,
    12003 => 58,
    12004 => 58,
    12005 => 58,
    12006 => 58,
    12007 => 58,
    12008 => 58,
    12009 => 58,
    12010 => 58,
    12011 => 58,
    12012 => 58,
    12013 => 58,
    12014 => 58,
    12015 => 58,
    12016 => 58,
    12017 => 58,
    12018 => 58,
    12019 => 58,
    12020 => 58,
    12021 => 58,
    12022 => 58,
    12023 => 58,
    12024 => 58,
    12025 => 58,
    12026 => 58,
    12027 => 58,
    12028 => 58,
    12029 => 58,
    12030 => 58,
    12031 => 58,
    12032 => 58,
    12033 => 58,
    12034 => 58,
    12035 => 58,
    12036 => 58,
    12037 => 58,
    12038 => 58,
    12039 => 58,
    12040 => 58,
    12041 => 58,
    12042 => 58,
    12043 => 58,
    12044 => 58,
    12045 => 58,
    12046 => 58,
    12047 => 58,
    12048 => 58,
    12049 => 58,
    12050 => 58,
    12051 => 58,
    12052 => 58,
    12053 => 58,
    12054 => 58,
    12055 => 58,
    12056 => 58,
    12057 => 58,
    12058 => 58,
    12059 => 58,
    12060 => 58,
    12061 => 58,
    12062 => 58,
    12063 => 58,
    12064 => 58,
    12065 => 58,
    12066 => 58,
    12067 => 58,
    12068 => 58,
    12069 => 58,
    12070 => 58,
    12071 => 58,
    12072 => 58,
    12073 => 58,
    12074 => 58,
    12075 => 58,
    12076 => 58,
    12077 => 58,
    12078 => 58,
    12079 => 58,
    12080 => 58,
    12081 => 58,
    12082 => 58,
    12083 => 58,
    12084 => 58,
    12085 => 58,
    12086 => 58,
    12087 => 58,
    12088 => 58,
    12089 => 58,
    12090 => 58,
    12091 => 58,
    12092 => 58,
    12093 => 58,
    12094 => 58,
    12095 => 58,
    12096 => 58,
    12097 => 58,
    12098 => 58,
    12099 => 58,
    12100 => 58,
    12101 => 58,
    12102 => 58,
    12103 => 58,
    12104 => 58,
    12105 => 58,
    12106 => 58,
    12107 => 58,
    12108 => 58,
    12109 => 58,
    12110 => 58,
    12111 => 58,
    12112 => 58,
    12113 => 58,
    12114 => 58,
    12115 => 58,
    12116 => 58,
    12117 => 58,
    12118 => 58,
    12119 => 58,
    12120 => 58,
    12121 => 58,
    12122 => 58,
    12123 => 58,
    12124 => 58,
    12125 => 58,
    12126 => 58,
    12127 => 58,
    12128 => 58,
    12129 => 58,
    12130 => 58,
    12131 => 58,
    12132 => 58,
    12133 => 58,
    12134 => 58,
    12135 => 58,
    12136 => 58,
    12137 => 58,
    12138 => 58,
    12139 => 58,
    12140 => 58,
    12141 => 58,
    12142 => 58,
    12143 => 58,
    12144 => 58,
    12145 => 58,
    12146 => 58,
    12147 => 58,
    12148 => 58,
    12149 => 58,
    12150 => 58,
    12151 => 58,
    12152 => 58,
    12153 => 58,
    12154 => 58,
    12155 => 58,
    12156 => 58,
    12157 => 58,
    12158 => 58,
    12159 => 58,
    12160 => 58,
    12161 => 58,
    12162 => 58,
    12163 => 58,
    12164 => 58,
    12165 => 58,
    12166 => 58,
    12167 => 58,
    12168 => 58,
    12169 => 58,
    12170 => 58,
    12171 => 58,
    12172 => 58,
    12173 => 58,
    12174 => 58,
    12175 => 58,
    12176 => 58,
    12177 => 58,
    12178 => 58,
    12179 => 58,
    12180 => 58,
    12181 => 58,
    12182 => 58,
    12183 => 58,
    12184 => 58,
    12185 => 58,
    12186 => 58,
    12187 => 58,
    12188 => 58,
    12189 => 58,
    12190 => 58,
    12191 => 58,
    12192 => 58,
    12193 => 58,
    12194 => 58,
    12195 => 58,
    12196 => 58,
    12197 => 58,
    12198 => 58,
    12199 => 58,
    12200 => 58,
    12201 => 58,
    12202 => 58,
    12203 => 58,
    12204 => 58,
    12205 => 58,
    12206 => 58,
    12207 => 58,
    12208 => 58,
    12209 => 58,
    12210 => 58,
    12211 => 58,
    12212 => 58,
    12213 => 58,
    12214 => 58,
    12215 => 58,
    12216 => 58,
    12217 => 58,
    12218 => 58,
    12219 => 58,
    12220 => 58,
    12221 => 58,
    12222 => 58,
    12223 => 58,
    12224 => 58,
    12225 => 58,
    12226 => 58,
    12227 => 58,
    12228 => 58,
    12229 => 58,
    12230 => 58,
    12231 => 58,
    12232 => 58,
    12233 => 58,
    12234 => 58,
    12235 => 58,
    12236 => 58,
    12237 => 58,
    12238 => 58,
    12239 => 58,
    12240 => 58,
    12241 => 58,
    12242 => 58,
    12243 => 58,
    12244 => 58,
    12245 => 58,
    12246 => 58,
    12247 => 58,
    12248 => 58,
    12249 => 58,
    12250 => 58,
    12251 => 58,
    12252 => 58,
    12253 => 58,
    12254 => 58,
    12255 => 58,
    12256 => 58,
    12257 => 58,
    12258 => 58,
    12259 => 58,
    12260 => 58,
    12261 => 58,
    12262 => 58,
    12263 => 58,
    12264 => 58,
    12265 => 58,
    12266 => 58,
    12267 => 58,
    12268 => 58,
    12269 => 58,
    12270 => 58,
    12271 => 58,
    12272 => 58,
    12273 => 58,
    12274 => 58,
    12275 => 58,
    12276 => 58,
    12277 => 58,
    12278 => 58,
    12279 => 58,
    12280 => 58,
    12281 => 58,
    12282 => 58,
    12283 => 58,
    12284 => 58,
    12285 => 58,
    12286 => 58,
    12287 => 58,
    12288 => 58,
    12289 => 58,
    12290 => 58,
    12291 => 58,
    12292 => 58,
    12293 => 58,
    12294 => 58,
    12295 => 58,
    12296 => 58,
    12297 => 58,
    12298 => 58,
    12299 => 58,
    12300 => 58,
    12301 => 58,
    12302 => 58,
    12303 => 58,
    12304 => 58,
    12305 => 58,
    12306 => 58,
    12307 => 58,
    12308 => 58,
    12309 => 58,
    12310 => 58,
    12311 => 58,
    12312 => 58,
    12313 => 58,
    12314 => 58,
    12315 => 58,
    12316 => 58,
    12317 => 58,
    12318 => 58,
    12319 => 58,
    12320 => 58,
    12321 => 58,
    12322 => 58,
    12323 => 58,
    12324 => 58,
    12325 => 58,
    12326 => 58,
    12327 => 58,
    12328 => 58,
    12329 => 58,
    12330 => 58,
    12331 => 58,
    12332 => 58,
    12333 => 58,
    12334 => 58,
    12335 => 58,
    12336 => 58,
    12337 => 58,
    12338 => 58,
    12339 => 58,
    12340 => 58,
    12341 => 58,
    12342 => 58,
    12343 => 58,
    12344 => 58,
    12345 => 58,
    12346 => 58,
    12347 => 58,
    12348 => 58,
    12349 => 58,
    12350 => 58,
    12351 => 58,
    12352 => 58,
    12353 => 58,
    12354 => 58,
    12355 => 58,
    12356 => 58,
    12357 => 58,
    12358 => 58,
    12359 => 58,
    12360 => 58,
    12361 => 58,
    12362 => 58,
    12363 => 58,
    12364 => 58,
    12365 => 58,
    12366 => 58,
    12367 => 58,
    12368 => 58,
    12369 => 58,
    12370 => 58,
    12371 => 58,
    12372 => 58,
    12373 => 58,
    12374 => 58,
    12375 => 58,
    12376 => 58,
    12377 => 58,
    12378 => 58,
    12379 => 58,
    12380 => 58,
    12381 => 58,
    12382 => 58,
    12383 => 58,
    12384 => 58,
    12385 => 58,
    12386 => 58,
    12387 => 58,
    12388 => 58,
    12389 => 58,
    12390 => 58,
    12391 => 58,
    12392 => 58,
    12393 => 58,
    12394 => 58,
    12395 => 58,
    12396 => 58,
    12397 => 58,
    12398 => 58,
    12399 => 58,
    12400 => 58,
    12401 => 58,
    12402 => 58,
    12403 => 58,
    12404 => 58,
    12405 => 58,
    12406 => 58,
    12407 => 58,
    12408 => 58,
    12409 => 58,
    12410 => 58,
    12411 => 58,
    12412 => 58,
    12413 => 58,
    12414 => 58,
    12415 => 58,
    12416 => 58,
    12417 => 58,
    12418 => 59,
    12419 => 59,
    12420 => 59,
    12421 => 59,
    12422 => 59,
    12423 => 59,
    12424 => 59,
    12425 => 59,
    12426 => 59,
    12427 => 59,
    12428 => 59,
    12429 => 59,
    12430 => 59,
    12431 => 59,
    12432 => 59,
    12433 => 59,
    12434 => 59,
    12435 => 59,
    12436 => 59,
    12437 => 59,
    12438 => 59,
    12439 => 59,
    12440 => 59,
    12441 => 59,
    12442 => 59,
    12443 => 59,
    12444 => 59,
    12445 => 59,
    12446 => 59,
    12447 => 59,
    12448 => 59,
    12449 => 59,
    12450 => 59,
    12451 => 59,
    12452 => 59,
    12453 => 59,
    12454 => 59,
    12455 => 59,
    12456 => 59,
    12457 => 59,
    12458 => 59,
    12459 => 59,
    12460 => 59,
    12461 => 59,
    12462 => 59,
    12463 => 59,
    12464 => 59,
    12465 => 59,
    12466 => 59,
    12467 => 59,
    12468 => 59,
    12469 => 59,
    12470 => 59,
    12471 => 59,
    12472 => 59,
    12473 => 59,
    12474 => 59,
    12475 => 59,
    12476 => 59,
    12477 => 59,
    12478 => 59,
    12479 => 59,
    12480 => 59,
    12481 => 59,
    12482 => 59,
    12483 => 59,
    12484 => 59,
    12485 => 59,
    12486 => 59,
    12487 => 59,
    12488 => 59,
    12489 => 59,
    12490 => 59,
    12491 => 59,
    12492 => 59,
    12493 => 59,
    12494 => 59,
    12495 => 59,
    12496 => 59,
    12497 => 59,
    12498 => 59,
    12499 => 59,
    12500 => 59,
    12501 => 59,
    12502 => 59,
    12503 => 59,
    12504 => 59,
    12505 => 59,
    12506 => 59,
    12507 => 59,
    12508 => 59,
    12509 => 59,
    12510 => 59,
    12511 => 59,
    12512 => 59,
    12513 => 59,
    12514 => 59,
    12515 => 59,
    12516 => 59,
    12517 => 59,
    12518 => 59,
    12519 => 59,
    12520 => 59,
    12521 => 59,
    12522 => 59,
    12523 => 59,
    12524 => 59,
    12525 => 59,
    12526 => 59,
    12527 => 59,
    12528 => 59,
    12529 => 59,
    12530 => 59,
    12531 => 59,
    12532 => 59,
    12533 => 59,
    12534 => 59,
    12535 => 59,
    12536 => 59,
    12537 => 59,
    12538 => 59,
    12539 => 59,
    12540 => 59,
    12541 => 59,
    12542 => 59,
    12543 => 59,
    12544 => 59,
    12545 => 59,
    12546 => 59,
    12547 => 59,
    12548 => 59,
    12549 => 59,
    12550 => 59,
    12551 => 59,
    12552 => 59,
    12553 => 59,
    12554 => 59,
    12555 => 59,
    12556 => 59,
    12557 => 59,
    12558 => 59,
    12559 => 59,
    12560 => 59,
    12561 => 59,
    12562 => 59,
    12563 => 59,
    12564 => 59,
    12565 => 59,
    12566 => 59,
    12567 => 59,
    12568 => 59,
    12569 => 59,
    12570 => 59,
    12571 => 59,
    12572 => 59,
    12573 => 59,
    12574 => 59,
    12575 => 59,
    12576 => 59,
    12577 => 59,
    12578 => 59,
    12579 => 59,
    12580 => 59,
    12581 => 59,
    12582 => 59,
    12583 => 59,
    12584 => 59,
    12585 => 59,
    12586 => 59,
    12587 => 59,
    12588 => 59,
    12589 => 59,
    12590 => 59,
    12591 => 59,
    12592 => 59,
    12593 => 59,
    12594 => 59,
    12595 => 59,
    12596 => 59,
    12597 => 59,
    12598 => 59,
    12599 => 59,
    12600 => 59,
    12601 => 59,
    12602 => 59,
    12603 => 59,
    12604 => 59,
    12605 => 59,
    12606 => 59,
    12607 => 59,
    12608 => 59,
    12609 => 59,
    12610 => 59,
    12611 => 59,
    12612 => 59,
    12613 => 59,
    12614 => 59,
    12615 => 59,
    12616 => 59,
    12617 => 59,
    12618 => 59,
    12619 => 59,
    12620 => 59,
    12621 => 59,
    12622 => 59,
    12623 => 59,
    12624 => 59,
    12625 => 59,
    12626 => 59,
    12627 => 59,
    12628 => 59,
    12629 => 59,
    12630 => 59,
    12631 => 59,
    12632 => 59,
    12633 => 59,
    12634 => 59,
    12635 => 59,
    12636 => 59,
    12637 => 59,
    12638 => 59,
    12639 => 59,
    12640 => 59,
    12641 => 59,
    12642 => 59,
    12643 => 59,
    12644 => 59,
    12645 => 59,
    12646 => 59,
    12647 => 59,
    12648 => 59,
    12649 => 59,
    12650 => 59,
    12651 => 59,
    12652 => 59,
    12653 => 59,
    12654 => 59,
    12655 => 59,
    12656 => 59,
    12657 => 59,
    12658 => 59,
    12659 => 59,
    12660 => 59,
    12661 => 59,
    12662 => 59,
    12663 => 59,
    12664 => 59,
    12665 => 59,
    12666 => 59,
    12667 => 59,
    12668 => 59,
    12669 => 59,
    12670 => 59,
    12671 => 59,
    12672 => 59,
    12673 => 59,
    12674 => 59,
    12675 => 59,
    12676 => 59,
    12677 => 59,
    12678 => 59,
    12679 => 59,
    12680 => 59,
    12681 => 59,
    12682 => 59,
    12683 => 59,
    12684 => 59,
    12685 => 59,
    12686 => 59,
    12687 => 59,
    12688 => 59,
    12689 => 59,
    12690 => 59,
    12691 => 59,
    12692 => 59,
    12693 => 59,
    12694 => 59,
    12695 => 59,
    12696 => 59,
    12697 => 59,
    12698 => 59,
    12699 => 59,
    12700 => 59,
    12701 => 59,
    12702 => 59,
    12703 => 59,
    12704 => 59,
    12705 => 59,
    12706 => 59,
    12707 => 59,
    12708 => 59,
    12709 => 59,
    12710 => 59,
    12711 => 59,
    12712 => 59,
    12713 => 59,
    12714 => 59,
    12715 => 59,
    12716 => 59,
    12717 => 59,
    12718 => 59,
    12719 => 59,
    12720 => 59,
    12721 => 59,
    12722 => 59,
    12723 => 59,
    12724 => 59,
    12725 => 59,
    12726 => 59,
    12727 => 59,
    12728 => 59,
    12729 => 59,
    12730 => 59,
    12731 => 59,
    12732 => 59,
    12733 => 59,
    12734 => 59,
    12735 => 59,
    12736 => 59,
    12737 => 59,
    12738 => 59,
    12739 => 59,
    12740 => 59,
    12741 => 59,
    12742 => 59,
    12743 => 59,
    12744 => 59,
    12745 => 59,
    12746 => 59,
    12747 => 59,
    12748 => 59,
    12749 => 59,
    12750 => 59,
    12751 => 59,
    12752 => 59,
    12753 => 59,
    12754 => 59,
    12755 => 59,
    12756 => 59,
    12757 => 59,
    12758 => 59,
    12759 => 59,
    12760 => 59,
    12761 => 59,
    12762 => 59,
    12763 => 59,
    12764 => 59,
    12765 => 59,
    12766 => 59,
    12767 => 59,
    12768 => 59,
    12769 => 59,
    12770 => 59,
    12771 => 59,
    12772 => 59,
    12773 => 59,
    12774 => 59,
    12775 => 59,
    12776 => 59,
    12777 => 59,
    12778 => 59,
    12779 => 59,
    12780 => 59,
    12781 => 59,
    12782 => 59,
    12783 => 59,
    12784 => 59,
    12785 => 59,
    12786 => 59,
    12787 => 59,
    12788 => 59,
    12789 => 59,
    12790 => 59,
    12791 => 59,
    12792 => 59,
    12793 => 59,
    12794 => 59,
    12795 => 59,
    12796 => 59,
    12797 => 59,
    12798 => 59,
    12799 => 59,
    12800 => 59,
    12801 => 59,
    12802 => 59,
    12803 => 59,
    12804 => 59,
    12805 => 59,
    12806 => 59,
    12807 => 59,
    12808 => 59,
    12809 => 59,
    12810 => 59,
    12811 => 59,
    12812 => 59,
    12813 => 59,
    12814 => 59,
    12815 => 59,
    12816 => 59,
    12817 => 59,
    12818 => 59,
    12819 => 59,
    12820 => 59,
    12821 => 59,
    12822 => 59,
    12823 => 59,
    12824 => 59,
    12825 => 59,
    12826 => 59,
    12827 => 59,
    12828 => 59,
    12829 => 59,
    12830 => 59,
    12831 => 59,
    12832 => 59,
    12833 => 59,
    12834 => 59,
    12835 => 59,
    12836 => 59,
    12837 => 59,
    12838 => 59,
    12839 => 59,
    12840 => 59,
    12841 => 59,
    12842 => 59,
    12843 => 59,
    12844 => 59,
    12845 => 59,
    12846 => 59,
    12847 => 59,
    12848 => 59,
    12849 => 59,
    12850 => 59,
    12851 => 59,
    12852 => 59,
    12853 => 59,
    12854 => 59,
    12855 => 59,
    12856 => 59,
    12857 => 59,
    12858 => 59,
    12859 => 59,
    12860 => 59,
    12861 => 59,
    12862 => 59,
    12863 => 59,
    12864 => 59,
    12865 => 59,
    12866 => 59,
    12867 => 59,
    12868 => 59,
    12869 => 59,
    12870 => 59,
    12871 => 59,
    12872 => 59,
    12873 => 59,
    12874 => 59,
    12875 => 59,
    12876 => 59,
    12877 => 59,
    12878 => 59,
    12879 => 59,
    12880 => 59,
    12881 => 59,
    12882 => 59,
    12883 => 59,
    12884 => 59,
    12885 => 59,
    12886 => 59,
    12887 => 59,
    12888 => 59,
    12889 => 59,
    12890 => 59,
    12891 => 60,
    12892 => 60,
    12893 => 60,
    12894 => 60,
    12895 => 60,
    12896 => 60,
    12897 => 60,
    12898 => 60,
    12899 => 60,
    12900 => 60,
    12901 => 60,
    12902 => 60,
    12903 => 60,
    12904 => 60,
    12905 => 60,
    12906 => 60,
    12907 => 60,
    12908 => 60,
    12909 => 60,
    12910 => 60,
    12911 => 60,
    12912 => 60,
    12913 => 60,
    12914 => 60,
    12915 => 60,
    12916 => 60,
    12917 => 60,
    12918 => 60,
    12919 => 60,
    12920 => 60,
    12921 => 60,
    12922 => 60,
    12923 => 60,
    12924 => 60,
    12925 => 60,
    12926 => 60,
    12927 => 60,
    12928 => 60,
    12929 => 60,
    12930 => 60,
    12931 => 60,
    12932 => 60,
    12933 => 60,
    12934 => 60,
    12935 => 60,
    12936 => 60,
    12937 => 60,
    12938 => 60,
    12939 => 60,
    12940 => 60,
    12941 => 60,
    12942 => 60,
    12943 => 60,
    12944 => 60,
    12945 => 60,
    12946 => 60,
    12947 => 60,
    12948 => 60,
    12949 => 60,
    12950 => 60,
    12951 => 60,
    12952 => 60,
    12953 => 60,
    12954 => 60,
    12955 => 60,
    12956 => 60,
    12957 => 60,
    12958 => 60,
    12959 => 60,
    12960 => 60,
    12961 => 60,
    12962 => 60,
    12963 => 60,
    12964 => 60,
    12965 => 60,
    12966 => 60,
    12967 => 60,
    12968 => 60,
    12969 => 60,
    12970 => 60,
    12971 => 60,
    12972 => 60,
    12973 => 60,
    12974 => 60,
    12975 => 60,
    12976 => 60,
    12977 => 60,
    12978 => 60,
    12979 => 60,
    12980 => 60,
    12981 => 60,
    12982 => 60,
    12983 => 60,
    12984 => 60,
    12985 => 60,
    12986 => 60,
    12987 => 60,
    12988 => 60,
    12989 => 60,
    12990 => 60,
    12991 => 60,
    12992 => 60,
    12993 => 60,
    12994 => 60,
    12995 => 60,
    12996 => 60,
    12997 => 60,
    12998 => 60,
    12999 => 60,
    13000 => 60,
    13001 => 60,
    13002 => 60,
    13003 => 60,
    13004 => 60,
    13005 => 60,
    13006 => 60,
    13007 => 60,
    13008 => 60,
    13009 => 60,
    13010 => 60,
    13011 => 60,
    13012 => 60,
    13013 => 60,
    13014 => 60,
    13015 => 60,
    13016 => 60,
    13017 => 60,
    13018 => 60,
    13019 => 60,
    13020 => 60,
    13021 => 60,
    13022 => 60,
    13023 => 60,
    13024 => 60,
    13025 => 60,
    13026 => 60,
    13027 => 60,
    13028 => 60,
    13029 => 60,
    13030 => 60,
    13031 => 60,
    13032 => 60,
    13033 => 60,
    13034 => 60,
    13035 => 60,
    13036 => 60,
    13037 => 60,
    13038 => 60,
    13039 => 60,
    13040 => 60,
    13041 => 60,
    13042 => 60,
    13043 => 60,
    13044 => 60,
    13045 => 60,
    13046 => 60,
    13047 => 60,
    13048 => 60,
    13049 => 60,
    13050 => 60,
    13051 => 60,
    13052 => 60,
    13053 => 60,
    13054 => 60,
    13055 => 60,
    13056 => 60,
    13057 => 60,
    13058 => 60,
    13059 => 60,
    13060 => 60,
    13061 => 60,
    13062 => 60,
    13063 => 60,
    13064 => 60,
    13065 => 60,
    13066 => 60,
    13067 => 60,
    13068 => 60,
    13069 => 60,
    13070 => 60,
    13071 => 60,
    13072 => 60,
    13073 => 60,
    13074 => 60,
    13075 => 60,
    13076 => 60,
    13077 => 60,
    13078 => 60,
    13079 => 60,
    13080 => 60,
    13081 => 60,
    13082 => 60,
    13083 => 60,
    13084 => 60,
    13085 => 60,
    13086 => 60,
    13087 => 60,
    13088 => 60,
    13089 => 60,
    13090 => 60,
    13091 => 60,
    13092 => 60,
    13093 => 60,
    13094 => 60,
    13095 => 60,
    13096 => 60,
    13097 => 60,
    13098 => 60,
    13099 => 60,
    13100 => 60,
    13101 => 60,
    13102 => 60,
    13103 => 60,
    13104 => 60,
    13105 => 60,
    13106 => 60,
    13107 => 60,
    13108 => 60,
    13109 => 60,
    13110 => 60,
    13111 => 60,
    13112 => 60,
    13113 => 60,
    13114 => 60,
    13115 => 60,
    13116 => 60,
    13117 => 60,
    13118 => 60,
    13119 => 60,
    13120 => 60,
    13121 => 60,
    13122 => 60,
    13123 => 60,
    13124 => 60,
    13125 => 60,
    13126 => 60,
    13127 => 60,
    13128 => 60,
    13129 => 60,
    13130 => 60,
    13131 => 60,
    13132 => 60,
    13133 => 60,
    13134 => 60,
    13135 => 60,
    13136 => 60,
    13137 => 60,
    13138 => 60,
    13139 => 60,
    13140 => 60,
    13141 => 60,
    13142 => 60,
    13143 => 60,
    13144 => 60,
    13145 => 60,
    13146 => 60,
    13147 => 60,
    13148 => 60,
    13149 => 60,
    13150 => 60,
    13151 => 60,
    13152 => 60,
    13153 => 60,
    13154 => 60,
    13155 => 60,
    13156 => 60,
    13157 => 60,
    13158 => 60,
    13159 => 60,
    13160 => 60,
    13161 => 60,
    13162 => 60,
    13163 => 60,
    13164 => 60,
    13165 => 60,
    13166 => 60,
    13167 => 60,
    13168 => 60,
    13169 => 60,
    13170 => 60,
    13171 => 60,
    13172 => 60,
    13173 => 60,
    13174 => 60,
    13175 => 60,
    13176 => 60,
    13177 => 60,
    13178 => 60,
    13179 => 60,
    13180 => 60,
    13181 => 60,
    13182 => 60,
    13183 => 60,
    13184 => 60,
    13185 => 60,
    13186 => 60,
    13187 => 60,
    13188 => 60,
    13189 => 60,
    13190 => 60,
    13191 => 60,
    13192 => 60,
    13193 => 60,
    13194 => 60,
    13195 => 60,
    13196 => 60,
    13197 => 60,
    13198 => 60,
    13199 => 60,
    13200 => 60,
    13201 => 60,
    13202 => 60,
    13203 => 60,
    13204 => 60,
    13205 => 60,
    13206 => 60,
    13207 => 60,
    13208 => 60,
    13209 => 60,
    13210 => 60,
    13211 => 60,
    13212 => 60,
    13213 => 60,
    13214 => 60,
    13215 => 60,
    13216 => 60,
    13217 => 60,
    13218 => 60,
    13219 => 60,
    13220 => 60,
    13221 => 60,
    13222 => 60,
    13223 => 60,
    13224 => 60,
    13225 => 60,
    13226 => 60,
    13227 => 60,
    13228 => 60,
    13229 => 60,
    13230 => 60,
    13231 => 60,
    13232 => 60,
    13233 => 60,
    13234 => 60,
    13235 => 60,
    13236 => 60,
    13237 => 60,
    13238 => 60,
    13239 => 60,
    13240 => 60,
    13241 => 60,
    13242 => 60,
    13243 => 60,
    13244 => 60,
    13245 => 60,
    13246 => 60,
    13247 => 60,
    13248 => 60,
    13249 => 60,
    13250 => 60,
    13251 => 60,
    13252 => 60,
    13253 => 60,
    13254 => 60,
    13255 => 60,
    13256 => 60,
    13257 => 60,
    13258 => 60,
    13259 => 60,
    13260 => 60,
    13261 => 60,
    13262 => 60,
    13263 => 60,
    13264 => 60,
    13265 => 60,
    13266 => 60,
    13267 => 60,
    13268 => 60,
    13269 => 60,
    13270 => 60,
    13271 => 60,
    13272 => 60,
    13273 => 60,
    13274 => 60,
    13275 => 60,
    13276 => 60,
    13277 => 60,
    13278 => 60,
    13279 => 60,
    13280 => 60,
    13281 => 60,
    13282 => 60,
    13283 => 60,
    13284 => 60,
    13285 => 60,
    13286 => 60,
    13287 => 60,
    13288 => 60,
    13289 => 60,
    13290 => 60,
    13291 => 60,
    13292 => 60,
    13293 => 60,
    13294 => 60,
    13295 => 60,
    13296 => 60,
    13297 => 60,
    13298 => 60,
    13299 => 60,
    13300 => 60,
    13301 => 60,
    13302 => 60,
    13303 => 60,
    13304 => 60,
    13305 => 60,
    13306 => 60,
    13307 => 60,
    13308 => 60,
    13309 => 60,
    13310 => 60,
    13311 => 60,
    13312 => 60,
    13313 => 60,
    13314 => 60,
    13315 => 60,
    13316 => 60,
    13317 => 60,
    13318 => 60,
    13319 => 60,
    13320 => 60,
    13321 => 60,
    13322 => 60,
    13323 => 60,
    13324 => 60,
    13325 => 60,
    13326 => 60,
    13327 => 60,
    13328 => 60,
    13329 => 60,
    13330 => 60,
    13331 => 60,
    13332 => 60,
    13333 => 60,
    13334 => 60,
    13335 => 60,
    13336 => 60,
    13337 => 60,
    13338 => 60,
    13339 => 60,
    13340 => 60,
    13341 => 60,
    13342 => 60,
    13343 => 60,
    13344 => 60,
    13345 => 60,
    13346 => 60,
    13347 => 60,
    13348 => 60,
    13349 => 60,
    13350 => 60,
    13351 => 60,
    13352 => 60,
    13353 => 60,
    13354 => 60,
    13355 => 60,
    13356 => 60,
    13357 => 60,
    13358 => 60,
    13359 => 60,
    13360 => 60,
    13361 => 60,
    13362 => 60,
    13363 => 60,
    13364 => 60,
    13365 => 60,
    13366 => 60,
    13367 => 60,
    13368 => 60,
    13369 => 60,
    13370 => 60,
    13371 => 60,
    13372 => 60,
    13373 => 60,
    13374 => 60,
    13375 => 60,
    13376 => 60,
    13377 => 60,
    13378 => 60,
    13379 => 60,
    13380 => 60,
    13381 => 60,
    13382 => 60,
    13383 => 60,
    13384 => 60,
    13385 => 60,
    13386 => 60,
    13387 => 60,
    13388 => 60,
    13389 => 60,
    13390 => 60,
    13391 => 60,
    13392 => 60,
    13393 => 60,
    13394 => 60,
    13395 => 60,
    13396 => 60,
    13397 => 60,
    13398 => 60,
    13399 => 60,
    13400 => 60,
    13401 => 60,
    13402 => 60,
    13403 => 60,
    13404 => 60,
    13405 => 60,
    13406 => 60,
    13407 => 60,
    13408 => 60,
    13409 => 60,
    13410 => 60,
    13411 => 60,
    13412 => 60,
    13413 => 60,
    13414 => 60,
    13415 => 60,
    13416 => 60,
    13417 => 60,
    13418 => 60,
    13419 => 60,
    13420 => 60,
    13421 => 60,
    13422 => 60,
    13423 => 60,
    13424 => 60,
    13425 => 60,
    13426 => 60,
    13427 => 60,
    13428 => 60,
    13429 => 60,
    13430 => 60,
    13431 => 60,
    13432 => 60,
    13433 => 60,
    13434 => 60,
    13435 => 60,
    13436 => 61,
    13437 => 61,
    13438 => 61,
    13439 => 61,
    13440 => 61,
    13441 => 61,
    13442 => 61,
    13443 => 61,
    13444 => 61,
    13445 => 61,
    13446 => 61,
    13447 => 61,
    13448 => 61,
    13449 => 61,
    13450 => 61,
    13451 => 61,
    13452 => 61,
    13453 => 61,
    13454 => 61,
    13455 => 61,
    13456 => 61,
    13457 => 61,
    13458 => 61,
    13459 => 61,
    13460 => 61,
    13461 => 61,
    13462 => 61,
    13463 => 61,
    13464 => 61,
    13465 => 61,
    13466 => 61,
    13467 => 61,
    13468 => 61,
    13469 => 61,
    13470 => 61,
    13471 => 61,
    13472 => 61,
    13473 => 61,
    13474 => 61,
    13475 => 61,
    13476 => 61,
    13477 => 61,
    13478 => 61,
    13479 => 61,
    13480 => 61,
    13481 => 61,
    13482 => 61,
    13483 => 61,
    13484 => 61,
    13485 => 61,
    13486 => 61,
    13487 => 61,
    13488 => 61,
    13489 => 61,
    13490 => 61,
    13491 => 61,
    13492 => 61,
    13493 => 61,
    13494 => 61,
    13495 => 61,
    13496 => 61,
    13497 => 61,
    13498 => 61,
    13499 => 61,
    13500 => 61,
    13501 => 61,
    13502 => 61,
    13503 => 61,
    13504 => 61,
    13505 => 61,
    13506 => 61,
    13507 => 61,
    13508 => 61,
    13509 => 61,
    13510 => 61,
    13511 => 61,
    13512 => 61,
    13513 => 61,
    13514 => 61,
    13515 => 61,
    13516 => 61,
    13517 => 61,
    13518 => 61,
    13519 => 61,
    13520 => 61,
    13521 => 61,
    13522 => 61,
    13523 => 61,
    13524 => 61,
    13525 => 61,
    13526 => 61,
    13527 => 61,
    13528 => 61,
    13529 => 61,
    13530 => 61,
    13531 => 61,
    13532 => 61,
    13533 => 61,
    13534 => 61,
    13535 => 61,
    13536 => 61,
    13537 => 61,
    13538 => 61,
    13539 => 61,
    13540 => 61,
    13541 => 61,
    13542 => 61,
    13543 => 61,
    13544 => 61,
    13545 => 61,
    13546 => 61,
    13547 => 61,
    13548 => 61,
    13549 => 61,
    13550 => 61,
    13551 => 61,
    13552 => 61,
    13553 => 61,
    13554 => 61,
    13555 => 61,
    13556 => 61,
    13557 => 61,
    13558 => 61,
    13559 => 61,
    13560 => 61,
    13561 => 61,
    13562 => 61,
    13563 => 61,
    13564 => 61,
    13565 => 61,
    13566 => 61,
    13567 => 61,
    13568 => 61,
    13569 => 61,
    13570 => 61,
    13571 => 61,
    13572 => 61,
    13573 => 61,
    13574 => 61,
    13575 => 61,
    13576 => 61,
    13577 => 61,
    13578 => 61,
    13579 => 61,
    13580 => 61,
    13581 => 61,
    13582 => 61,
    13583 => 61,
    13584 => 61,
    13585 => 61,
    13586 => 61,
    13587 => 61,
    13588 => 61,
    13589 => 61,
    13590 => 61,
    13591 => 61,
    13592 => 61,
    13593 => 61,
    13594 => 61,
    13595 => 61,
    13596 => 61,
    13597 => 61,
    13598 => 61,
    13599 => 61,
    13600 => 61,
    13601 => 61,
    13602 => 61,
    13603 => 61,
    13604 => 61,
    13605 => 61,
    13606 => 61,
    13607 => 61,
    13608 => 61,
    13609 => 61,
    13610 => 61,
    13611 => 61,
    13612 => 61,
    13613 => 61,
    13614 => 61,
    13615 => 61,
    13616 => 61,
    13617 => 61,
    13618 => 61,
    13619 => 61,
    13620 => 61,
    13621 => 61,
    13622 => 61,
    13623 => 61,
    13624 => 61,
    13625 => 61,
    13626 => 61,
    13627 => 61,
    13628 => 61,
    13629 => 61,
    13630 => 61,
    13631 => 61,
    13632 => 61,
    13633 => 61,
    13634 => 61,
    13635 => 61,
    13636 => 61,
    13637 => 61,
    13638 => 61,
    13639 => 61,
    13640 => 61,
    13641 => 61,
    13642 => 61,
    13643 => 61,
    13644 => 61,
    13645 => 61,
    13646 => 61,
    13647 => 61,
    13648 => 61,
    13649 => 61,
    13650 => 61,
    13651 => 61,
    13652 => 61,
    13653 => 61,
    13654 => 61,
    13655 => 61,
    13656 => 61,
    13657 => 61,
    13658 => 61,
    13659 => 61,
    13660 => 61,
    13661 => 61,
    13662 => 61,
    13663 => 61,
    13664 => 61,
    13665 => 61,
    13666 => 61,
    13667 => 61,
    13668 => 61,
    13669 => 61,
    13670 => 61,
    13671 => 61,
    13672 => 61,
    13673 => 61,
    13674 => 61,
    13675 => 61,
    13676 => 61,
    13677 => 61,
    13678 => 61,
    13679 => 61,
    13680 => 61,
    13681 => 61,
    13682 => 61,
    13683 => 61,
    13684 => 61,
    13685 => 61,
    13686 => 61,
    13687 => 61,
    13688 => 61,
    13689 => 61,
    13690 => 61,
    13691 => 61,
    13692 => 61,
    13693 => 61,
    13694 => 61,
    13695 => 61,
    13696 => 61,
    13697 => 61,
    13698 => 61,
    13699 => 61,
    13700 => 61,
    13701 => 61,
    13702 => 61,
    13703 => 61,
    13704 => 61,
    13705 => 61,
    13706 => 61,
    13707 => 61,
    13708 => 61,
    13709 => 61,
    13710 => 61,
    13711 => 61,
    13712 => 61,
    13713 => 61,
    13714 => 61,
    13715 => 61,
    13716 => 61,
    13717 => 61,
    13718 => 61,
    13719 => 61,
    13720 => 61,
    13721 => 61,
    13722 => 61,
    13723 => 61,
    13724 => 61,
    13725 => 61,
    13726 => 61,
    13727 => 61,
    13728 => 61,
    13729 => 61,
    13730 => 61,
    13731 => 61,
    13732 => 61,
    13733 => 61,
    13734 => 61,
    13735 => 61,
    13736 => 61,
    13737 => 61,
    13738 => 61,
    13739 => 61,
    13740 => 61,
    13741 => 61,
    13742 => 61,
    13743 => 61,
    13744 => 61,
    13745 => 61,
    13746 => 61,
    13747 => 61,
    13748 => 61,
    13749 => 61,
    13750 => 61,
    13751 => 61,
    13752 => 61,
    13753 => 61,
    13754 => 61,
    13755 => 61,
    13756 => 61,
    13757 => 61,
    13758 => 61,
    13759 => 61,
    13760 => 61,
    13761 => 61,
    13762 => 61,
    13763 => 61,
    13764 => 61,
    13765 => 61,
    13766 => 61,
    13767 => 61,
    13768 => 61,
    13769 => 61,
    13770 => 61,
    13771 => 61,
    13772 => 61,
    13773 => 61,
    13774 => 61,
    13775 => 61,
    13776 => 61,
    13777 => 61,
    13778 => 61,
    13779 => 61,
    13780 => 61,
    13781 => 61,
    13782 => 61,
    13783 => 61,
    13784 => 61,
    13785 => 61,
    13786 => 61,
    13787 => 61,
    13788 => 61,
    13789 => 61,
    13790 => 61,
    13791 => 61,
    13792 => 61,
    13793 => 61,
    13794 => 61,
    13795 => 61,
    13796 => 61,
    13797 => 61,
    13798 => 61,
    13799 => 61,
    13800 => 61,
    13801 => 61,
    13802 => 61,
    13803 => 61,
    13804 => 61,
    13805 => 61,
    13806 => 61,
    13807 => 61,
    13808 => 61,
    13809 => 61,
    13810 => 61,
    13811 => 61,
    13812 => 61,
    13813 => 61,
    13814 => 61,
    13815 => 61,
    13816 => 61,
    13817 => 61,
    13818 => 61,
    13819 => 61,
    13820 => 61,
    13821 => 61,
    13822 => 61,
    13823 => 61,
    13824 => 61,
    13825 => 61,
    13826 => 61,
    13827 => 61,
    13828 => 61,
    13829 => 61,
    13830 => 61,
    13831 => 61,
    13832 => 61,
    13833 => 61,
    13834 => 61,
    13835 => 61,
    13836 => 61,
    13837 => 61,
    13838 => 61,
    13839 => 61,
    13840 => 61,
    13841 => 61,
    13842 => 61,
    13843 => 61,
    13844 => 61,
    13845 => 61,
    13846 => 61,
    13847 => 61,
    13848 => 61,
    13849 => 61,
    13850 => 61,
    13851 => 61,
    13852 => 61,
    13853 => 61,
    13854 => 61,
    13855 => 61,
    13856 => 61,
    13857 => 61,
    13858 => 61,
    13859 => 61,
    13860 => 61,
    13861 => 61,
    13862 => 61,
    13863 => 61,
    13864 => 61,
    13865 => 61,
    13866 => 61,
    13867 => 61,
    13868 => 61,
    13869 => 61,
    13870 => 61,
    13871 => 61,
    13872 => 61,
    13873 => 61,
    13874 => 61,
    13875 => 61,
    13876 => 61,
    13877 => 61,
    13878 => 61,
    13879 => 61,
    13880 => 61,
    13881 => 61,
    13882 => 61,
    13883 => 61,
    13884 => 61,
    13885 => 61,
    13886 => 61,
    13887 => 61,
    13888 => 61,
    13889 => 61,
    13890 => 61,
    13891 => 61,
    13892 => 61,
    13893 => 61,
    13894 => 61,
    13895 => 61,
    13896 => 61,
    13897 => 61,
    13898 => 61,
    13899 => 61,
    13900 => 61,
    13901 => 61,
    13902 => 61,
    13903 => 61,
    13904 => 61,
    13905 => 61,
    13906 => 61,
    13907 => 61,
    13908 => 61,
    13909 => 61,
    13910 => 61,
    13911 => 61,
    13912 => 61,
    13913 => 61,
    13914 => 61,
    13915 => 61,
    13916 => 61,
    13917 => 61,
    13918 => 61,
    13919 => 61,
    13920 => 61,
    13921 => 61,
    13922 => 61,
    13923 => 61,
    13924 => 61,
    13925 => 61,
    13926 => 61,
    13927 => 61,
    13928 => 61,
    13929 => 61,
    13930 => 61,
    13931 => 61,
    13932 => 61,
    13933 => 61,
    13934 => 61,
    13935 => 61,
    13936 => 61,
    13937 => 61,
    13938 => 61,
    13939 => 61,
    13940 => 61,
    13941 => 61,
    13942 => 61,
    13943 => 61,
    13944 => 61,
    13945 => 61,
    13946 => 61,
    13947 => 61,
    13948 => 61,
    13949 => 61,
    13950 => 61,
    13951 => 61,
    13952 => 61,
    13953 => 61,
    13954 => 61,
    13955 => 61,
    13956 => 61,
    13957 => 61,
    13958 => 61,
    13959 => 61,
    13960 => 61,
    13961 => 61,
    13962 => 61,
    13963 => 61,
    13964 => 61,
    13965 => 61,
    13966 => 61,
    13967 => 61,
    13968 => 61,
    13969 => 61,
    13970 => 61,
    13971 => 61,
    13972 => 61,
    13973 => 61,
    13974 => 61,
    13975 => 61,
    13976 => 61,
    13977 => 61,
    13978 => 61,
    13979 => 61,
    13980 => 61,
    13981 => 61,
    13982 => 61,
    13983 => 61,
    13984 => 61,
    13985 => 61,
    13986 => 61,
    13987 => 61,
    13988 => 61,
    13989 => 61,
    13990 => 61,
    13991 => 61,
    13992 => 61,
    13993 => 61,
    13994 => 61,
    13995 => 61,
    13996 => 61,
    13997 => 61,
    13998 => 61,
    13999 => 61,
    14000 => 61,
    14001 => 61,
    14002 => 61,
    14003 => 61,
    14004 => 61,
    14005 => 61,
    14006 => 61,
    14007 => 61,
    14008 => 61,
    14009 => 61,
    14010 => 61,
    14011 => 61,
    14012 => 61,
    14013 => 61,
    14014 => 61,
    14015 => 61,
    14016 => 61,
    14017 => 61,
    14018 => 61,
    14019 => 61,
    14020 => 61,
    14021 => 61,
    14022 => 61,
    14023 => 61,
    14024 => 61,
    14025 => 61,
    14026 => 61,
    14027 => 61,
    14028 => 61,
    14029 => 61,
    14030 => 61,
    14031 => 61,
    14032 => 61,
    14033 => 61,
    14034 => 61,
    14035 => 61,
    14036 => 61,
    14037 => 61,
    14038 => 61,
    14039 => 61,
    14040 => 61,
    14041 => 61,
    14042 => 61,
    14043 => 61,
    14044 => 61,
    14045 => 61,
    14046 => 61,
    14047 => 61,
    14048 => 61,
    14049 => 61,
    14050 => 61,
    14051 => 61,
    14052 => 61,
    14053 => 61,
    14054 => 61,
    14055 => 61,
    14056 => 61,
    14057 => 61,
    14058 => 61,
    14059 => 61,
    14060 => 61,
    14061 => 61,
    14062 => 61,
    14063 => 61,
    14064 => 61,
    14065 => 61,
    14066 => 61,
    14067 => 61,
    14068 => 61,
    14069 => 61,
    14070 => 61,
    14071 => 61,
    14072 => 61,
    14073 => 61,
    14074 => 61,
    14075 => 61,
    14076 => 61,
    14077 => 61,
    14078 => 61,
    14079 => 61,
    14080 => 61,
    14081 => 61,
    14082 => 61,
    14083 => 61,
    14084 => 61,
    14085 => 61,
    14086 => 61,
    14087 => 61,
    14088 => 61,
    14089 => 61,
    14090 => 61,
    14091 => 61,
    14092 => 61,
    14093 => 61,
    14094 => 61,
    14095 => 61,
    14096 => 61,
    14097 => 61,
    14098 => 61,
    14099 => 61,
    14100 => 61,
    14101 => 61,
    14102 => 61,
    14103 => 61,
    14104 => 62,
    14105 => 62,
    14106 => 62,
    14107 => 62,
    14108 => 62,
    14109 => 62,
    14110 => 62,
    14111 => 62,
    14112 => 62,
    14113 => 62,
    14114 => 62,
    14115 => 62,
    14116 => 62,
    14117 => 62,
    14118 => 62,
    14119 => 62,
    14120 => 62,
    14121 => 62,
    14122 => 62,
    14123 => 62,
    14124 => 62,
    14125 => 62,
    14126 => 62,
    14127 => 62,
    14128 => 62,
    14129 => 62,
    14130 => 62,
    14131 => 62,
    14132 => 62,
    14133 => 62,
    14134 => 62,
    14135 => 62,
    14136 => 62,
    14137 => 62,
    14138 => 62,
    14139 => 62,
    14140 => 62,
    14141 => 62,
    14142 => 62,
    14143 => 62,
    14144 => 62,
    14145 => 62,
    14146 => 62,
    14147 => 62,
    14148 => 62,
    14149 => 62,
    14150 => 62,
    14151 => 62,
    14152 => 62,
    14153 => 62,
    14154 => 62,
    14155 => 62,
    14156 => 62,
    14157 => 62,
    14158 => 62,
    14159 => 62,
    14160 => 62,
    14161 => 62,
    14162 => 62,
    14163 => 62,
    14164 => 62,
    14165 => 62,
    14166 => 62,
    14167 => 62,
    14168 => 62,
    14169 => 62,
    14170 => 62,
    14171 => 62,
    14172 => 62,
    14173 => 62,
    14174 => 62,
    14175 => 62,
    14176 => 62,
    14177 => 62,
    14178 => 62,
    14179 => 62,
    14180 => 62,
    14181 => 62,
    14182 => 62,
    14183 => 62,
    14184 => 62,
    14185 => 62,
    14186 => 62,
    14187 => 62,
    14188 => 62,
    14189 => 62,
    14190 => 62,
    14191 => 62,
    14192 => 62,
    14193 => 62,
    14194 => 62,
    14195 => 62,
    14196 => 62,
    14197 => 62,
    14198 => 62,
    14199 => 62,
    14200 => 62,
    14201 => 62,
    14202 => 62,
    14203 => 62,
    14204 => 62,
    14205 => 62,
    14206 => 62,
    14207 => 62,
    14208 => 62,
    14209 => 62,
    14210 => 62,
    14211 => 62,
    14212 => 62,
    14213 => 62,
    14214 => 62,
    14215 => 62,
    14216 => 62,
    14217 => 62,
    14218 => 62,
    14219 => 62,
    14220 => 62,
    14221 => 62,
    14222 => 62,
    14223 => 62,
    14224 => 62,
    14225 => 62,
    14226 => 62,
    14227 => 62,
    14228 => 62,
    14229 => 62,
    14230 => 62,
    14231 => 62,
    14232 => 62,
    14233 => 62,
    14234 => 62,
    14235 => 62,
    14236 => 62,
    14237 => 62,
    14238 => 62,
    14239 => 62,
    14240 => 62,
    14241 => 62,
    14242 => 62,
    14243 => 62,
    14244 => 62,
    14245 => 62,
    14246 => 62,
    14247 => 62,
    14248 => 62,
    14249 => 62,
    14250 => 62,
    14251 => 62,
    14252 => 62,
    14253 => 62,
    14254 => 62,
    14255 => 62,
    14256 => 62,
    14257 => 62,
    14258 => 62,
    14259 => 62,
    14260 => 62,
    14261 => 62,
    14262 => 62,
    14263 => 62,
    14264 => 62,
    14265 => 62,
    14266 => 62,
    14267 => 62,
    14268 => 62,
    14269 => 62,
    14270 => 62,
    14271 => 62,
    14272 => 62,
    14273 => 62,
    14274 => 62,
    14275 => 62,
    14276 => 62,
    14277 => 62,
    14278 => 62,
    14279 => 62,
    14280 => 62,
    14281 => 62,
    14282 => 62,
    14283 => 62,
    14284 => 62,
    14285 => 62,
    14286 => 62,
    14287 => 62,
    14288 => 62,
    14289 => 62,
    14290 => 62,
    14291 => 62,
    14292 => 62,
    14293 => 62,
    14294 => 62,
    14295 => 62,
    14296 => 62,
    14297 => 62,
    14298 => 62,
    14299 => 62,
    14300 => 62,
    14301 => 62,
    14302 => 62,
    14303 => 62,
    14304 => 62,
    14305 => 62,
    14306 => 62,
    14307 => 62,
    14308 => 62,
    14309 => 62,
    14310 => 62,
    14311 => 62,
    14312 => 62,
    14313 => 62,
    14314 => 62,
    14315 => 62,
    14316 => 62,
    14317 => 62,
    14318 => 62,
    14319 => 62,
    14320 => 62,
    14321 => 62,
    14322 => 62,
    14323 => 62,
    14324 => 62,
    14325 => 62,
    14326 => 62,
    14327 => 62,
    14328 => 62,
    14329 => 62,
    14330 => 62,
    14331 => 62,
    14332 => 62,
    14333 => 62,
    14334 => 62,
    14335 => 62,
    14336 => 62,
    14337 => 62,
    14338 => 62,
    14339 => 62,
    14340 => 62,
    14341 => 62,
    14342 => 62,
    14343 => 62,
    14344 => 62,
    14345 => 62,
    14346 => 62,
    14347 => 62,
    14348 => 62,
    14349 => 62,
    14350 => 62,
    14351 => 62,
    14352 => 62,
    14353 => 62,
    14354 => 62,
    14355 => 62,
    14356 => 62,
    14357 => 62,
    14358 => 62,
    14359 => 62,
    14360 => 62,
    14361 => 62,
    14362 => 62,
    14363 => 62,
    14364 => 62,
    14365 => 62,
    14366 => 62,
    14367 => 62,
    14368 => 62,
    14369 => 62,
    14370 => 62,
    14371 => 62,
    14372 => 62,
    14373 => 62,
    14374 => 62,
    14375 => 62,
    14376 => 62,
    14377 => 62,
    14378 => 62,
    14379 => 62,
    14380 => 62,
    14381 => 62,
    14382 => 62,
    14383 => 62,
    14384 => 62,
    14385 => 62,
    14386 => 62,
    14387 => 62,
    14388 => 62,
    14389 => 62,
    14390 => 62,
    14391 => 62,
    14392 => 62,
    14393 => 62,
    14394 => 62,
    14395 => 62,
    14396 => 62,
    14397 => 62,
    14398 => 62,
    14399 => 62,
    14400 => 62,
    14401 => 62,
    14402 => 62,
    14403 => 62,
    14404 => 62,
    14405 => 62,
    14406 => 62,
    14407 => 62,
    14408 => 62,
    14409 => 62,
    14410 => 62,
    14411 => 62,
    14412 => 62,
    14413 => 62,
    14414 => 62,
    14415 => 62,
    14416 => 62,
    14417 => 62,
    14418 => 62,
    14419 => 62,
    14420 => 62,
    14421 => 62,
    14422 => 62,
    14423 => 62,
    14424 => 62,
    14425 => 62,
    14426 => 62,
    14427 => 62,
    14428 => 62,
    14429 => 62,
    14430 => 62,
    14431 => 62,
    14432 => 62,
    14433 => 62,
    14434 => 62,
    14435 => 62,
    14436 => 62,
    14437 => 62,
    14438 => 62,
    14439 => 62,
    14440 => 62,
    14441 => 62,
    14442 => 62,
    14443 => 62,
    14444 => 62,
    14445 => 62,
    14446 => 62,
    14447 => 62,
    14448 => 62,
    14449 => 62,
    14450 => 62,
    14451 => 62,
    14452 => 62,
    14453 => 62,
    14454 => 62,
    14455 => 62,
    14456 => 62,
    14457 => 62,
    14458 => 62,
    14459 => 62,
    14460 => 62,
    14461 => 62,
    14462 => 62,
    14463 => 62,
    14464 => 62,
    14465 => 62,
    14466 => 62,
    14467 => 62,
    14468 => 62,
    14469 => 62,
    14470 => 62,
    14471 => 62,
    14472 => 62,
    14473 => 62,
    14474 => 62,
    14475 => 62,
    14476 => 62,
    14477 => 62,
    14478 => 62,
    14479 => 62,
    14480 => 62,
    14481 => 62,
    14482 => 62,
    14483 => 62,
    14484 => 62,
    14485 => 62,
    14486 => 62,
    14487 => 62,
    14488 => 62,
    14489 => 62,
    14490 => 62,
    14491 => 62,
    14492 => 62,
    14493 => 62,
    14494 => 62,
    14495 => 62,
    14496 => 62,
    14497 => 62,
    14498 => 62,
    14499 => 62,
    14500 => 62,
    14501 => 62,
    14502 => 62,
    14503 => 62,
    14504 => 62,
    14505 => 62,
    14506 => 62,
    14507 => 62,
    14508 => 62,
    14509 => 62,
    14510 => 62,
    14511 => 62,
    14512 => 62,
    14513 => 62,
    14514 => 62,
    14515 => 62,
    14516 => 62,
    14517 => 62,
    14518 => 62,
    14519 => 62,
    14520 => 62,
    14521 => 62,
    14522 => 62,
    14523 => 62,
    14524 => 62,
    14525 => 62,
    14526 => 62,
    14527 => 62,
    14528 => 62,
    14529 => 62,
    14530 => 62,
    14531 => 62,
    14532 => 62,
    14533 => 62,
    14534 => 62,
    14535 => 62,
    14536 => 62,
    14537 => 62,
    14538 => 62,
    14539 => 62,
    14540 => 62,
    14541 => 62,
    14542 => 62,
    14543 => 62,
    14544 => 62,
    14545 => 62,
    14546 => 62,
    14547 => 62,
    14548 => 62,
    14549 => 62,
    14550 => 62,
    14551 => 62,
    14552 => 62,
    14553 => 62,
    14554 => 62,
    14555 => 62,
    14556 => 62,
    14557 => 62,
    14558 => 62,
    14559 => 62,
    14560 => 62,
    14561 => 62,
    14562 => 62,
    14563 => 62,
    14564 => 62,
    14565 => 62,
    14566 => 62,
    14567 => 62,
    14568 => 62,
    14569 => 62,
    14570 => 62,
    14571 => 62,
    14572 => 62,
    14573 => 62,
    14574 => 62,
    14575 => 62,
    14576 => 62,
    14577 => 62,
    14578 => 62,
    14579 => 62,
    14580 => 62,
    14581 => 62,
    14582 => 62,
    14583 => 62,
    14584 => 62,
    14585 => 62,
    14586 => 62,
    14587 => 62,
    14588 => 62,
    14589 => 62,
    14590 => 62,
    14591 => 62,
    14592 => 62,
    14593 => 62,
    14594 => 62,
    14595 => 62,
    14596 => 62,
    14597 => 62,
    14598 => 62,
    14599 => 62,
    14600 => 62,
    14601 => 62,
    14602 => 62,
    14603 => 62,
    14604 => 62,
    14605 => 62,
    14606 => 62,
    14607 => 62,
    14608 => 62,
    14609 => 62,
    14610 => 62,
    14611 => 62,
    14612 => 62,
    14613 => 62,
    14614 => 62,
    14615 => 62,
    14616 => 62,
    14617 => 62,
    14618 => 62,
    14619 => 62,
    14620 => 62,
    14621 => 62,
    14622 => 62,
    14623 => 62,
    14624 => 62,
    14625 => 62,
    14626 => 62,
    14627 => 62,
    14628 => 62,
    14629 => 62,
    14630 => 62,
    14631 => 62,
    14632 => 62,
    14633 => 62,
    14634 => 62,
    14635 => 62,
    14636 => 62,
    14637 => 62,
    14638 => 62,
    14639 => 62,
    14640 => 62,
    14641 => 62,
    14642 => 62,
    14643 => 62,
    14644 => 62,
    14645 => 62,
    14646 => 62,
    14647 => 62,
    14648 => 62,
    14649 => 62,
    14650 => 62,
    14651 => 62,
    14652 => 62,
    14653 => 62,
    14654 => 62,
    14655 => 62,
    14656 => 62,
    14657 => 62,
    14658 => 62,
    14659 => 62,
    14660 => 62,
    14661 => 62,
    14662 => 62,
    14663 => 62,
    14664 => 62,
    14665 => 62,
    14666 => 62,
    14667 => 62,
    14668 => 62,
    14669 => 62,
    14670 => 62,
    14671 => 62,
    14672 => 62,
    14673 => 62,
    14674 => 62,
    14675 => 62,
    14676 => 62,
    14677 => 62,
    14678 => 62,
    14679 => 62,
    14680 => 62,
    14681 => 62,
    14682 => 62,
    14683 => 62,
    14684 => 62,
    14685 => 62,
    14686 => 62,
    14687 => 62,
    14688 => 62,
    14689 => 62,
    14690 => 62,
    14691 => 62,
    14692 => 62,
    14693 => 62,
    14694 => 62,
    14695 => 62,
    14696 => 62,
    14697 => 62,
    14698 => 62,
    14699 => 62,
    14700 => 62,
    14701 => 62,
    14702 => 62,
    14703 => 62,
    14704 => 62,
    14705 => 62,
    14706 => 62,
    14707 => 62,
    14708 => 62,
    14709 => 62,
    14710 => 62,
    14711 => 62,
    14712 => 62,
    14713 => 62,
    14714 => 62,
    14715 => 62,
    14716 => 62,
    14717 => 62,
    14718 => 62,
    14719 => 62,
    14720 => 62,
    14721 => 62,
    14722 => 62,
    14723 => 62,
    14724 => 62,
    14725 => 62,
    14726 => 62,
    14727 => 62,
    14728 => 62,
    14729 => 62,
    14730 => 62,
    14731 => 62,
    14732 => 62,
    14733 => 62,
    14734 => 62,
    14735 => 62,
    14736 => 62,
    14737 => 62,
    14738 => 62,
    14739 => 62,
    14740 => 62,
    14741 => 62,
    14742 => 62,
    14743 => 62,
    14744 => 62,
    14745 => 62,
    14746 => 62,
    14747 => 62,
    14748 => 62,
    14749 => 62,
    14750 => 62,
    14751 => 62,
    14752 => 62,
    14753 => 62,
    14754 => 62,
    14755 => 62,
    14756 => 62,
    14757 => 62,
    14758 => 62,
    14759 => 62,
    14760 => 62,
    14761 => 62,
    14762 => 62,
    14763 => 62,
    14764 => 62,
    14765 => 62,
    14766 => 62,
    14767 => 62,
    14768 => 62,
    14769 => 62,
    14770 => 62,
    14771 => 62,
    14772 => 62,
    14773 => 62,
    14774 => 62,
    14775 => 62,
    14776 => 62,
    14777 => 62,
    14778 => 62,
    14779 => 62,
    14780 => 62,
    14781 => 62,
    14782 => 62,
    14783 => 62,
    14784 => 62,
    14785 => 62,
    14786 => 62,
    14787 => 62,
    14788 => 62,
    14789 => 62,
    14790 => 62,
    14791 => 62,
    14792 => 62,
    14793 => 62,
    14794 => 62,
    14795 => 62,
    14796 => 62,
    14797 => 62,
    14798 => 62,
    14799 => 62,
    14800 => 62,
    14801 => 62,
    14802 => 62,
    14803 => 62,
    14804 => 62,
    14805 => 62,
    14806 => 62,
    14807 => 62,
    14808 => 62,
    14809 => 62,
    14810 => 62,
    14811 => 62,
    14812 => 62,
    14813 => 62,
    14814 => 62,
    14815 => 62,
    14816 => 62,
    14817 => 62,
    14818 => 62,
    14819 => 62,
    14820 => 62,
    14821 => 62,
    14822 => 62,
    14823 => 62,
    14824 => 62,
    14825 => 62,
    14826 => 62,
    14827 => 62,
    14828 => 62,
    14829 => 62,
    14830 => 62,
    14831 => 62,
    14832 => 62,
    14833 => 62,
    14834 => 62,
    14835 => 62,
    14836 => 62,
    14837 => 62,
    14838 => 62,
    14839 => 62,
    14840 => 62,
    14841 => 62,
    14842 => 62,
    14843 => 62,
    14844 => 62,
    14845 => 62,
    14846 => 62,
    14847 => 62,
    14848 => 62,
    14849 => 62,
    14850 => 62,
    14851 => 62,
    14852 => 62,
    14853 => 62,
    14854 => 62,
    14855 => 62,
    14856 => 62,
    14857 => 62,
    14858 => 62,
    14859 => 62,
    14860 => 62,
    14861 => 62,
    14862 => 62,
    14863 => 62,
    14864 => 62,
    14865 => 62,
    14866 => 62,
    14867 => 62,
    14868 => 62,
    14869 => 62,
    14870 => 62,
    14871 => 62,
    14872 => 62,
    14873 => 62,
    14874 => 62,
    14875 => 62,
    14876 => 62,
    14877 => 62,
    14878 => 62,
    14879 => 62,
    14880 => 62,
    14881 => 62,
    14882 => 62,
    14883 => 62,
    14884 => 62,
    14885 => 62,
    14886 => 62,
    14887 => 62,
    14888 => 62,
    14889 => 62,
    14890 => 62,
    14891 => 62,
    14892 => 62,
    14893 => 62,
    14894 => 62,
    14895 => 62,
    14896 => 62,
    14897 => 62,
    14898 => 62,
    14899 => 62,
    14900 => 62,
    14901 => 62,
    14902 => 62,
    14903 => 62,
    14904 => 62,
    14905 => 62,
    14906 => 62,
    14907 => 62,
    14908 => 62,
    14909 => 62,
    14910 => 62,
    14911 => 62,
    14912 => 62,
    14913 => 62,
    14914 => 62,
    14915 => 62,
    14916 => 62,
    14917 => 62,
    14918 => 62,
    14919 => 62,
    14920 => 62,
    14921 => 62,
    14922 => 62,
    14923 => 62,
    14924 => 62,
    14925 => 62,
    14926 => 62,
    14927 => 62,
    14928 => 62,
    14929 => 62,
    14930 => 62,
    14931 => 62,
    14932 => 62,
    14933 => 62,
    14934 => 62,
    14935 => 62,
    14936 => 62,
    14937 => 62,
    14938 => 62,
    14939 => 62,
    14940 => 62,
    14941 => 62,
    14942 => 62,
    14943 => 62,
    14944 => 62,
    14945 => 62,
    14946 => 62,
    14947 => 62,
    14948 => 62,
    14949 => 62,
    14950 => 62,
    14951 => 62,
    14952 => 62,
    14953 => 62,
    14954 => 62,
    14955 => 62,
    14956 => 62,
    14957 => 62,
    14958 => 62,
    14959 => 62,
    14960 => 62,
    14961 => 62,
    14962 => 62,
    14963 => 62,
    14964 => 62,
    14965 => 62,
    14966 => 62,
    14967 => 62,
    14968 => 62,
    14969 => 62,
    14970 => 62,
    14971 => 62,
    14972 => 62,
    14973 => 62,
    14974 => 62,
    14975 => 62,
    14976 => 62,
    14977 => 62,
    14978 => 62,
    14979 => 62,
    14980 => 62,
    14981 => 62,
    14982 => 62,
    14983 => 62,
    14984 => 62,
    14985 => 62,
    14986 => 62,
    14987 => 62,
    14988 => 62,
    14989 => 62,
    14990 => 62,
    14991 => 62,
    14992 => 62,
    14993 => 62,
    14994 => 62,
    14995 => 62,
    14996 => 62,
    14997 => 62,
    14998 => 62,
    14999 => 62,
    15000 => 62,
    15001 => 62,
    15002 => 62,
    15003 => 62,
    15004 => 62,
    15005 => 62,
    15006 => 62,
    15007 => 62,
    15008 => 62,
    15009 => 62,
    15010 => 62,
    15011 => 62,
    15012 => 62,
    15013 => 62,
    15014 => 62,
    15015 => 62,
    15016 => 62,
    15017 => 62,
    15018 => 62,
    15019 => 62,
    15020 => 62,
    15021 => 62,
    15022 => 62,
    15023 => 62,
    15024 => 62,
    15025 => 62,
    15026 => 62,
    15027 => 62,
    15028 => 62,
    15029 => 62,
    15030 => 62,
    15031 => 62,
    15032 => 62,
    15033 => 62,
    15034 => 62,
    15035 => 62,
    15036 => 62,
    15037 => 62,
    15038 => 62,
    15039 => 62,
    15040 => 62,
    15041 => 62,
    15042 => 62,
    15043 => 62,
    15044 => 62,
    15045 => 62,
    15046 => 62,
    15047 => 62,
    15048 => 62,
    15049 => 62,
    15050 => 62,
    15051 => 62,
    15052 => 62,
    15053 => 62,
    15054 => 62,
    15055 => 62,
    15056 => 62,
    15057 => 62,
    15058 => 62,
    15059 => 62,
    15060 => 62,
    15061 => 62,
    15062 => 62,
    15063 => 62,
    15064 => 62,
    15065 => 62,
    15066 => 62,
    15067 => 62,
    15068 => 62,
    15069 => 62,
    15070 => 63,
    15071 => 63,
    15072 => 63,
    15073 => 63,
    15074 => 63,
    15075 => 63,
    15076 => 63,
    15077 => 63,
    15078 => 63,
    15079 => 63,
    15080 => 63,
    15081 => 63,
    15082 => 63,
    15083 => 63,
    15084 => 63,
    15085 => 63,
    15086 => 63,
    15087 => 63,
    15088 => 63,
    15089 => 63,
    15090 => 63,
    15091 => 63,
    15092 => 63,
    15093 => 63,
    15094 => 63,
    15095 => 63,
    15096 => 63,
    15097 => 63,
    15098 => 63,
    15099 => 63,
    15100 => 63,
    15101 => 63,
    15102 => 63,
    15103 => 63,
    15104 => 63,
    15105 => 63,
    15106 => 63,
    15107 => 63,
    15108 => 63,
    15109 => 63,
    15110 => 63,
    15111 => 63,
    15112 => 63,
    15113 => 63,
    15114 => 63,
    15115 => 63,
    15116 => 63,
    15117 => 63,
    15118 => 63,
    15119 => 63,
    15120 => 63,
    15121 => 63,
    15122 => 63,
    15123 => 63,
    15124 => 63,
    15125 => 63,
    15126 => 63,
    15127 => 63,
    15128 => 63,
    15129 => 63,
    15130 => 63,
    15131 => 63,
    15132 => 63,
    15133 => 63,
    15134 => 63,
    15135 => 63,
    15136 => 63,
    15137 => 63,
    15138 => 63,
    15139 => 63,
    15140 => 63,
    15141 => 63,
    15142 => 63,
    15143 => 63,
    15144 => 63,
    15145 => 63,
    15146 => 63,
    15147 => 63,
    15148 => 63,
    15149 => 63,
    15150 => 63,
    15151 => 63,
    15152 => 63,
    15153 => 63,
    15154 => 63,
    15155 => 63,
    15156 => 63,
    15157 => 63,
    15158 => 63,
    15159 => 63,
    15160 => 63,
    15161 => 63,
    15162 => 63,
    15163 => 63,
    15164 => 63,
    15165 => 63,
    15166 => 63,
    15167 => 63,
    15168 => 63,
    15169 => 63,
    15170 => 63,
    15171 => 63,
    15172 => 63,
    15173 => 63,
    15174 => 63,
    15175 => 63,
    15176 => 63,
    15177 => 63,
    15178 => 63,
    15179 => 63,
    15180 => 63,
    15181 => 63,
    15182 => 63,
    15183 => 63,
    15184 => 63,
    15185 => 63,
    15186 => 63,
    15187 => 63,
    15188 => 63,
    15189 => 63,
    15190 => 63,
    15191 => 63,
    15192 => 63,
    15193 => 63,
    15194 => 63,
    15195 => 63,
    15196 => 63,
    15197 => 63,
    15198 => 63,
    15199 => 63,
    15200 => 63,
    15201 => 63,
    15202 => 63,
    15203 => 63,
    15204 => 63,
    15205 => 63,
    15206 => 63,
    15207 => 63,
    15208 => 63,
    15209 => 63,
    15210 => 63,
    15211 => 63,
    15212 => 63,
    15213 => 63,
    15214 => 63,
    15215 => 63,
    15216 => 63,
    15217 => 63,
    15218 => 63,
    15219 => 63,
    15220 => 63,
    15221 => 63,
    15222 => 63,
    15223 => 63,
    15224 => 63,
    15225 => 63,
    15226 => 63,
    15227 => 63,
    15228 => 63,
    15229 => 63,
    15230 => 63,
    15231 => 63,
    15232 => 63,
    15233 => 63,
    15234 => 63,
    15235 => 63,
    15236 => 63,
    15237 => 63,
    15238 => 63,
    15239 => 63,
    15240 => 63,
    15241 => 63,
    15242 => 63,
    15243 => 63,
    15244 => 63,
    15245 => 63,
    15246 => 63,
    15247 => 63,
    15248 => 63,
    15249 => 63,
    15250 => 63,
    15251 => 63,
    15252 => 63,
    15253 => 63,
    15254 => 63,
    15255 => 63,
    15256 => 63,
    15257 => 63,
    15258 => 63,
    15259 => 63,
    15260 => 63,
    15261 => 63,
    15262 => 63,
    15263 => 63,
    15264 => 63,
    15265 => 63,
    15266 => 63,
    15267 => 63,
    15268 => 63,
    15269 => 63,
    15270 => 63,
    15271 => 63,
    15272 => 63,
    15273 => 63,
    15274 => 63,
    15275 => 63,
    15276 => 63,
    15277 => 63,
    15278 => 63,
    15279 => 63,
    15280 => 63,
    15281 => 63,
    15282 => 63,
    15283 => 63,
    15284 => 63,
    15285 => 63,
    15286 => 63,
    15287 => 63,
    15288 => 63,
    15289 => 63,
    15290 => 63,
    15291 => 63,
    15292 => 63,
    15293 => 63,
    15294 => 63,
    15295 => 63,
    15296 => 63,
    15297 => 63,
    15298 => 63,
    15299 => 63,
    15300 => 63,
    15301 => 63,
    15302 => 63,
    15303 => 63,
    15304 => 63,
    15305 => 63,
    15306 => 63,
    15307 => 63,
    15308 => 63,
    15309 => 63,
    15310 => 63,
    15311 => 63,
    15312 => 63,
    15313 => 63,
    15314 => 63,
    15315 => 63,
    15316 => 63,
    15317 => 63,
    15318 => 63,
    15319 => 63,
    15320 => 63,
    15321 => 63,
    15322 => 63,
    15323 => 63,
    15324 => 63,
    15325 => 63,
    15326 => 63,
    15327 => 63,
    15328 => 63,
    15329 => 63,
    15330 => 63,
    15331 => 63,
    15332 => 63,
    15333 => 63,
    15334 => 63,
    15335 => 63,
    15336 => 63,
    15337 => 63,
    15338 => 63,
    15339 => 63,
    15340 => 63,
    15341 => 63,
    15342 => 63,
    15343 => 63,
    15344 => 63,
    15345 => 63,
    15346 => 63,
    15347 => 63,
    15348 => 63,
    15349 => 63,
    15350 => 63,
    15351 => 63,
    15352 => 63,
    15353 => 63,
    15354 => 63,
    15355 => 63,
    15356 => 63,
    15357 => 63,
    15358 => 63,
    15359 => 63,
    15360 => 63,
    15361 => 63,
    15362 => 63,
    15363 => 63,
    15364 => 63,
    15365 => 63,
    15366 => 63,
    15367 => 63,
    15368 => 63,
    15369 => 63,
    15370 => 63,
    15371 => 63,
    15372 => 63,
    15373 => 63,
    15374 => 63,
    15375 => 63,
    15376 => 63,
    15377 => 63,
    15378 => 63,
    15379 => 63,
    15380 => 63,
    15381 => 63,
    15382 => 63,
    15383 => 63,
    15384 => 63,
    15385 => 63,
    15386 => 63,
    15387 => 63,
    15388 => 63,
    15389 => 63,
    15390 => 63,
    15391 => 63,
    15392 => 63,
    15393 => 63,
    15394 => 63,
    15395 => 63,
    15396 => 63,
    15397 => 63,
    15398 => 63,
    15399 => 63,
    15400 => 63,
    15401 => 63,
    15402 => 63,
    15403 => 63,
    15404 => 63,
    15405 => 63,
    15406 => 63,
    15407 => 63,
    15408 => 63,
    15409 => 63,
    15410 => 63,
    15411 => 63,
    15412 => 63,
    15413 => 63,
    15414 => 63,
    15415 => 63,
    15416 => 63,
    15417 => 63,
    15418 => 63,
    15419 => 63,
    15420 => 63,
    15421 => 63,
    15422 => 63,
    15423 => 63,
    15424 => 63,
    15425 => 63,
    15426 => 63,
    15427 => 63,
    15428 => 63,
    15429 => 63,
    15430 => 63,
    15431 => 63,
    15432 => 63,
    15433 => 63,
    15434 => 63,
    15435 => 63,
    15436 => 63,
    15437 => 63,
    15438 => 63,
    15439 => 63,
    15440 => 63,
    15441 => 63,
    15442 => 63,
    15443 => 63,
    15444 => 63,
    15445 => 63,
    15446 => 63,
    15447 => 63,
    15448 => 63,
    15449 => 63,
    15450 => 63,
    15451 => 63,
    15452 => 63,
    15453 => 63,
    15454 => 63,
    15455 => 63,
    15456 => 63,
    15457 => 63,
    15458 => 63,
    15459 => 63,
    15460 => 63,
    15461 => 63,
    15462 => 63,
    15463 => 63,
    15464 => 63,
    15465 => 63,
    15466 => 63,
    15467 => 63,
    15468 => 63,
    15469 => 63,
    15470 => 63,
    15471 => 63,
    15472 => 63,
    15473 => 63,
    15474 => 63,
    15475 => 63,
    15476 => 63,
    15477 => 63,
    15478 => 63,
    15479 => 63,
    15480 => 63,
    15481 => 63,
    15482 => 63,
    15483 => 63,
    15484 => 63,
    15485 => 63,
    15486 => 63,
    15487 => 63,
    15488 => 63,
    15489 => 63,
    15490 => 63,
    15491 => 63,
    15492 => 63,
    15493 => 63,
    15494 => 63,
    15495 => 63,
    15496 => 63,
    15497 => 63,
    15498 => 63,
    15499 => 63,
    15500 => 63,
    15501 => 63,
    15502 => 63,
    15503 => 63,
    15504 => 63,
    15505 => 63,
    15506 => 63,
    15507 => 63,
    15508 => 63,
    15509 => 63,
    15510 => 63,
    15511 => 63,
    15512 => 63,
    15513 => 63,
    15514 => 63,
    15515 => 63,
    15516 => 63,
    15517 => 63,
    15518 => 63,
    15519 => 63,
    15520 => 63,
    15521 => 63,
    15522 => 63,
    15523 => 63,
    15524 => 63,
    15525 => 63,
    15526 => 63,
    15527 => 63,
    15528 => 63,
    15529 => 63,
    15530 => 63,
    15531 => 63,
    15532 => 63,
    15533 => 63,
    15534 => 63,
    15535 => 63,
    15536 => 63,
    15537 => 63,
    15538 => 63,
    15539 => 63,
    15540 => 63,
    15541 => 63,
    15542 => 63,
    15543 => 63,
    15544 => 63,
    15545 => 63,
    15546 => 63,
    15547 => 63,
    15548 => 63,
    15549 => 63,
    15550 => 63,
    15551 => 63,
    15552 => 63,
    15553 => 63,
    15554 => 63,
    15555 => 63,
    15556 => 63,
    15557 => 63,
    15558 => 63,
    15559 => 63,
    15560 => 63,
    15561 => 63,
    15562 => 63,
    15563 => 63,
    15564 => 63,
    15565 => 63,
    15566 => 63,
    15567 => 63,
    15568 => 63,
    15569 => 63,
    15570 => 63,
    15571 => 63,
    15572 => 63,
    15573 => 63,
    15574 => 63,
    15575 => 63,
    15576 => 63,
    15577 => 63,
    15578 => 63,
    15579 => 63,
    15580 => 63,
    15581 => 63,
    15582 => 63,
    15583 => 63,
    15584 => 63,
    15585 => 63,
    15586 => 63,
    15587 => 63,
    15588 => 63,
    15589 => 63,
    15590 => 63,
    15591 => 63,
    15592 => 63,
    15593 => 63,
    15594 => 63,
    15595 => 63,
    15596 => 63,
    15597 => 63,
    15598 => 63,
    15599 => 63,
    15600 => 63,
    15601 => 63,
    15602 => 63,
    15603 => 63,
    15604 => 63,
    15605 => 63,
    15606 => 63,
    15607 => 63,
    15608 => 63,
    15609 => 63,
    15610 => 63,
    15611 => 63,
    15612 => 63,
    15613 => 63,
    15614 => 63,
    15615 => 63,
    15616 => 63,
    15617 => 63,
    15618 => 63,
    15619 => 63,
    15620 => 63,
    15621 => 63,
    15622 => 63,
    15623 => 63,
    15624 => 63,
    15625 => 63,
    15626 => 63,
    15627 => 63,
    15628 => 63,
    15629 => 63,
    15630 => 63,
    15631 => 63,
    15632 => 63,
    15633 => 63,
    15634 => 63,
    15635 => 63,
    15636 => 63,
    15637 => 63,
    15638 => 63,
    15639 => 63,
    15640 => 63,
    15641 => 63,
    15642 => 63,
    15643 => 63,
    15644 => 63,
    15645 => 63,
    15646 => 63,
    15647 => 63,
    15648 => 63,
    15649 => 63,
    15650 => 63,
    15651 => 63,
    15652 => 63,
    15653 => 63,
    15654 => 63,
    15655 => 63,
    15656 => 63,
    15657 => 63,
    15658 => 63,
    15659 => 63,
    15660 => 63,
    15661 => 63,
    15662 => 63,
    15663 => 63,
    15664 => 63,
    15665 => 63,
    15666 => 63,
    15667 => 63,
    15668 => 63,
    15669 => 63,
    15670 => 63,
    15671 => 63,
    15672 => 63,
    15673 => 63,
    15674 => 63,
    15675 => 63,
    15676 => 63,
    15677 => 63,
    15678 => 63,
    15679 => 63,
    15680 => 63,
    15681 => 63,
    15682 => 63,
    15683 => 63,
    15684 => 63,
    15685 => 63,
    15686 => 63,
    15687 => 63,
    15688 => 63,
    15689 => 63,
    15690 => 63,
    15691 => 63,
    15692 => 63,
    15693 => 63,
    15694 => 63,
    15695 => 63,
    15696 => 63,
    15697 => 63,
    15698 => 63,
    15699 => 63,
    15700 => 63,
    15701 => 63,
    15702 => 63,
    15703 => 63,
    15704 => 63,
    15705 => 63,
    15706 => 63,
    15707 => 63,
    15708 => 63,
    15709 => 63,
    15710 => 63,
    15711 => 63,
    15712 => 63,
    15713 => 63,
    15714 => 63,
    15715 => 63,
    15716 => 63,
    15717 => 63,
    15718 => 63,
    15719 => 63,
    15720 => 63,
    15721 => 63,
    15722 => 63,
    15723 => 63,
    15724 => 63,
    15725 => 63,
    15726 => 63,
    15727 => 63,
    15728 => 63,
    15729 => 63,
    15730 => 63,
    15731 => 63,
    15732 => 63,
    15733 => 63,
    15734 => 63,
    15735 => 63,
    15736 => 63,
    15737 => 63,
    15738 => 63,
    15739 => 63,
    15740 => 63,
    15741 => 63,
    15742 => 63,
    15743 => 63,
    15744 => 63,
    15745 => 63,
    15746 => 63,
    15747 => 63,
    15748 => 63,
    15749 => 63,
    15750 => 63,
    15751 => 63,
    15752 => 63,
    15753 => 63,
    15754 => 63,
    15755 => 63,
    15756 => 63,
    15757 => 63,
    15758 => 63,
    15759 => 63,
    15760 => 63,
    15761 => 63,
    15762 => 63,
    15763 => 63,
    15764 => 63,
    15765 => 63,
    15766 => 63,
    15767 => 63,
    15768 => 63,
    15769 => 63,
    15770 => 63,
    15771 => 63,
    15772 => 63,
    15773 => 63,
    15774 => 63,
    15775 => 63,
    15776 => 63,
    15777 => 63,
    15778 => 63,
    15779 => 63,
    15780 => 63,
    15781 => 63,
    15782 => 63,
    15783 => 63,
    15784 => 63,
    15785 => 63,
    15786 => 63,
    15787 => 63,
    15788 => 63,
    15789 => 63,
    15790 => 63,
    15791 => 63,
    15792 => 63,
    15793 => 63,
    15794 => 63,
    15795 => 63,
    15796 => 63,
    15797 => 63,
    15798 => 63,
    15799 => 63,
    15800 => 63,
    15801 => 63,
    15802 => 63,
    15803 => 63,
    15804 => 63,
    15805 => 63,
    15806 => 63,
    15807 => 63,
    15808 => 63,
    15809 => 63,
    15810 => 63,
    15811 => 63,
    15812 => 63,
    15813 => 63,
    15814 => 63,
    15815 => 63,
    15816 => 63,
    15817 => 63,
    15818 => 63,
    15819 => 63,
    15820 => 63,
    15821 => 63,
    15822 => 63,
    15823 => 63,
    15824 => 63,
    15825 => 63,
    15826 => 63,
    15827 => 63,
    15828 => 63,
    15829 => 63,
    15830 => 63,
    15831 => 63,
    15832 => 63,
    15833 => 63,
    15834 => 63,
    15835 => 63,
    15836 => 63,
    15837 => 63,
    15838 => 63,
    15839 => 63,
    15840 => 63,
    15841 => 63,
    15842 => 63,
    15843 => 63,
    15844 => 63,
    15845 => 63,
    15846 => 63,
    15847 => 63,
    15848 => 63,
    15849 => 63,
    15850 => 63,
    15851 => 63,
    15852 => 63,
    15853 => 63,
    15854 => 63,
    15855 => 63,
    15856 => 63,
    15857 => 63,
    15858 => 63,
    15859 => 63,
    15860 => 63,
    15861 => 63,
    15862 => 63,
    15863 => 63,
    15864 => 63,
    15865 => 63,
    15866 => 63,
    15867 => 63,
    15868 => 63,
    15869 => 63,
    15870 => 63,
    15871 => 63,
    15872 => 63,
    15873 => 63,
    15874 => 63,
    15875 => 63,
    15876 => 63,
    15877 => 63,
    15878 => 63,
    15879 => 63,
    15880 => 63,
    15881 => 63,
    15882 => 63,
    15883 => 63,
    15884 => 63,
    15885 => 63,
    15886 => 63,
    15887 => 63,
    15888 => 63,
    15889 => 63,
    15890 => 63,
    15891 => 63,
    15892 => 63,
    15893 => 63,
    15894 => 63,
    15895 => 63,
    15896 => 63,
    15897 => 63,
    15898 => 63,
    15899 => 63,
    15900 => 63,
    15901 => 63,
    15902 => 63,
    15903 => 63,
    15904 => 63,
    15905 => 63,
    15906 => 63,
    15907 => 63,
    15908 => 63,
    15909 => 63,
    15910 => 63,
    15911 => 63,
    15912 => 63,
    15913 => 63,
    15914 => 63,
    15915 => 63,
    15916 => 63,
    15917 => 63,
    15918 => 63,
    15919 => 63,
    15920 => 63,
    15921 => 63,
    15922 => 63,
    15923 => 63,
    15924 => 63,
    15925 => 63,
    15926 => 63,
    15927 => 63,
    15928 => 63,
    15929 => 63,
    15930 => 63,
    15931 => 63,
    15932 => 63,
    15933 => 63,
    15934 => 63,
    15935 => 63,
    15936 => 63,
    15937 => 63,
    15938 => 63,
    15939 => 63,
    15940 => 63,
    15941 => 63,
    15942 => 63,
    15943 => 63,
    15944 => 63,
    15945 => 63,
    15946 => 63,
    15947 => 63,
    15948 => 63,
    15949 => 63,
    15950 => 63,
    15951 => 63,
    15952 => 63,
    15953 => 63,
    15954 => 63,
    15955 => 63,
    15956 => 63,
    15957 => 63,
    15958 => 63,
    15959 => 63,
    15960 => 63,
    15961 => 63,
    15962 => 63,
    15963 => 63,
    15964 => 63,
    15965 => 63,
    15966 => 63,
    15967 => 63,
    15968 => 63,
    15969 => 63,
    15970 => 63,
    15971 => 63,
    15972 => 63,
    15973 => 63,
    15974 => 63,
    15975 => 63,
    15976 => 63,
    15977 => 63,
    15978 => 63,
    15979 => 63,
    15980 => 63,
    15981 => 63,
    15982 => 63,
    15983 => 63,
    15984 => 63,
    15985 => 63,
    15986 => 63,
    15987 => 63,
    15988 => 63,
    15989 => 63,
    15990 => 63,
    15991 => 63,
    15992 => 63,
    15993 => 63,
    15994 => 63,
    15995 => 63,
    15996 => 63,
    15997 => 63,
    15998 => 63,
    15999 => 63,
    16000 => 63,
    16001 => 63,
    16002 => 63,
    16003 => 63,
    16004 => 63,
    16005 => 63,
    16006 => 63,
    16007 => 63,
    16008 => 63,
    16009 => 63,
    16010 => 63,
    16011 => 63,
    16012 => 63,
    16013 => 63,
    16014 => 63,
    16015 => 63,
    16016 => 63,
    16017 => 63,
    16018 => 63,
    16019 => 63,
    16020 => 63,
    16021 => 63,
    16022 => 63,
    16023 => 63,
    16024 => 63,
    16025 => 63,
    16026 => 63,
    16027 => 63,
    16028 => 63,
    16029 => 63,
    16030 => 63,
    16031 => 63,
    16032 => 63,
    16033 => 63,
    16034 => 63,
    16035 => 63,
    16036 => 63,
    16037 => 63,
    16038 => 63,
    16039 => 63,
    16040 => 63,
    16041 => 63,
    16042 => 63,
    16043 => 63,
    16044 => 63,
    16045 => 63,
    16046 => 63,
    16047 => 63,
    16048 => 63,
    16049 => 63,
    16050 => 63,
    16051 => 63,
    16052 => 63,
    16053 => 63,
    16054 => 63,
    16055 => 63,
    16056 => 63,
    16057 => 63,
    16058 => 63,
    16059 => 63,
    16060 => 63,
    16061 => 63,
    16062 => 63,
    16063 => 63,
    16064 => 63,
    16065 => 63,
    16066 => 63,
    16067 => 63,
    16068 => 63,
    16069 => 63,
    16070 => 63,
    16071 => 63,
    16072 => 63,
    16073 => 63,
    16074 => 63,
    16075 => 63,
    16076 => 63,
    16077 => 63,
    16078 => 63,
    16079 => 63,
    16080 => 63,
    16081 => 63,
    16082 => 63,
    16083 => 63,
    16084 => 63,
    16085 => 63,
    16086 => 63,
    16087 => 63,
    16088 => 63,
    16089 => 63,
    16090 => 63,
    16091 => 63,
    16092 => 63,
    16093 => 63,
    16094 => 63,
    16095 => 63,
    16096 => 63,
    16097 => 63,
    16098 => 63,
    16099 => 63,
    16100 => 63,
    16101 => 63,
    16102 => 63,
    16103 => 63,
    16104 => 63,
    16105 => 63,
    16106 => 63,
    16107 => 63,
    16108 => 63,
    16109 => 63,
    16110 => 63,
    16111 => 63,
    16112 => 63,
    16113 => 63,
    16114 => 63,
    16115 => 63,
    16116 => 63,
    16117 => 63,
    16118 => 63,
    16119 => 63,
    16120 => 63,
    16121 => 63,
    16122 => 63,
    16123 => 63,
    16124 => 63,
    16125 => 63,
    16126 => 63,
    16127 => 63,
    16128 => 63,
    16129 => 63,
    16130 => 63,
    16131 => 63,
    16132 => 63,
    16133 => 63,
    16134 => 63,
    16135 => 63,
    16136 => 63,
    16137 => 63,
    16138 => 63,
    16139 => 63,
    16140 => 63,
    16141 => 63,
    16142 => 63,
    16143 => 63,
    16144 => 63,
    16145 => 63,
    16146 => 63,
    16147 => 63,
    16148 => 63,
    16149 => 63,
    16150 => 63,
    16151 => 63,
    16152 => 63,
    16153 => 63,
    16154 => 63,
    16155 => 63,
    16156 => 63,
    16157 => 63,
    16158 => 63,
    16159 => 63,
    16160 => 63,
    16161 => 63,
    16162 => 63,
    16163 => 63,
    16164 => 63,
    16165 => 63,
    16166 => 63,
    16167 => 63,
    16168 => 63,
    16169 => 63,
    16170 => 63,
    16171 => 63,
    16172 => 63,
    16173 => 63,
    16174 => 63,
    16175 => 63,
    16176 => 63,
    16177 => 63,
    16178 => 63,
    16179 => 63,
    16180 => 63,
    16181 => 63,
    16182 => 63,
    16183 => 63,
    16184 => 63,
    16185 => 63,
    16186 => 63,
    16187 => 63,
    16188 => 63,
    16189 => 63,
    16190 => 63,
    16191 => 63,
    16192 => 63,
    16193 => 63,
    16194 => 63,
    16195 => 63,
    16196 => 63,
    16197 => 63,
    16198 => 63,
    16199 => 63,
    16200 => 63,
    16201 => 63,
    16202 => 63,
    16203 => 63,
    16204 => 63,
    16205 => 63,
    16206 => 63,
    16207 => 63,
    16208 => 63,
    16209 => 63,
    16210 => 63,
    16211 => 63,
    16212 => 63,
    16213 => 63,
    16214 => 63,
    16215 => 63,
    16216 => 63,
    16217 => 63,
    16218 => 63,
    16219 => 63,
    16220 => 63,
    16221 => 63,
    16222 => 63,
    16223 => 63,
    16224 => 63,
    16225 => 63,
    16226 => 63,
    16227 => 63,
    16228 => 63,
    16229 => 63,
    16230 => 63,
    16231 => 63,
    16232 => 63,
    16233 => 63,
    16234 => 63,
    16235 => 63,
    16236 => 63,
    16237 => 63,
    16238 => 63,
    16239 => 63,
    16240 => 63,
    16241 => 63,
    16242 => 63,
    16243 => 63,
    16244 => 63,
    16245 => 63,
    16246 => 63,
    16247 => 63,
    16248 => 63,
    16249 => 63,
    16250 => 63,
    16251 => 63,
    16252 => 63,
    16253 => 63,
    16254 => 63,
    16255 => 63,
    16256 => 63,
    16257 => 63,
    16258 => 63,
    16259 => 63,
    16260 => 63,
    16261 => 63,
    16262 => 63,
    16263 => 63,
    16264 => 63,
    16265 => 63,
    16266 => 63,
    16267 => 63,
    16268 => 63,
    16269 => 63,
    16270 => 63,
    16271 => 63,
    16272 => 63,
    16273 => 63,
    16274 => 63,
    16275 => 63,
    16276 => 63,
    16277 => 63,
    16278 => 63,
    16279 => 63,
    16280 => 63,
    16281 => 63,
    16282 => 63,
    16283 => 63,
    16284 => 63,
    16285 => 63,
    16286 => 63,
    16287 => 63,
    16288 => 63,
    16289 => 63,
    16290 => 63,
    16291 => 63,
    16292 => 63,
    16293 => 63,
    16294 => 63,
    16295 => 63,
    16296 => 63,
    16297 => 63,
    16298 => 63,
    16299 => 63,
    16300 => 63,
    16301 => 63,
    16302 => 63,
    16303 => 63,
    16304 => 63,
    16305 => 63,
    16306 => 63,
    16307 => 63,
    16308 => 63,
    16309 => 63,
    16310 => 63,
    16311 => 63,
    16312 => 63,
    16313 => 63,
    16314 => 63,
    16315 => 63,
    16316 => 63,
    16317 => 63,
    16318 => 63,
    16319 => 63,
    16320 => 63,
    16321 => 63,
    16322 => 63,
    16323 => 63,
    16324 => 63,
    16325 => 63,
    16326 => 63,
    16327 => 63,
    16328 => 63,
    16329 => 63,
    16330 => 63,
    16331 => 63,
    16332 => 63,
    16333 => 63,
    16334 => 63,
    16335 => 63,
    16336 => 63,
    16337 => 63,
    16338 => 63,
    16339 => 63,
    16340 => 63,
    16341 => 63,
    16342 => 63,
    16343 => 63,
    16344 => 63,
    16345 => 63,
    16346 => 63,
    16347 => 63,
    16348 => 63,
    16349 => 63,
    16350 => 63,
    16351 => 63,
    16352 => 63,
    16353 => 63,
    16354 => 63,
    16355 => 63,
    16356 => 63,
    16357 => 63,
    16358 => 63,
    16359 => 63,
    16360 => 63,
    16361 => 63,
    16362 => 63,
    16363 => 63,
    16364 => 63,
    16365 => 63,
    16366 => 63,
    16367 => 63,
    16368 => 63,
    16369 => 63,
    16370 => 63,
    16371 => 63,
    16372 => 63,
    16373 => 63,
    16374 => 63,
    16375 => 63,
    16376 => 63,
    16377 => 63,
    16378 => 63,
    16379 => 63,
    16380 => 63,
    16381 => 63,
    16382 => 63,
    16383 => 63
  );

  begin
    -- Process to output LUT data based on address input
    lut_out <= std_logic_vector(to_signed(LUT(to_integer(unsigned(address))), P));
  end architecture;
