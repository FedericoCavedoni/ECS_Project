library IEEE;
  use IEEE.std_logic_1164.all;
  use IEEE.numeric_std.all;

entity lut_table_65536_7bit is
  generic (
    N : integer := 16;
    P : integer := 7
  );
  port (
    address  : in  std_logic_vector(N-1 downto 0);
    lut_out : out std_logic_vector(P-1 downto 0)
  );
end entity;

architecture behavior of lut_table_65536_7bit is

  type LUT_t is array (natural range 0 to 65535) of integer;
  constant LUT: LUT_t := (
    0 => 0,
    1 => 0,
    2 => 0,
    3 => 0,
    4 => 0,
    5 => 0,
    6 => 0,
    7 => 0,
    8 => 0,
    9 => 0,
    10 => 0,
    11 => 0,
    12 => 0,
    13 => 0,
    14 => 0,
    15 => 0,
    16 => 0,
    17 => 0,
    18 => 0,
    19 => 0,
    20 => 0,
    21 => 0,
    22 => 0,
    23 => 0,
    24 => 0,
    25 => 0,
    26 => 0,
    27 => 0,
    28 => 0,
    29 => 0,
    30 => 0,
    31 => 0,
    32 => 0,
    33 => 0,
    34 => 0,
    35 => 0,
    36 => 0,
    37 => 0,
    38 => 0,
    39 => 0,
    40 => 0,
    41 => 0,
    42 => 0,
    43 => 0,
    44 => 0,
    45 => 0,
    46 => 0,
    47 => 0,
    48 => 0,
    49 => 0,
    50 => 0,
    51 => 0,
    52 => 0,
    53 => 0,
    54 => 0,
    55 => 0,
    56 => 0,
    57 => 0,
    58 => 0,
    59 => 0,
    60 => 0,
    61 => 0,
    62 => 0,
    63 => 0,
    64 => 0,
    65 => 0,
    66 => 0,
    67 => 0,
    68 => 0,
    69 => 0,
    70 => 0,
    71 => 0,
    72 => 0,
    73 => 0,
    74 => 0,
    75 => 0,
    76 => 0,
    77 => 0,
    78 => 0,
    79 => 0,
    80 => 0,
    81 => 0,
    82 => 0,
    83 => 1,
    84 => 1,
    85 => 1,
    86 => 1,
    87 => 1,
    88 => 1,
    89 => 1,
    90 => 1,
    91 => 1,
    92 => 1,
    93 => 1,
    94 => 1,
    95 => 1,
    96 => 1,
    97 => 1,
    98 => 1,
    99 => 1,
    100 => 1,
    101 => 1,
    102 => 1,
    103 => 1,
    104 => 1,
    105 => 1,
    106 => 1,
    107 => 1,
    108 => 1,
    109 => 1,
    110 => 1,
    111 => 1,
    112 => 1,
    113 => 1,
    114 => 1,
    115 => 1,
    116 => 1,
    117 => 1,
    118 => 1,
    119 => 1,
    120 => 1,
    121 => 1,
    122 => 1,
    123 => 1,
    124 => 1,
    125 => 1,
    126 => 1,
    127 => 1,
    128 => 1,
    129 => 1,
    130 => 1,
    131 => 1,
    132 => 1,
    133 => 1,
    134 => 1,
    135 => 1,
    136 => 1,
    137 => 1,
    138 => 1,
    139 => 1,
    140 => 1,
    141 => 1,
    142 => 1,
    143 => 1,
    144 => 1,
    145 => 1,
    146 => 1,
    147 => 1,
    148 => 1,
    149 => 1,
    150 => 1,
    151 => 1,
    152 => 1,
    153 => 1,
    154 => 1,
    155 => 1,
    156 => 1,
    157 => 1,
    158 => 1,
    159 => 1,
    160 => 1,
    161 => 1,
    162 => 1,
    163 => 1,
    164 => 1,
    165 => 1,
    166 => 1,
    167 => 1,
    168 => 1,
    169 => 1,
    170 => 1,
    171 => 1,
    172 => 1,
    173 => 1,
    174 => 1,
    175 => 1,
    176 => 1,
    177 => 1,
    178 => 1,
    179 => 1,
    180 => 1,
    181 => 1,
    182 => 1,
    183 => 1,
    184 => 1,
    185 => 1,
    186 => 1,
    187 => 1,
    188 => 1,
    189 => 1,
    190 => 1,
    191 => 1,
    192 => 1,
    193 => 1,
    194 => 1,
    195 => 1,
    196 => 1,
    197 => 1,
    198 => 1,
    199 => 1,
    200 => 1,
    201 => 1,
    202 => 1,
    203 => 1,
    204 => 1,
    205 => 1,
    206 => 1,
    207 => 1,
    208 => 1,
    209 => 1,
    210 => 1,
    211 => 1,
    212 => 1,
    213 => 1,
    214 => 1,
    215 => 1,
    216 => 1,
    217 => 1,
    218 => 1,
    219 => 1,
    220 => 1,
    221 => 1,
    222 => 1,
    223 => 1,
    224 => 1,
    225 => 1,
    226 => 1,
    227 => 1,
    228 => 1,
    229 => 1,
    230 => 1,
    231 => 1,
    232 => 1,
    233 => 1,
    234 => 1,
    235 => 1,
    236 => 1,
    237 => 1,
    238 => 1,
    239 => 1,
    240 => 1,
    241 => 1,
    242 => 1,
    243 => 1,
    244 => 1,
    245 => 1,
    246 => 1,
    247 => 1,
    248 => 1,
    249 => 2,
    250 => 2,
    251 => 2,
    252 => 2,
    253 => 2,
    254 => 2,
    255 => 2,
    256 => 2,
    257 => 2,
    258 => 2,
    259 => 2,
    260 => 2,
    261 => 2,
    262 => 2,
    263 => 2,
    264 => 2,
    265 => 2,
    266 => 2,
    267 => 2,
    268 => 2,
    269 => 2,
    270 => 2,
    271 => 2,
    272 => 2,
    273 => 2,
    274 => 2,
    275 => 2,
    276 => 2,
    277 => 2,
    278 => 2,
    279 => 2,
    280 => 2,
    281 => 2,
    282 => 2,
    283 => 2,
    284 => 2,
    285 => 2,
    286 => 2,
    287 => 2,
    288 => 2,
    289 => 2,
    290 => 2,
    291 => 2,
    292 => 2,
    293 => 2,
    294 => 2,
    295 => 2,
    296 => 2,
    297 => 2,
    298 => 2,
    299 => 2,
    300 => 2,
    301 => 2,
    302 => 2,
    303 => 2,
    304 => 2,
    305 => 2,
    306 => 2,
    307 => 2,
    308 => 2,
    309 => 2,
    310 => 2,
    311 => 2,
    312 => 2,
    313 => 2,
    314 => 2,
    315 => 2,
    316 => 2,
    317 => 2,
    318 => 2,
    319 => 2,
    320 => 2,
    321 => 2,
    322 => 2,
    323 => 2,
    324 => 2,
    325 => 2,
    326 => 2,
    327 => 2,
    328 => 2,
    329 => 2,
    330 => 2,
    331 => 2,
    332 => 2,
    333 => 2,
    334 => 2,
    335 => 2,
    336 => 2,
    337 => 2,
    338 => 2,
    339 => 2,
    340 => 2,
    341 => 2,
    342 => 2,
    343 => 2,
    344 => 2,
    345 => 2,
    346 => 2,
    347 => 2,
    348 => 2,
    349 => 2,
    350 => 2,
    351 => 2,
    352 => 2,
    353 => 2,
    354 => 2,
    355 => 2,
    356 => 2,
    357 => 2,
    358 => 2,
    359 => 2,
    360 => 2,
    361 => 2,
    362 => 2,
    363 => 2,
    364 => 2,
    365 => 2,
    366 => 2,
    367 => 2,
    368 => 2,
    369 => 2,
    370 => 2,
    371 => 2,
    372 => 2,
    373 => 2,
    374 => 2,
    375 => 2,
    376 => 2,
    377 => 2,
    378 => 2,
    379 => 2,
    380 => 2,
    381 => 2,
    382 => 2,
    383 => 2,
    384 => 2,
    385 => 2,
    386 => 2,
    387 => 2,
    388 => 2,
    389 => 2,
    390 => 2,
    391 => 2,
    392 => 2,
    393 => 2,
    394 => 2,
    395 => 2,
    396 => 2,
    397 => 2,
    398 => 2,
    399 => 2,
    400 => 2,
    401 => 2,
    402 => 2,
    403 => 2,
    404 => 2,
    405 => 2,
    406 => 2,
    407 => 2,
    408 => 2,
    409 => 2,
    410 => 2,
    411 => 2,
    412 => 2,
    413 => 2,
    414 => 2,
    415 => 3,
    416 => 3,
    417 => 3,
    418 => 3,
    419 => 3,
    420 => 3,
    421 => 3,
    422 => 3,
    423 => 3,
    424 => 3,
    425 => 3,
    426 => 3,
    427 => 3,
    428 => 3,
    429 => 3,
    430 => 3,
    431 => 3,
    432 => 3,
    433 => 3,
    434 => 3,
    435 => 3,
    436 => 3,
    437 => 3,
    438 => 3,
    439 => 3,
    440 => 3,
    441 => 3,
    442 => 3,
    443 => 3,
    444 => 3,
    445 => 3,
    446 => 3,
    447 => 3,
    448 => 3,
    449 => 3,
    450 => 3,
    451 => 3,
    452 => 3,
    453 => 3,
    454 => 3,
    455 => 3,
    456 => 3,
    457 => 3,
    458 => 3,
    459 => 3,
    460 => 3,
    461 => 3,
    462 => 3,
    463 => 3,
    464 => 3,
    465 => 3,
    466 => 3,
    467 => 3,
    468 => 3,
    469 => 3,
    470 => 3,
    471 => 3,
    472 => 3,
    473 => 3,
    474 => 3,
    475 => 3,
    476 => 3,
    477 => 3,
    478 => 3,
    479 => 3,
    480 => 3,
    481 => 3,
    482 => 3,
    483 => 3,
    484 => 3,
    485 => 3,
    486 => 3,
    487 => 3,
    488 => 3,
    489 => 3,
    490 => 3,
    491 => 3,
    492 => 3,
    493 => 3,
    494 => 3,
    495 => 3,
    496 => 3,
    497 => 3,
    498 => 3,
    499 => 3,
    500 => 3,
    501 => 3,
    502 => 3,
    503 => 3,
    504 => 3,
    505 => 3,
    506 => 3,
    507 => 3,
    508 => 3,
    509 => 3,
    510 => 3,
    511 => 3,
    512 => 3,
    513 => 3,
    514 => 3,
    515 => 3,
    516 => 3,
    517 => 3,
    518 => 3,
    519 => 3,
    520 => 3,
    521 => 3,
    522 => 3,
    523 => 3,
    524 => 3,
    525 => 3,
    526 => 3,
    527 => 3,
    528 => 3,
    529 => 3,
    530 => 3,
    531 => 3,
    532 => 3,
    533 => 3,
    534 => 3,
    535 => 3,
    536 => 3,
    537 => 3,
    538 => 3,
    539 => 3,
    540 => 3,
    541 => 3,
    542 => 3,
    543 => 3,
    544 => 3,
    545 => 3,
    546 => 3,
    547 => 3,
    548 => 3,
    549 => 3,
    550 => 3,
    551 => 3,
    552 => 3,
    553 => 3,
    554 => 3,
    555 => 3,
    556 => 3,
    557 => 3,
    558 => 3,
    559 => 3,
    560 => 3,
    561 => 3,
    562 => 3,
    563 => 3,
    564 => 3,
    565 => 3,
    566 => 3,
    567 => 3,
    568 => 3,
    569 => 3,
    570 => 3,
    571 => 3,
    572 => 3,
    573 => 3,
    574 => 3,
    575 => 3,
    576 => 3,
    577 => 3,
    578 => 3,
    579 => 3,
    580 => 4,
    581 => 4,
    582 => 4,
    583 => 4,
    584 => 4,
    585 => 4,
    586 => 4,
    587 => 4,
    588 => 4,
    589 => 4,
    590 => 4,
    591 => 4,
    592 => 4,
    593 => 4,
    594 => 4,
    595 => 4,
    596 => 4,
    597 => 4,
    598 => 4,
    599 => 4,
    600 => 4,
    601 => 4,
    602 => 4,
    603 => 4,
    604 => 4,
    605 => 4,
    606 => 4,
    607 => 4,
    608 => 4,
    609 => 4,
    610 => 4,
    611 => 4,
    612 => 4,
    613 => 4,
    614 => 4,
    615 => 4,
    616 => 4,
    617 => 4,
    618 => 4,
    619 => 4,
    620 => 4,
    621 => 4,
    622 => 4,
    623 => 4,
    624 => 4,
    625 => 4,
    626 => 4,
    627 => 4,
    628 => 4,
    629 => 4,
    630 => 4,
    631 => 4,
    632 => 4,
    633 => 4,
    634 => 4,
    635 => 4,
    636 => 4,
    637 => 4,
    638 => 4,
    639 => 4,
    640 => 4,
    641 => 4,
    642 => 4,
    643 => 4,
    644 => 4,
    645 => 4,
    646 => 4,
    647 => 4,
    648 => 4,
    649 => 4,
    650 => 4,
    651 => 4,
    652 => 4,
    653 => 4,
    654 => 4,
    655 => 4,
    656 => 4,
    657 => 4,
    658 => 4,
    659 => 4,
    660 => 4,
    661 => 4,
    662 => 4,
    663 => 4,
    664 => 4,
    665 => 4,
    666 => 4,
    667 => 4,
    668 => 4,
    669 => 4,
    670 => 4,
    671 => 4,
    672 => 4,
    673 => 4,
    674 => 4,
    675 => 4,
    676 => 4,
    677 => 4,
    678 => 4,
    679 => 4,
    680 => 4,
    681 => 4,
    682 => 4,
    683 => 4,
    684 => 4,
    685 => 4,
    686 => 4,
    687 => 4,
    688 => 4,
    689 => 4,
    690 => 4,
    691 => 4,
    692 => 4,
    693 => 4,
    694 => 4,
    695 => 4,
    696 => 4,
    697 => 4,
    698 => 4,
    699 => 4,
    700 => 4,
    701 => 4,
    702 => 4,
    703 => 4,
    704 => 4,
    705 => 4,
    706 => 4,
    707 => 4,
    708 => 4,
    709 => 4,
    710 => 4,
    711 => 4,
    712 => 4,
    713 => 4,
    714 => 4,
    715 => 4,
    716 => 4,
    717 => 4,
    718 => 4,
    719 => 4,
    720 => 4,
    721 => 4,
    722 => 4,
    723 => 4,
    724 => 4,
    725 => 4,
    726 => 4,
    727 => 4,
    728 => 4,
    729 => 4,
    730 => 4,
    731 => 4,
    732 => 4,
    733 => 4,
    734 => 4,
    735 => 4,
    736 => 4,
    737 => 4,
    738 => 4,
    739 => 4,
    740 => 4,
    741 => 4,
    742 => 4,
    743 => 4,
    744 => 4,
    745 => 4,
    746 => 5,
    747 => 5,
    748 => 5,
    749 => 5,
    750 => 5,
    751 => 5,
    752 => 5,
    753 => 5,
    754 => 5,
    755 => 5,
    756 => 5,
    757 => 5,
    758 => 5,
    759 => 5,
    760 => 5,
    761 => 5,
    762 => 5,
    763 => 5,
    764 => 5,
    765 => 5,
    766 => 5,
    767 => 5,
    768 => 5,
    769 => 5,
    770 => 5,
    771 => 5,
    772 => 5,
    773 => 5,
    774 => 5,
    775 => 5,
    776 => 5,
    777 => 5,
    778 => 5,
    779 => 5,
    780 => 5,
    781 => 5,
    782 => 5,
    783 => 5,
    784 => 5,
    785 => 5,
    786 => 5,
    787 => 5,
    788 => 5,
    789 => 5,
    790 => 5,
    791 => 5,
    792 => 5,
    793 => 5,
    794 => 5,
    795 => 5,
    796 => 5,
    797 => 5,
    798 => 5,
    799 => 5,
    800 => 5,
    801 => 5,
    802 => 5,
    803 => 5,
    804 => 5,
    805 => 5,
    806 => 5,
    807 => 5,
    808 => 5,
    809 => 5,
    810 => 5,
    811 => 5,
    812 => 5,
    813 => 5,
    814 => 5,
    815 => 5,
    816 => 5,
    817 => 5,
    818 => 5,
    819 => 5,
    820 => 5,
    821 => 5,
    822 => 5,
    823 => 5,
    824 => 5,
    825 => 5,
    826 => 5,
    827 => 5,
    828 => 5,
    829 => 5,
    830 => 5,
    831 => 5,
    832 => 5,
    833 => 5,
    834 => 5,
    835 => 5,
    836 => 5,
    837 => 5,
    838 => 5,
    839 => 5,
    840 => 5,
    841 => 5,
    842 => 5,
    843 => 5,
    844 => 5,
    845 => 5,
    846 => 5,
    847 => 5,
    848 => 5,
    849 => 5,
    850 => 5,
    851 => 5,
    852 => 5,
    853 => 5,
    854 => 5,
    855 => 5,
    856 => 5,
    857 => 5,
    858 => 5,
    859 => 5,
    860 => 5,
    861 => 5,
    862 => 5,
    863 => 5,
    864 => 5,
    865 => 5,
    866 => 5,
    867 => 5,
    868 => 5,
    869 => 5,
    870 => 5,
    871 => 5,
    872 => 5,
    873 => 5,
    874 => 5,
    875 => 5,
    876 => 5,
    877 => 5,
    878 => 5,
    879 => 5,
    880 => 5,
    881 => 5,
    882 => 5,
    883 => 5,
    884 => 5,
    885 => 5,
    886 => 5,
    887 => 5,
    888 => 5,
    889 => 5,
    890 => 5,
    891 => 5,
    892 => 5,
    893 => 5,
    894 => 5,
    895 => 5,
    896 => 5,
    897 => 5,
    898 => 5,
    899 => 5,
    900 => 5,
    901 => 5,
    902 => 5,
    903 => 5,
    904 => 5,
    905 => 5,
    906 => 5,
    907 => 5,
    908 => 5,
    909 => 5,
    910 => 5,
    911 => 5,
    912 => 6,
    913 => 6,
    914 => 6,
    915 => 6,
    916 => 6,
    917 => 6,
    918 => 6,
    919 => 6,
    920 => 6,
    921 => 6,
    922 => 6,
    923 => 6,
    924 => 6,
    925 => 6,
    926 => 6,
    927 => 6,
    928 => 6,
    929 => 6,
    930 => 6,
    931 => 6,
    932 => 6,
    933 => 6,
    934 => 6,
    935 => 6,
    936 => 6,
    937 => 6,
    938 => 6,
    939 => 6,
    940 => 6,
    941 => 6,
    942 => 6,
    943 => 6,
    944 => 6,
    945 => 6,
    946 => 6,
    947 => 6,
    948 => 6,
    949 => 6,
    950 => 6,
    951 => 6,
    952 => 6,
    953 => 6,
    954 => 6,
    955 => 6,
    956 => 6,
    957 => 6,
    958 => 6,
    959 => 6,
    960 => 6,
    961 => 6,
    962 => 6,
    963 => 6,
    964 => 6,
    965 => 6,
    966 => 6,
    967 => 6,
    968 => 6,
    969 => 6,
    970 => 6,
    971 => 6,
    972 => 6,
    973 => 6,
    974 => 6,
    975 => 6,
    976 => 6,
    977 => 6,
    978 => 6,
    979 => 6,
    980 => 6,
    981 => 6,
    982 => 6,
    983 => 6,
    984 => 6,
    985 => 6,
    986 => 6,
    987 => 6,
    988 => 6,
    989 => 6,
    990 => 6,
    991 => 6,
    992 => 6,
    993 => 6,
    994 => 6,
    995 => 6,
    996 => 6,
    997 => 6,
    998 => 6,
    999 => 6,
    1000 => 6,
    1001 => 6,
    1002 => 6,
    1003 => 6,
    1004 => 6,
    1005 => 6,
    1006 => 6,
    1007 => 6,
    1008 => 6,
    1009 => 6,
    1010 => 6,
    1011 => 6,
    1012 => 6,
    1013 => 6,
    1014 => 6,
    1015 => 6,
    1016 => 6,
    1017 => 6,
    1018 => 6,
    1019 => 6,
    1020 => 6,
    1021 => 6,
    1022 => 6,
    1023 => 6,
    1024 => 6,
    1025 => 6,
    1026 => 6,
    1027 => 6,
    1028 => 6,
    1029 => 6,
    1030 => 6,
    1031 => 6,
    1032 => 6,
    1033 => 6,
    1034 => 6,
    1035 => 6,
    1036 => 6,
    1037 => 6,
    1038 => 6,
    1039 => 6,
    1040 => 6,
    1041 => 6,
    1042 => 6,
    1043 => 6,
    1044 => 6,
    1045 => 6,
    1046 => 6,
    1047 => 6,
    1048 => 6,
    1049 => 6,
    1050 => 6,
    1051 => 6,
    1052 => 6,
    1053 => 6,
    1054 => 6,
    1055 => 6,
    1056 => 6,
    1057 => 6,
    1058 => 6,
    1059 => 6,
    1060 => 6,
    1061 => 6,
    1062 => 6,
    1063 => 6,
    1064 => 6,
    1065 => 6,
    1066 => 6,
    1067 => 6,
    1068 => 6,
    1069 => 6,
    1070 => 6,
    1071 => 6,
    1072 => 6,
    1073 => 6,
    1074 => 6,
    1075 => 6,
    1076 => 6,
    1077 => 6,
    1078 => 6,
    1079 => 7,
    1080 => 7,
    1081 => 7,
    1082 => 7,
    1083 => 7,
    1084 => 7,
    1085 => 7,
    1086 => 7,
    1087 => 7,
    1088 => 7,
    1089 => 7,
    1090 => 7,
    1091 => 7,
    1092 => 7,
    1093 => 7,
    1094 => 7,
    1095 => 7,
    1096 => 7,
    1097 => 7,
    1098 => 7,
    1099 => 7,
    1100 => 7,
    1101 => 7,
    1102 => 7,
    1103 => 7,
    1104 => 7,
    1105 => 7,
    1106 => 7,
    1107 => 7,
    1108 => 7,
    1109 => 7,
    1110 => 7,
    1111 => 7,
    1112 => 7,
    1113 => 7,
    1114 => 7,
    1115 => 7,
    1116 => 7,
    1117 => 7,
    1118 => 7,
    1119 => 7,
    1120 => 7,
    1121 => 7,
    1122 => 7,
    1123 => 7,
    1124 => 7,
    1125 => 7,
    1126 => 7,
    1127 => 7,
    1128 => 7,
    1129 => 7,
    1130 => 7,
    1131 => 7,
    1132 => 7,
    1133 => 7,
    1134 => 7,
    1135 => 7,
    1136 => 7,
    1137 => 7,
    1138 => 7,
    1139 => 7,
    1140 => 7,
    1141 => 7,
    1142 => 7,
    1143 => 7,
    1144 => 7,
    1145 => 7,
    1146 => 7,
    1147 => 7,
    1148 => 7,
    1149 => 7,
    1150 => 7,
    1151 => 7,
    1152 => 7,
    1153 => 7,
    1154 => 7,
    1155 => 7,
    1156 => 7,
    1157 => 7,
    1158 => 7,
    1159 => 7,
    1160 => 7,
    1161 => 7,
    1162 => 7,
    1163 => 7,
    1164 => 7,
    1165 => 7,
    1166 => 7,
    1167 => 7,
    1168 => 7,
    1169 => 7,
    1170 => 7,
    1171 => 7,
    1172 => 7,
    1173 => 7,
    1174 => 7,
    1175 => 7,
    1176 => 7,
    1177 => 7,
    1178 => 7,
    1179 => 7,
    1180 => 7,
    1181 => 7,
    1182 => 7,
    1183 => 7,
    1184 => 7,
    1185 => 7,
    1186 => 7,
    1187 => 7,
    1188 => 7,
    1189 => 7,
    1190 => 7,
    1191 => 7,
    1192 => 7,
    1193 => 7,
    1194 => 7,
    1195 => 7,
    1196 => 7,
    1197 => 7,
    1198 => 7,
    1199 => 7,
    1200 => 7,
    1201 => 7,
    1202 => 7,
    1203 => 7,
    1204 => 7,
    1205 => 7,
    1206 => 7,
    1207 => 7,
    1208 => 7,
    1209 => 7,
    1210 => 7,
    1211 => 7,
    1212 => 7,
    1213 => 7,
    1214 => 7,
    1215 => 7,
    1216 => 7,
    1217 => 7,
    1218 => 7,
    1219 => 7,
    1220 => 7,
    1221 => 7,
    1222 => 7,
    1223 => 7,
    1224 => 7,
    1225 => 7,
    1226 => 7,
    1227 => 7,
    1228 => 7,
    1229 => 7,
    1230 => 7,
    1231 => 7,
    1232 => 7,
    1233 => 7,
    1234 => 7,
    1235 => 7,
    1236 => 7,
    1237 => 7,
    1238 => 7,
    1239 => 7,
    1240 => 7,
    1241 => 7,
    1242 => 7,
    1243 => 7,
    1244 => 7,
    1245 => 8,
    1246 => 8,
    1247 => 8,
    1248 => 8,
    1249 => 8,
    1250 => 8,
    1251 => 8,
    1252 => 8,
    1253 => 8,
    1254 => 8,
    1255 => 8,
    1256 => 8,
    1257 => 8,
    1258 => 8,
    1259 => 8,
    1260 => 8,
    1261 => 8,
    1262 => 8,
    1263 => 8,
    1264 => 8,
    1265 => 8,
    1266 => 8,
    1267 => 8,
    1268 => 8,
    1269 => 8,
    1270 => 8,
    1271 => 8,
    1272 => 8,
    1273 => 8,
    1274 => 8,
    1275 => 8,
    1276 => 8,
    1277 => 8,
    1278 => 8,
    1279 => 8,
    1280 => 8,
    1281 => 8,
    1282 => 8,
    1283 => 8,
    1284 => 8,
    1285 => 8,
    1286 => 8,
    1287 => 8,
    1288 => 8,
    1289 => 8,
    1290 => 8,
    1291 => 8,
    1292 => 8,
    1293 => 8,
    1294 => 8,
    1295 => 8,
    1296 => 8,
    1297 => 8,
    1298 => 8,
    1299 => 8,
    1300 => 8,
    1301 => 8,
    1302 => 8,
    1303 => 8,
    1304 => 8,
    1305 => 8,
    1306 => 8,
    1307 => 8,
    1308 => 8,
    1309 => 8,
    1310 => 8,
    1311 => 8,
    1312 => 8,
    1313 => 8,
    1314 => 8,
    1315 => 8,
    1316 => 8,
    1317 => 8,
    1318 => 8,
    1319 => 8,
    1320 => 8,
    1321 => 8,
    1322 => 8,
    1323 => 8,
    1324 => 8,
    1325 => 8,
    1326 => 8,
    1327 => 8,
    1328 => 8,
    1329 => 8,
    1330 => 8,
    1331 => 8,
    1332 => 8,
    1333 => 8,
    1334 => 8,
    1335 => 8,
    1336 => 8,
    1337 => 8,
    1338 => 8,
    1339 => 8,
    1340 => 8,
    1341 => 8,
    1342 => 8,
    1343 => 8,
    1344 => 8,
    1345 => 8,
    1346 => 8,
    1347 => 8,
    1348 => 8,
    1349 => 8,
    1350 => 8,
    1351 => 8,
    1352 => 8,
    1353 => 8,
    1354 => 8,
    1355 => 8,
    1356 => 8,
    1357 => 8,
    1358 => 8,
    1359 => 8,
    1360 => 8,
    1361 => 8,
    1362 => 8,
    1363 => 8,
    1364 => 8,
    1365 => 8,
    1366 => 8,
    1367 => 8,
    1368 => 8,
    1369 => 8,
    1370 => 8,
    1371 => 8,
    1372 => 8,
    1373 => 8,
    1374 => 8,
    1375 => 8,
    1376 => 8,
    1377 => 8,
    1378 => 8,
    1379 => 8,
    1380 => 8,
    1381 => 8,
    1382 => 8,
    1383 => 8,
    1384 => 8,
    1385 => 8,
    1386 => 8,
    1387 => 8,
    1388 => 8,
    1389 => 8,
    1390 => 8,
    1391 => 8,
    1392 => 8,
    1393 => 8,
    1394 => 8,
    1395 => 8,
    1396 => 8,
    1397 => 8,
    1398 => 8,
    1399 => 8,
    1400 => 8,
    1401 => 8,
    1402 => 8,
    1403 => 8,
    1404 => 8,
    1405 => 8,
    1406 => 8,
    1407 => 8,
    1408 => 8,
    1409 => 8,
    1410 => 8,
    1411 => 8,
    1412 => 9,
    1413 => 9,
    1414 => 9,
    1415 => 9,
    1416 => 9,
    1417 => 9,
    1418 => 9,
    1419 => 9,
    1420 => 9,
    1421 => 9,
    1422 => 9,
    1423 => 9,
    1424 => 9,
    1425 => 9,
    1426 => 9,
    1427 => 9,
    1428 => 9,
    1429 => 9,
    1430 => 9,
    1431 => 9,
    1432 => 9,
    1433 => 9,
    1434 => 9,
    1435 => 9,
    1436 => 9,
    1437 => 9,
    1438 => 9,
    1439 => 9,
    1440 => 9,
    1441 => 9,
    1442 => 9,
    1443 => 9,
    1444 => 9,
    1445 => 9,
    1446 => 9,
    1447 => 9,
    1448 => 9,
    1449 => 9,
    1450 => 9,
    1451 => 9,
    1452 => 9,
    1453 => 9,
    1454 => 9,
    1455 => 9,
    1456 => 9,
    1457 => 9,
    1458 => 9,
    1459 => 9,
    1460 => 9,
    1461 => 9,
    1462 => 9,
    1463 => 9,
    1464 => 9,
    1465 => 9,
    1466 => 9,
    1467 => 9,
    1468 => 9,
    1469 => 9,
    1470 => 9,
    1471 => 9,
    1472 => 9,
    1473 => 9,
    1474 => 9,
    1475 => 9,
    1476 => 9,
    1477 => 9,
    1478 => 9,
    1479 => 9,
    1480 => 9,
    1481 => 9,
    1482 => 9,
    1483 => 9,
    1484 => 9,
    1485 => 9,
    1486 => 9,
    1487 => 9,
    1488 => 9,
    1489 => 9,
    1490 => 9,
    1491 => 9,
    1492 => 9,
    1493 => 9,
    1494 => 9,
    1495 => 9,
    1496 => 9,
    1497 => 9,
    1498 => 9,
    1499 => 9,
    1500 => 9,
    1501 => 9,
    1502 => 9,
    1503 => 9,
    1504 => 9,
    1505 => 9,
    1506 => 9,
    1507 => 9,
    1508 => 9,
    1509 => 9,
    1510 => 9,
    1511 => 9,
    1512 => 9,
    1513 => 9,
    1514 => 9,
    1515 => 9,
    1516 => 9,
    1517 => 9,
    1518 => 9,
    1519 => 9,
    1520 => 9,
    1521 => 9,
    1522 => 9,
    1523 => 9,
    1524 => 9,
    1525 => 9,
    1526 => 9,
    1527 => 9,
    1528 => 9,
    1529 => 9,
    1530 => 9,
    1531 => 9,
    1532 => 9,
    1533 => 9,
    1534 => 9,
    1535 => 9,
    1536 => 9,
    1537 => 9,
    1538 => 9,
    1539 => 9,
    1540 => 9,
    1541 => 9,
    1542 => 9,
    1543 => 9,
    1544 => 9,
    1545 => 9,
    1546 => 9,
    1547 => 9,
    1548 => 9,
    1549 => 9,
    1550 => 9,
    1551 => 9,
    1552 => 9,
    1553 => 9,
    1554 => 9,
    1555 => 9,
    1556 => 9,
    1557 => 9,
    1558 => 9,
    1559 => 9,
    1560 => 9,
    1561 => 9,
    1562 => 9,
    1563 => 9,
    1564 => 9,
    1565 => 9,
    1566 => 9,
    1567 => 9,
    1568 => 9,
    1569 => 9,
    1570 => 9,
    1571 => 9,
    1572 => 9,
    1573 => 9,
    1574 => 9,
    1575 => 9,
    1576 => 9,
    1577 => 9,
    1578 => 9,
    1579 => 10,
    1580 => 10,
    1581 => 10,
    1582 => 10,
    1583 => 10,
    1584 => 10,
    1585 => 10,
    1586 => 10,
    1587 => 10,
    1588 => 10,
    1589 => 10,
    1590 => 10,
    1591 => 10,
    1592 => 10,
    1593 => 10,
    1594 => 10,
    1595 => 10,
    1596 => 10,
    1597 => 10,
    1598 => 10,
    1599 => 10,
    1600 => 10,
    1601 => 10,
    1602 => 10,
    1603 => 10,
    1604 => 10,
    1605 => 10,
    1606 => 10,
    1607 => 10,
    1608 => 10,
    1609 => 10,
    1610 => 10,
    1611 => 10,
    1612 => 10,
    1613 => 10,
    1614 => 10,
    1615 => 10,
    1616 => 10,
    1617 => 10,
    1618 => 10,
    1619 => 10,
    1620 => 10,
    1621 => 10,
    1622 => 10,
    1623 => 10,
    1624 => 10,
    1625 => 10,
    1626 => 10,
    1627 => 10,
    1628 => 10,
    1629 => 10,
    1630 => 10,
    1631 => 10,
    1632 => 10,
    1633 => 10,
    1634 => 10,
    1635 => 10,
    1636 => 10,
    1637 => 10,
    1638 => 10,
    1639 => 10,
    1640 => 10,
    1641 => 10,
    1642 => 10,
    1643 => 10,
    1644 => 10,
    1645 => 10,
    1646 => 10,
    1647 => 10,
    1648 => 10,
    1649 => 10,
    1650 => 10,
    1651 => 10,
    1652 => 10,
    1653 => 10,
    1654 => 10,
    1655 => 10,
    1656 => 10,
    1657 => 10,
    1658 => 10,
    1659 => 10,
    1660 => 10,
    1661 => 10,
    1662 => 10,
    1663 => 10,
    1664 => 10,
    1665 => 10,
    1666 => 10,
    1667 => 10,
    1668 => 10,
    1669 => 10,
    1670 => 10,
    1671 => 10,
    1672 => 10,
    1673 => 10,
    1674 => 10,
    1675 => 10,
    1676 => 10,
    1677 => 10,
    1678 => 10,
    1679 => 10,
    1680 => 10,
    1681 => 10,
    1682 => 10,
    1683 => 10,
    1684 => 10,
    1685 => 10,
    1686 => 10,
    1687 => 10,
    1688 => 10,
    1689 => 10,
    1690 => 10,
    1691 => 10,
    1692 => 10,
    1693 => 10,
    1694 => 10,
    1695 => 10,
    1696 => 10,
    1697 => 10,
    1698 => 10,
    1699 => 10,
    1700 => 10,
    1701 => 10,
    1702 => 10,
    1703 => 10,
    1704 => 10,
    1705 => 10,
    1706 => 10,
    1707 => 10,
    1708 => 10,
    1709 => 10,
    1710 => 10,
    1711 => 10,
    1712 => 10,
    1713 => 10,
    1714 => 10,
    1715 => 10,
    1716 => 10,
    1717 => 10,
    1718 => 10,
    1719 => 10,
    1720 => 10,
    1721 => 10,
    1722 => 10,
    1723 => 10,
    1724 => 10,
    1725 => 10,
    1726 => 10,
    1727 => 10,
    1728 => 10,
    1729 => 10,
    1730 => 10,
    1731 => 10,
    1732 => 10,
    1733 => 10,
    1734 => 10,
    1735 => 10,
    1736 => 10,
    1737 => 10,
    1738 => 10,
    1739 => 10,
    1740 => 10,
    1741 => 10,
    1742 => 10,
    1743 => 10,
    1744 => 10,
    1745 => 10,
    1746 => 10,
    1747 => 11,
    1748 => 11,
    1749 => 11,
    1750 => 11,
    1751 => 11,
    1752 => 11,
    1753 => 11,
    1754 => 11,
    1755 => 11,
    1756 => 11,
    1757 => 11,
    1758 => 11,
    1759 => 11,
    1760 => 11,
    1761 => 11,
    1762 => 11,
    1763 => 11,
    1764 => 11,
    1765 => 11,
    1766 => 11,
    1767 => 11,
    1768 => 11,
    1769 => 11,
    1770 => 11,
    1771 => 11,
    1772 => 11,
    1773 => 11,
    1774 => 11,
    1775 => 11,
    1776 => 11,
    1777 => 11,
    1778 => 11,
    1779 => 11,
    1780 => 11,
    1781 => 11,
    1782 => 11,
    1783 => 11,
    1784 => 11,
    1785 => 11,
    1786 => 11,
    1787 => 11,
    1788 => 11,
    1789 => 11,
    1790 => 11,
    1791 => 11,
    1792 => 11,
    1793 => 11,
    1794 => 11,
    1795 => 11,
    1796 => 11,
    1797 => 11,
    1798 => 11,
    1799 => 11,
    1800 => 11,
    1801 => 11,
    1802 => 11,
    1803 => 11,
    1804 => 11,
    1805 => 11,
    1806 => 11,
    1807 => 11,
    1808 => 11,
    1809 => 11,
    1810 => 11,
    1811 => 11,
    1812 => 11,
    1813 => 11,
    1814 => 11,
    1815 => 11,
    1816 => 11,
    1817 => 11,
    1818 => 11,
    1819 => 11,
    1820 => 11,
    1821 => 11,
    1822 => 11,
    1823 => 11,
    1824 => 11,
    1825 => 11,
    1826 => 11,
    1827 => 11,
    1828 => 11,
    1829 => 11,
    1830 => 11,
    1831 => 11,
    1832 => 11,
    1833 => 11,
    1834 => 11,
    1835 => 11,
    1836 => 11,
    1837 => 11,
    1838 => 11,
    1839 => 11,
    1840 => 11,
    1841 => 11,
    1842 => 11,
    1843 => 11,
    1844 => 11,
    1845 => 11,
    1846 => 11,
    1847 => 11,
    1848 => 11,
    1849 => 11,
    1850 => 11,
    1851 => 11,
    1852 => 11,
    1853 => 11,
    1854 => 11,
    1855 => 11,
    1856 => 11,
    1857 => 11,
    1858 => 11,
    1859 => 11,
    1860 => 11,
    1861 => 11,
    1862 => 11,
    1863 => 11,
    1864 => 11,
    1865 => 11,
    1866 => 11,
    1867 => 11,
    1868 => 11,
    1869 => 11,
    1870 => 11,
    1871 => 11,
    1872 => 11,
    1873 => 11,
    1874 => 11,
    1875 => 11,
    1876 => 11,
    1877 => 11,
    1878 => 11,
    1879 => 11,
    1880 => 11,
    1881 => 11,
    1882 => 11,
    1883 => 11,
    1884 => 11,
    1885 => 11,
    1886 => 11,
    1887 => 11,
    1888 => 11,
    1889 => 11,
    1890 => 11,
    1891 => 11,
    1892 => 11,
    1893 => 11,
    1894 => 11,
    1895 => 11,
    1896 => 11,
    1897 => 11,
    1898 => 11,
    1899 => 11,
    1900 => 11,
    1901 => 11,
    1902 => 11,
    1903 => 11,
    1904 => 11,
    1905 => 11,
    1906 => 11,
    1907 => 11,
    1908 => 11,
    1909 => 11,
    1910 => 11,
    1911 => 11,
    1912 => 11,
    1913 => 11,
    1914 => 11,
    1915 => 12,
    1916 => 12,
    1917 => 12,
    1918 => 12,
    1919 => 12,
    1920 => 12,
    1921 => 12,
    1922 => 12,
    1923 => 12,
    1924 => 12,
    1925 => 12,
    1926 => 12,
    1927 => 12,
    1928 => 12,
    1929 => 12,
    1930 => 12,
    1931 => 12,
    1932 => 12,
    1933 => 12,
    1934 => 12,
    1935 => 12,
    1936 => 12,
    1937 => 12,
    1938 => 12,
    1939 => 12,
    1940 => 12,
    1941 => 12,
    1942 => 12,
    1943 => 12,
    1944 => 12,
    1945 => 12,
    1946 => 12,
    1947 => 12,
    1948 => 12,
    1949 => 12,
    1950 => 12,
    1951 => 12,
    1952 => 12,
    1953 => 12,
    1954 => 12,
    1955 => 12,
    1956 => 12,
    1957 => 12,
    1958 => 12,
    1959 => 12,
    1960 => 12,
    1961 => 12,
    1962 => 12,
    1963 => 12,
    1964 => 12,
    1965 => 12,
    1966 => 12,
    1967 => 12,
    1968 => 12,
    1969 => 12,
    1970 => 12,
    1971 => 12,
    1972 => 12,
    1973 => 12,
    1974 => 12,
    1975 => 12,
    1976 => 12,
    1977 => 12,
    1978 => 12,
    1979 => 12,
    1980 => 12,
    1981 => 12,
    1982 => 12,
    1983 => 12,
    1984 => 12,
    1985 => 12,
    1986 => 12,
    1987 => 12,
    1988 => 12,
    1989 => 12,
    1990 => 12,
    1991 => 12,
    1992 => 12,
    1993 => 12,
    1994 => 12,
    1995 => 12,
    1996 => 12,
    1997 => 12,
    1998 => 12,
    1999 => 12,
    2000 => 12,
    2001 => 12,
    2002 => 12,
    2003 => 12,
    2004 => 12,
    2005 => 12,
    2006 => 12,
    2007 => 12,
    2008 => 12,
    2009 => 12,
    2010 => 12,
    2011 => 12,
    2012 => 12,
    2013 => 12,
    2014 => 12,
    2015 => 12,
    2016 => 12,
    2017 => 12,
    2018 => 12,
    2019 => 12,
    2020 => 12,
    2021 => 12,
    2022 => 12,
    2023 => 12,
    2024 => 12,
    2025 => 12,
    2026 => 12,
    2027 => 12,
    2028 => 12,
    2029 => 12,
    2030 => 12,
    2031 => 12,
    2032 => 12,
    2033 => 12,
    2034 => 12,
    2035 => 12,
    2036 => 12,
    2037 => 12,
    2038 => 12,
    2039 => 12,
    2040 => 12,
    2041 => 12,
    2042 => 12,
    2043 => 12,
    2044 => 12,
    2045 => 12,
    2046 => 12,
    2047 => 12,
    2048 => 12,
    2049 => 12,
    2050 => 12,
    2051 => 12,
    2052 => 12,
    2053 => 12,
    2054 => 12,
    2055 => 12,
    2056 => 12,
    2057 => 12,
    2058 => 12,
    2059 => 12,
    2060 => 12,
    2061 => 12,
    2062 => 12,
    2063 => 12,
    2064 => 12,
    2065 => 12,
    2066 => 12,
    2067 => 12,
    2068 => 12,
    2069 => 12,
    2070 => 12,
    2071 => 12,
    2072 => 12,
    2073 => 12,
    2074 => 12,
    2075 => 12,
    2076 => 12,
    2077 => 12,
    2078 => 12,
    2079 => 12,
    2080 => 12,
    2081 => 12,
    2082 => 12,
    2083 => 12,
    2084 => 13,
    2085 => 13,
    2086 => 13,
    2087 => 13,
    2088 => 13,
    2089 => 13,
    2090 => 13,
    2091 => 13,
    2092 => 13,
    2093 => 13,
    2094 => 13,
    2095 => 13,
    2096 => 13,
    2097 => 13,
    2098 => 13,
    2099 => 13,
    2100 => 13,
    2101 => 13,
    2102 => 13,
    2103 => 13,
    2104 => 13,
    2105 => 13,
    2106 => 13,
    2107 => 13,
    2108 => 13,
    2109 => 13,
    2110 => 13,
    2111 => 13,
    2112 => 13,
    2113 => 13,
    2114 => 13,
    2115 => 13,
    2116 => 13,
    2117 => 13,
    2118 => 13,
    2119 => 13,
    2120 => 13,
    2121 => 13,
    2122 => 13,
    2123 => 13,
    2124 => 13,
    2125 => 13,
    2126 => 13,
    2127 => 13,
    2128 => 13,
    2129 => 13,
    2130 => 13,
    2131 => 13,
    2132 => 13,
    2133 => 13,
    2134 => 13,
    2135 => 13,
    2136 => 13,
    2137 => 13,
    2138 => 13,
    2139 => 13,
    2140 => 13,
    2141 => 13,
    2142 => 13,
    2143 => 13,
    2144 => 13,
    2145 => 13,
    2146 => 13,
    2147 => 13,
    2148 => 13,
    2149 => 13,
    2150 => 13,
    2151 => 13,
    2152 => 13,
    2153 => 13,
    2154 => 13,
    2155 => 13,
    2156 => 13,
    2157 => 13,
    2158 => 13,
    2159 => 13,
    2160 => 13,
    2161 => 13,
    2162 => 13,
    2163 => 13,
    2164 => 13,
    2165 => 13,
    2166 => 13,
    2167 => 13,
    2168 => 13,
    2169 => 13,
    2170 => 13,
    2171 => 13,
    2172 => 13,
    2173 => 13,
    2174 => 13,
    2175 => 13,
    2176 => 13,
    2177 => 13,
    2178 => 13,
    2179 => 13,
    2180 => 13,
    2181 => 13,
    2182 => 13,
    2183 => 13,
    2184 => 13,
    2185 => 13,
    2186 => 13,
    2187 => 13,
    2188 => 13,
    2189 => 13,
    2190 => 13,
    2191 => 13,
    2192 => 13,
    2193 => 13,
    2194 => 13,
    2195 => 13,
    2196 => 13,
    2197 => 13,
    2198 => 13,
    2199 => 13,
    2200 => 13,
    2201 => 13,
    2202 => 13,
    2203 => 13,
    2204 => 13,
    2205 => 13,
    2206 => 13,
    2207 => 13,
    2208 => 13,
    2209 => 13,
    2210 => 13,
    2211 => 13,
    2212 => 13,
    2213 => 13,
    2214 => 13,
    2215 => 13,
    2216 => 13,
    2217 => 13,
    2218 => 13,
    2219 => 13,
    2220 => 13,
    2221 => 13,
    2222 => 13,
    2223 => 13,
    2224 => 13,
    2225 => 13,
    2226 => 13,
    2227 => 13,
    2228 => 13,
    2229 => 13,
    2230 => 13,
    2231 => 13,
    2232 => 13,
    2233 => 13,
    2234 => 13,
    2235 => 13,
    2236 => 13,
    2237 => 13,
    2238 => 13,
    2239 => 13,
    2240 => 13,
    2241 => 13,
    2242 => 13,
    2243 => 13,
    2244 => 13,
    2245 => 13,
    2246 => 13,
    2247 => 13,
    2248 => 13,
    2249 => 13,
    2250 => 13,
    2251 => 13,
    2252 => 13,
    2253 => 14,
    2254 => 14,
    2255 => 14,
    2256 => 14,
    2257 => 14,
    2258 => 14,
    2259 => 14,
    2260 => 14,
    2261 => 14,
    2262 => 14,
    2263 => 14,
    2264 => 14,
    2265 => 14,
    2266 => 14,
    2267 => 14,
    2268 => 14,
    2269 => 14,
    2270 => 14,
    2271 => 14,
    2272 => 14,
    2273 => 14,
    2274 => 14,
    2275 => 14,
    2276 => 14,
    2277 => 14,
    2278 => 14,
    2279 => 14,
    2280 => 14,
    2281 => 14,
    2282 => 14,
    2283 => 14,
    2284 => 14,
    2285 => 14,
    2286 => 14,
    2287 => 14,
    2288 => 14,
    2289 => 14,
    2290 => 14,
    2291 => 14,
    2292 => 14,
    2293 => 14,
    2294 => 14,
    2295 => 14,
    2296 => 14,
    2297 => 14,
    2298 => 14,
    2299 => 14,
    2300 => 14,
    2301 => 14,
    2302 => 14,
    2303 => 14,
    2304 => 14,
    2305 => 14,
    2306 => 14,
    2307 => 14,
    2308 => 14,
    2309 => 14,
    2310 => 14,
    2311 => 14,
    2312 => 14,
    2313 => 14,
    2314 => 14,
    2315 => 14,
    2316 => 14,
    2317 => 14,
    2318 => 14,
    2319 => 14,
    2320 => 14,
    2321 => 14,
    2322 => 14,
    2323 => 14,
    2324 => 14,
    2325 => 14,
    2326 => 14,
    2327 => 14,
    2328 => 14,
    2329 => 14,
    2330 => 14,
    2331 => 14,
    2332 => 14,
    2333 => 14,
    2334 => 14,
    2335 => 14,
    2336 => 14,
    2337 => 14,
    2338 => 14,
    2339 => 14,
    2340 => 14,
    2341 => 14,
    2342 => 14,
    2343 => 14,
    2344 => 14,
    2345 => 14,
    2346 => 14,
    2347 => 14,
    2348 => 14,
    2349 => 14,
    2350 => 14,
    2351 => 14,
    2352 => 14,
    2353 => 14,
    2354 => 14,
    2355 => 14,
    2356 => 14,
    2357 => 14,
    2358 => 14,
    2359 => 14,
    2360 => 14,
    2361 => 14,
    2362 => 14,
    2363 => 14,
    2364 => 14,
    2365 => 14,
    2366 => 14,
    2367 => 14,
    2368 => 14,
    2369 => 14,
    2370 => 14,
    2371 => 14,
    2372 => 14,
    2373 => 14,
    2374 => 14,
    2375 => 14,
    2376 => 14,
    2377 => 14,
    2378 => 14,
    2379 => 14,
    2380 => 14,
    2381 => 14,
    2382 => 14,
    2383 => 14,
    2384 => 14,
    2385 => 14,
    2386 => 14,
    2387 => 14,
    2388 => 14,
    2389 => 14,
    2390 => 14,
    2391 => 14,
    2392 => 14,
    2393 => 14,
    2394 => 14,
    2395 => 14,
    2396 => 14,
    2397 => 14,
    2398 => 14,
    2399 => 14,
    2400 => 14,
    2401 => 14,
    2402 => 14,
    2403 => 14,
    2404 => 14,
    2405 => 14,
    2406 => 14,
    2407 => 14,
    2408 => 14,
    2409 => 14,
    2410 => 14,
    2411 => 14,
    2412 => 14,
    2413 => 14,
    2414 => 14,
    2415 => 14,
    2416 => 14,
    2417 => 14,
    2418 => 14,
    2419 => 14,
    2420 => 14,
    2421 => 14,
    2422 => 14,
    2423 => 15,
    2424 => 15,
    2425 => 15,
    2426 => 15,
    2427 => 15,
    2428 => 15,
    2429 => 15,
    2430 => 15,
    2431 => 15,
    2432 => 15,
    2433 => 15,
    2434 => 15,
    2435 => 15,
    2436 => 15,
    2437 => 15,
    2438 => 15,
    2439 => 15,
    2440 => 15,
    2441 => 15,
    2442 => 15,
    2443 => 15,
    2444 => 15,
    2445 => 15,
    2446 => 15,
    2447 => 15,
    2448 => 15,
    2449 => 15,
    2450 => 15,
    2451 => 15,
    2452 => 15,
    2453 => 15,
    2454 => 15,
    2455 => 15,
    2456 => 15,
    2457 => 15,
    2458 => 15,
    2459 => 15,
    2460 => 15,
    2461 => 15,
    2462 => 15,
    2463 => 15,
    2464 => 15,
    2465 => 15,
    2466 => 15,
    2467 => 15,
    2468 => 15,
    2469 => 15,
    2470 => 15,
    2471 => 15,
    2472 => 15,
    2473 => 15,
    2474 => 15,
    2475 => 15,
    2476 => 15,
    2477 => 15,
    2478 => 15,
    2479 => 15,
    2480 => 15,
    2481 => 15,
    2482 => 15,
    2483 => 15,
    2484 => 15,
    2485 => 15,
    2486 => 15,
    2487 => 15,
    2488 => 15,
    2489 => 15,
    2490 => 15,
    2491 => 15,
    2492 => 15,
    2493 => 15,
    2494 => 15,
    2495 => 15,
    2496 => 15,
    2497 => 15,
    2498 => 15,
    2499 => 15,
    2500 => 15,
    2501 => 15,
    2502 => 15,
    2503 => 15,
    2504 => 15,
    2505 => 15,
    2506 => 15,
    2507 => 15,
    2508 => 15,
    2509 => 15,
    2510 => 15,
    2511 => 15,
    2512 => 15,
    2513 => 15,
    2514 => 15,
    2515 => 15,
    2516 => 15,
    2517 => 15,
    2518 => 15,
    2519 => 15,
    2520 => 15,
    2521 => 15,
    2522 => 15,
    2523 => 15,
    2524 => 15,
    2525 => 15,
    2526 => 15,
    2527 => 15,
    2528 => 15,
    2529 => 15,
    2530 => 15,
    2531 => 15,
    2532 => 15,
    2533 => 15,
    2534 => 15,
    2535 => 15,
    2536 => 15,
    2537 => 15,
    2538 => 15,
    2539 => 15,
    2540 => 15,
    2541 => 15,
    2542 => 15,
    2543 => 15,
    2544 => 15,
    2545 => 15,
    2546 => 15,
    2547 => 15,
    2548 => 15,
    2549 => 15,
    2550 => 15,
    2551 => 15,
    2552 => 15,
    2553 => 15,
    2554 => 15,
    2555 => 15,
    2556 => 15,
    2557 => 15,
    2558 => 15,
    2559 => 15,
    2560 => 15,
    2561 => 15,
    2562 => 15,
    2563 => 15,
    2564 => 15,
    2565 => 15,
    2566 => 15,
    2567 => 15,
    2568 => 15,
    2569 => 15,
    2570 => 15,
    2571 => 15,
    2572 => 15,
    2573 => 15,
    2574 => 15,
    2575 => 15,
    2576 => 15,
    2577 => 15,
    2578 => 15,
    2579 => 15,
    2580 => 15,
    2581 => 15,
    2582 => 15,
    2583 => 15,
    2584 => 15,
    2585 => 15,
    2586 => 15,
    2587 => 15,
    2588 => 15,
    2589 => 15,
    2590 => 15,
    2591 => 15,
    2592 => 15,
    2593 => 16,
    2594 => 16,
    2595 => 16,
    2596 => 16,
    2597 => 16,
    2598 => 16,
    2599 => 16,
    2600 => 16,
    2601 => 16,
    2602 => 16,
    2603 => 16,
    2604 => 16,
    2605 => 16,
    2606 => 16,
    2607 => 16,
    2608 => 16,
    2609 => 16,
    2610 => 16,
    2611 => 16,
    2612 => 16,
    2613 => 16,
    2614 => 16,
    2615 => 16,
    2616 => 16,
    2617 => 16,
    2618 => 16,
    2619 => 16,
    2620 => 16,
    2621 => 16,
    2622 => 16,
    2623 => 16,
    2624 => 16,
    2625 => 16,
    2626 => 16,
    2627 => 16,
    2628 => 16,
    2629 => 16,
    2630 => 16,
    2631 => 16,
    2632 => 16,
    2633 => 16,
    2634 => 16,
    2635 => 16,
    2636 => 16,
    2637 => 16,
    2638 => 16,
    2639 => 16,
    2640 => 16,
    2641 => 16,
    2642 => 16,
    2643 => 16,
    2644 => 16,
    2645 => 16,
    2646 => 16,
    2647 => 16,
    2648 => 16,
    2649 => 16,
    2650 => 16,
    2651 => 16,
    2652 => 16,
    2653 => 16,
    2654 => 16,
    2655 => 16,
    2656 => 16,
    2657 => 16,
    2658 => 16,
    2659 => 16,
    2660 => 16,
    2661 => 16,
    2662 => 16,
    2663 => 16,
    2664 => 16,
    2665 => 16,
    2666 => 16,
    2667 => 16,
    2668 => 16,
    2669 => 16,
    2670 => 16,
    2671 => 16,
    2672 => 16,
    2673 => 16,
    2674 => 16,
    2675 => 16,
    2676 => 16,
    2677 => 16,
    2678 => 16,
    2679 => 16,
    2680 => 16,
    2681 => 16,
    2682 => 16,
    2683 => 16,
    2684 => 16,
    2685 => 16,
    2686 => 16,
    2687 => 16,
    2688 => 16,
    2689 => 16,
    2690 => 16,
    2691 => 16,
    2692 => 16,
    2693 => 16,
    2694 => 16,
    2695 => 16,
    2696 => 16,
    2697 => 16,
    2698 => 16,
    2699 => 16,
    2700 => 16,
    2701 => 16,
    2702 => 16,
    2703 => 16,
    2704 => 16,
    2705 => 16,
    2706 => 16,
    2707 => 16,
    2708 => 16,
    2709 => 16,
    2710 => 16,
    2711 => 16,
    2712 => 16,
    2713 => 16,
    2714 => 16,
    2715 => 16,
    2716 => 16,
    2717 => 16,
    2718 => 16,
    2719 => 16,
    2720 => 16,
    2721 => 16,
    2722 => 16,
    2723 => 16,
    2724 => 16,
    2725 => 16,
    2726 => 16,
    2727 => 16,
    2728 => 16,
    2729 => 16,
    2730 => 16,
    2731 => 16,
    2732 => 16,
    2733 => 16,
    2734 => 16,
    2735 => 16,
    2736 => 16,
    2737 => 16,
    2738 => 16,
    2739 => 16,
    2740 => 16,
    2741 => 16,
    2742 => 16,
    2743 => 16,
    2744 => 16,
    2745 => 16,
    2746 => 16,
    2747 => 16,
    2748 => 16,
    2749 => 16,
    2750 => 16,
    2751 => 16,
    2752 => 16,
    2753 => 16,
    2754 => 16,
    2755 => 16,
    2756 => 16,
    2757 => 16,
    2758 => 16,
    2759 => 16,
    2760 => 16,
    2761 => 16,
    2762 => 16,
    2763 => 16,
    2764 => 16,
    2765 => 17,
    2766 => 17,
    2767 => 17,
    2768 => 17,
    2769 => 17,
    2770 => 17,
    2771 => 17,
    2772 => 17,
    2773 => 17,
    2774 => 17,
    2775 => 17,
    2776 => 17,
    2777 => 17,
    2778 => 17,
    2779 => 17,
    2780 => 17,
    2781 => 17,
    2782 => 17,
    2783 => 17,
    2784 => 17,
    2785 => 17,
    2786 => 17,
    2787 => 17,
    2788 => 17,
    2789 => 17,
    2790 => 17,
    2791 => 17,
    2792 => 17,
    2793 => 17,
    2794 => 17,
    2795 => 17,
    2796 => 17,
    2797 => 17,
    2798 => 17,
    2799 => 17,
    2800 => 17,
    2801 => 17,
    2802 => 17,
    2803 => 17,
    2804 => 17,
    2805 => 17,
    2806 => 17,
    2807 => 17,
    2808 => 17,
    2809 => 17,
    2810 => 17,
    2811 => 17,
    2812 => 17,
    2813 => 17,
    2814 => 17,
    2815 => 17,
    2816 => 17,
    2817 => 17,
    2818 => 17,
    2819 => 17,
    2820 => 17,
    2821 => 17,
    2822 => 17,
    2823 => 17,
    2824 => 17,
    2825 => 17,
    2826 => 17,
    2827 => 17,
    2828 => 17,
    2829 => 17,
    2830 => 17,
    2831 => 17,
    2832 => 17,
    2833 => 17,
    2834 => 17,
    2835 => 17,
    2836 => 17,
    2837 => 17,
    2838 => 17,
    2839 => 17,
    2840 => 17,
    2841 => 17,
    2842 => 17,
    2843 => 17,
    2844 => 17,
    2845 => 17,
    2846 => 17,
    2847 => 17,
    2848 => 17,
    2849 => 17,
    2850 => 17,
    2851 => 17,
    2852 => 17,
    2853 => 17,
    2854 => 17,
    2855 => 17,
    2856 => 17,
    2857 => 17,
    2858 => 17,
    2859 => 17,
    2860 => 17,
    2861 => 17,
    2862 => 17,
    2863 => 17,
    2864 => 17,
    2865 => 17,
    2866 => 17,
    2867 => 17,
    2868 => 17,
    2869 => 17,
    2870 => 17,
    2871 => 17,
    2872 => 17,
    2873 => 17,
    2874 => 17,
    2875 => 17,
    2876 => 17,
    2877 => 17,
    2878 => 17,
    2879 => 17,
    2880 => 17,
    2881 => 17,
    2882 => 17,
    2883 => 17,
    2884 => 17,
    2885 => 17,
    2886 => 17,
    2887 => 17,
    2888 => 17,
    2889 => 17,
    2890 => 17,
    2891 => 17,
    2892 => 17,
    2893 => 17,
    2894 => 17,
    2895 => 17,
    2896 => 17,
    2897 => 17,
    2898 => 17,
    2899 => 17,
    2900 => 17,
    2901 => 17,
    2902 => 17,
    2903 => 17,
    2904 => 17,
    2905 => 17,
    2906 => 17,
    2907 => 17,
    2908 => 17,
    2909 => 17,
    2910 => 17,
    2911 => 17,
    2912 => 17,
    2913 => 17,
    2914 => 17,
    2915 => 17,
    2916 => 17,
    2917 => 17,
    2918 => 17,
    2919 => 17,
    2920 => 17,
    2921 => 17,
    2922 => 17,
    2923 => 17,
    2924 => 17,
    2925 => 17,
    2926 => 17,
    2927 => 17,
    2928 => 17,
    2929 => 17,
    2930 => 17,
    2931 => 17,
    2932 => 17,
    2933 => 17,
    2934 => 17,
    2935 => 17,
    2936 => 18,
    2937 => 18,
    2938 => 18,
    2939 => 18,
    2940 => 18,
    2941 => 18,
    2942 => 18,
    2943 => 18,
    2944 => 18,
    2945 => 18,
    2946 => 18,
    2947 => 18,
    2948 => 18,
    2949 => 18,
    2950 => 18,
    2951 => 18,
    2952 => 18,
    2953 => 18,
    2954 => 18,
    2955 => 18,
    2956 => 18,
    2957 => 18,
    2958 => 18,
    2959 => 18,
    2960 => 18,
    2961 => 18,
    2962 => 18,
    2963 => 18,
    2964 => 18,
    2965 => 18,
    2966 => 18,
    2967 => 18,
    2968 => 18,
    2969 => 18,
    2970 => 18,
    2971 => 18,
    2972 => 18,
    2973 => 18,
    2974 => 18,
    2975 => 18,
    2976 => 18,
    2977 => 18,
    2978 => 18,
    2979 => 18,
    2980 => 18,
    2981 => 18,
    2982 => 18,
    2983 => 18,
    2984 => 18,
    2985 => 18,
    2986 => 18,
    2987 => 18,
    2988 => 18,
    2989 => 18,
    2990 => 18,
    2991 => 18,
    2992 => 18,
    2993 => 18,
    2994 => 18,
    2995 => 18,
    2996 => 18,
    2997 => 18,
    2998 => 18,
    2999 => 18,
    3000 => 18,
    3001 => 18,
    3002 => 18,
    3003 => 18,
    3004 => 18,
    3005 => 18,
    3006 => 18,
    3007 => 18,
    3008 => 18,
    3009 => 18,
    3010 => 18,
    3011 => 18,
    3012 => 18,
    3013 => 18,
    3014 => 18,
    3015 => 18,
    3016 => 18,
    3017 => 18,
    3018 => 18,
    3019 => 18,
    3020 => 18,
    3021 => 18,
    3022 => 18,
    3023 => 18,
    3024 => 18,
    3025 => 18,
    3026 => 18,
    3027 => 18,
    3028 => 18,
    3029 => 18,
    3030 => 18,
    3031 => 18,
    3032 => 18,
    3033 => 18,
    3034 => 18,
    3035 => 18,
    3036 => 18,
    3037 => 18,
    3038 => 18,
    3039 => 18,
    3040 => 18,
    3041 => 18,
    3042 => 18,
    3043 => 18,
    3044 => 18,
    3045 => 18,
    3046 => 18,
    3047 => 18,
    3048 => 18,
    3049 => 18,
    3050 => 18,
    3051 => 18,
    3052 => 18,
    3053 => 18,
    3054 => 18,
    3055 => 18,
    3056 => 18,
    3057 => 18,
    3058 => 18,
    3059 => 18,
    3060 => 18,
    3061 => 18,
    3062 => 18,
    3063 => 18,
    3064 => 18,
    3065 => 18,
    3066 => 18,
    3067 => 18,
    3068 => 18,
    3069 => 18,
    3070 => 18,
    3071 => 18,
    3072 => 18,
    3073 => 18,
    3074 => 18,
    3075 => 18,
    3076 => 18,
    3077 => 18,
    3078 => 18,
    3079 => 18,
    3080 => 18,
    3081 => 18,
    3082 => 18,
    3083 => 18,
    3084 => 18,
    3085 => 18,
    3086 => 18,
    3087 => 18,
    3088 => 18,
    3089 => 18,
    3090 => 18,
    3091 => 18,
    3092 => 18,
    3093 => 18,
    3094 => 18,
    3095 => 18,
    3096 => 18,
    3097 => 18,
    3098 => 18,
    3099 => 18,
    3100 => 18,
    3101 => 18,
    3102 => 18,
    3103 => 18,
    3104 => 18,
    3105 => 18,
    3106 => 18,
    3107 => 18,
    3108 => 18,
    3109 => 19,
    3110 => 19,
    3111 => 19,
    3112 => 19,
    3113 => 19,
    3114 => 19,
    3115 => 19,
    3116 => 19,
    3117 => 19,
    3118 => 19,
    3119 => 19,
    3120 => 19,
    3121 => 19,
    3122 => 19,
    3123 => 19,
    3124 => 19,
    3125 => 19,
    3126 => 19,
    3127 => 19,
    3128 => 19,
    3129 => 19,
    3130 => 19,
    3131 => 19,
    3132 => 19,
    3133 => 19,
    3134 => 19,
    3135 => 19,
    3136 => 19,
    3137 => 19,
    3138 => 19,
    3139 => 19,
    3140 => 19,
    3141 => 19,
    3142 => 19,
    3143 => 19,
    3144 => 19,
    3145 => 19,
    3146 => 19,
    3147 => 19,
    3148 => 19,
    3149 => 19,
    3150 => 19,
    3151 => 19,
    3152 => 19,
    3153 => 19,
    3154 => 19,
    3155 => 19,
    3156 => 19,
    3157 => 19,
    3158 => 19,
    3159 => 19,
    3160 => 19,
    3161 => 19,
    3162 => 19,
    3163 => 19,
    3164 => 19,
    3165 => 19,
    3166 => 19,
    3167 => 19,
    3168 => 19,
    3169 => 19,
    3170 => 19,
    3171 => 19,
    3172 => 19,
    3173 => 19,
    3174 => 19,
    3175 => 19,
    3176 => 19,
    3177 => 19,
    3178 => 19,
    3179 => 19,
    3180 => 19,
    3181 => 19,
    3182 => 19,
    3183 => 19,
    3184 => 19,
    3185 => 19,
    3186 => 19,
    3187 => 19,
    3188 => 19,
    3189 => 19,
    3190 => 19,
    3191 => 19,
    3192 => 19,
    3193 => 19,
    3194 => 19,
    3195 => 19,
    3196 => 19,
    3197 => 19,
    3198 => 19,
    3199 => 19,
    3200 => 19,
    3201 => 19,
    3202 => 19,
    3203 => 19,
    3204 => 19,
    3205 => 19,
    3206 => 19,
    3207 => 19,
    3208 => 19,
    3209 => 19,
    3210 => 19,
    3211 => 19,
    3212 => 19,
    3213 => 19,
    3214 => 19,
    3215 => 19,
    3216 => 19,
    3217 => 19,
    3218 => 19,
    3219 => 19,
    3220 => 19,
    3221 => 19,
    3222 => 19,
    3223 => 19,
    3224 => 19,
    3225 => 19,
    3226 => 19,
    3227 => 19,
    3228 => 19,
    3229 => 19,
    3230 => 19,
    3231 => 19,
    3232 => 19,
    3233 => 19,
    3234 => 19,
    3235 => 19,
    3236 => 19,
    3237 => 19,
    3238 => 19,
    3239 => 19,
    3240 => 19,
    3241 => 19,
    3242 => 19,
    3243 => 19,
    3244 => 19,
    3245 => 19,
    3246 => 19,
    3247 => 19,
    3248 => 19,
    3249 => 19,
    3250 => 19,
    3251 => 19,
    3252 => 19,
    3253 => 19,
    3254 => 19,
    3255 => 19,
    3256 => 19,
    3257 => 19,
    3258 => 19,
    3259 => 19,
    3260 => 19,
    3261 => 19,
    3262 => 19,
    3263 => 19,
    3264 => 19,
    3265 => 19,
    3266 => 19,
    3267 => 19,
    3268 => 19,
    3269 => 19,
    3270 => 19,
    3271 => 19,
    3272 => 19,
    3273 => 19,
    3274 => 19,
    3275 => 19,
    3276 => 19,
    3277 => 19,
    3278 => 19,
    3279 => 19,
    3280 => 19,
    3281 => 19,
    3282 => 19,
    3283 => 20,
    3284 => 20,
    3285 => 20,
    3286 => 20,
    3287 => 20,
    3288 => 20,
    3289 => 20,
    3290 => 20,
    3291 => 20,
    3292 => 20,
    3293 => 20,
    3294 => 20,
    3295 => 20,
    3296 => 20,
    3297 => 20,
    3298 => 20,
    3299 => 20,
    3300 => 20,
    3301 => 20,
    3302 => 20,
    3303 => 20,
    3304 => 20,
    3305 => 20,
    3306 => 20,
    3307 => 20,
    3308 => 20,
    3309 => 20,
    3310 => 20,
    3311 => 20,
    3312 => 20,
    3313 => 20,
    3314 => 20,
    3315 => 20,
    3316 => 20,
    3317 => 20,
    3318 => 20,
    3319 => 20,
    3320 => 20,
    3321 => 20,
    3322 => 20,
    3323 => 20,
    3324 => 20,
    3325 => 20,
    3326 => 20,
    3327 => 20,
    3328 => 20,
    3329 => 20,
    3330 => 20,
    3331 => 20,
    3332 => 20,
    3333 => 20,
    3334 => 20,
    3335 => 20,
    3336 => 20,
    3337 => 20,
    3338 => 20,
    3339 => 20,
    3340 => 20,
    3341 => 20,
    3342 => 20,
    3343 => 20,
    3344 => 20,
    3345 => 20,
    3346 => 20,
    3347 => 20,
    3348 => 20,
    3349 => 20,
    3350 => 20,
    3351 => 20,
    3352 => 20,
    3353 => 20,
    3354 => 20,
    3355 => 20,
    3356 => 20,
    3357 => 20,
    3358 => 20,
    3359 => 20,
    3360 => 20,
    3361 => 20,
    3362 => 20,
    3363 => 20,
    3364 => 20,
    3365 => 20,
    3366 => 20,
    3367 => 20,
    3368 => 20,
    3369 => 20,
    3370 => 20,
    3371 => 20,
    3372 => 20,
    3373 => 20,
    3374 => 20,
    3375 => 20,
    3376 => 20,
    3377 => 20,
    3378 => 20,
    3379 => 20,
    3380 => 20,
    3381 => 20,
    3382 => 20,
    3383 => 20,
    3384 => 20,
    3385 => 20,
    3386 => 20,
    3387 => 20,
    3388 => 20,
    3389 => 20,
    3390 => 20,
    3391 => 20,
    3392 => 20,
    3393 => 20,
    3394 => 20,
    3395 => 20,
    3396 => 20,
    3397 => 20,
    3398 => 20,
    3399 => 20,
    3400 => 20,
    3401 => 20,
    3402 => 20,
    3403 => 20,
    3404 => 20,
    3405 => 20,
    3406 => 20,
    3407 => 20,
    3408 => 20,
    3409 => 20,
    3410 => 20,
    3411 => 20,
    3412 => 20,
    3413 => 20,
    3414 => 20,
    3415 => 20,
    3416 => 20,
    3417 => 20,
    3418 => 20,
    3419 => 20,
    3420 => 20,
    3421 => 20,
    3422 => 20,
    3423 => 20,
    3424 => 20,
    3425 => 20,
    3426 => 20,
    3427 => 20,
    3428 => 20,
    3429 => 20,
    3430 => 20,
    3431 => 20,
    3432 => 20,
    3433 => 20,
    3434 => 20,
    3435 => 20,
    3436 => 20,
    3437 => 20,
    3438 => 20,
    3439 => 20,
    3440 => 20,
    3441 => 20,
    3442 => 20,
    3443 => 20,
    3444 => 20,
    3445 => 20,
    3446 => 20,
    3447 => 20,
    3448 => 20,
    3449 => 20,
    3450 => 20,
    3451 => 20,
    3452 => 20,
    3453 => 20,
    3454 => 20,
    3455 => 20,
    3456 => 20,
    3457 => 21,
    3458 => 21,
    3459 => 21,
    3460 => 21,
    3461 => 21,
    3462 => 21,
    3463 => 21,
    3464 => 21,
    3465 => 21,
    3466 => 21,
    3467 => 21,
    3468 => 21,
    3469 => 21,
    3470 => 21,
    3471 => 21,
    3472 => 21,
    3473 => 21,
    3474 => 21,
    3475 => 21,
    3476 => 21,
    3477 => 21,
    3478 => 21,
    3479 => 21,
    3480 => 21,
    3481 => 21,
    3482 => 21,
    3483 => 21,
    3484 => 21,
    3485 => 21,
    3486 => 21,
    3487 => 21,
    3488 => 21,
    3489 => 21,
    3490 => 21,
    3491 => 21,
    3492 => 21,
    3493 => 21,
    3494 => 21,
    3495 => 21,
    3496 => 21,
    3497 => 21,
    3498 => 21,
    3499 => 21,
    3500 => 21,
    3501 => 21,
    3502 => 21,
    3503 => 21,
    3504 => 21,
    3505 => 21,
    3506 => 21,
    3507 => 21,
    3508 => 21,
    3509 => 21,
    3510 => 21,
    3511 => 21,
    3512 => 21,
    3513 => 21,
    3514 => 21,
    3515 => 21,
    3516 => 21,
    3517 => 21,
    3518 => 21,
    3519 => 21,
    3520 => 21,
    3521 => 21,
    3522 => 21,
    3523 => 21,
    3524 => 21,
    3525 => 21,
    3526 => 21,
    3527 => 21,
    3528 => 21,
    3529 => 21,
    3530 => 21,
    3531 => 21,
    3532 => 21,
    3533 => 21,
    3534 => 21,
    3535 => 21,
    3536 => 21,
    3537 => 21,
    3538 => 21,
    3539 => 21,
    3540 => 21,
    3541 => 21,
    3542 => 21,
    3543 => 21,
    3544 => 21,
    3545 => 21,
    3546 => 21,
    3547 => 21,
    3548 => 21,
    3549 => 21,
    3550 => 21,
    3551 => 21,
    3552 => 21,
    3553 => 21,
    3554 => 21,
    3555 => 21,
    3556 => 21,
    3557 => 21,
    3558 => 21,
    3559 => 21,
    3560 => 21,
    3561 => 21,
    3562 => 21,
    3563 => 21,
    3564 => 21,
    3565 => 21,
    3566 => 21,
    3567 => 21,
    3568 => 21,
    3569 => 21,
    3570 => 21,
    3571 => 21,
    3572 => 21,
    3573 => 21,
    3574 => 21,
    3575 => 21,
    3576 => 21,
    3577 => 21,
    3578 => 21,
    3579 => 21,
    3580 => 21,
    3581 => 21,
    3582 => 21,
    3583 => 21,
    3584 => 21,
    3585 => 21,
    3586 => 21,
    3587 => 21,
    3588 => 21,
    3589 => 21,
    3590 => 21,
    3591 => 21,
    3592 => 21,
    3593 => 21,
    3594 => 21,
    3595 => 21,
    3596 => 21,
    3597 => 21,
    3598 => 21,
    3599 => 21,
    3600 => 21,
    3601 => 21,
    3602 => 21,
    3603 => 21,
    3604 => 21,
    3605 => 21,
    3606 => 21,
    3607 => 21,
    3608 => 21,
    3609 => 21,
    3610 => 21,
    3611 => 21,
    3612 => 21,
    3613 => 21,
    3614 => 21,
    3615 => 21,
    3616 => 21,
    3617 => 21,
    3618 => 21,
    3619 => 21,
    3620 => 21,
    3621 => 21,
    3622 => 21,
    3623 => 21,
    3624 => 21,
    3625 => 21,
    3626 => 21,
    3627 => 21,
    3628 => 21,
    3629 => 21,
    3630 => 21,
    3631 => 21,
    3632 => 21,
    3633 => 22,
    3634 => 22,
    3635 => 22,
    3636 => 22,
    3637 => 22,
    3638 => 22,
    3639 => 22,
    3640 => 22,
    3641 => 22,
    3642 => 22,
    3643 => 22,
    3644 => 22,
    3645 => 22,
    3646 => 22,
    3647 => 22,
    3648 => 22,
    3649 => 22,
    3650 => 22,
    3651 => 22,
    3652 => 22,
    3653 => 22,
    3654 => 22,
    3655 => 22,
    3656 => 22,
    3657 => 22,
    3658 => 22,
    3659 => 22,
    3660 => 22,
    3661 => 22,
    3662 => 22,
    3663 => 22,
    3664 => 22,
    3665 => 22,
    3666 => 22,
    3667 => 22,
    3668 => 22,
    3669 => 22,
    3670 => 22,
    3671 => 22,
    3672 => 22,
    3673 => 22,
    3674 => 22,
    3675 => 22,
    3676 => 22,
    3677 => 22,
    3678 => 22,
    3679 => 22,
    3680 => 22,
    3681 => 22,
    3682 => 22,
    3683 => 22,
    3684 => 22,
    3685 => 22,
    3686 => 22,
    3687 => 22,
    3688 => 22,
    3689 => 22,
    3690 => 22,
    3691 => 22,
    3692 => 22,
    3693 => 22,
    3694 => 22,
    3695 => 22,
    3696 => 22,
    3697 => 22,
    3698 => 22,
    3699 => 22,
    3700 => 22,
    3701 => 22,
    3702 => 22,
    3703 => 22,
    3704 => 22,
    3705 => 22,
    3706 => 22,
    3707 => 22,
    3708 => 22,
    3709 => 22,
    3710 => 22,
    3711 => 22,
    3712 => 22,
    3713 => 22,
    3714 => 22,
    3715 => 22,
    3716 => 22,
    3717 => 22,
    3718 => 22,
    3719 => 22,
    3720 => 22,
    3721 => 22,
    3722 => 22,
    3723 => 22,
    3724 => 22,
    3725 => 22,
    3726 => 22,
    3727 => 22,
    3728 => 22,
    3729 => 22,
    3730 => 22,
    3731 => 22,
    3732 => 22,
    3733 => 22,
    3734 => 22,
    3735 => 22,
    3736 => 22,
    3737 => 22,
    3738 => 22,
    3739 => 22,
    3740 => 22,
    3741 => 22,
    3742 => 22,
    3743 => 22,
    3744 => 22,
    3745 => 22,
    3746 => 22,
    3747 => 22,
    3748 => 22,
    3749 => 22,
    3750 => 22,
    3751 => 22,
    3752 => 22,
    3753 => 22,
    3754 => 22,
    3755 => 22,
    3756 => 22,
    3757 => 22,
    3758 => 22,
    3759 => 22,
    3760 => 22,
    3761 => 22,
    3762 => 22,
    3763 => 22,
    3764 => 22,
    3765 => 22,
    3766 => 22,
    3767 => 22,
    3768 => 22,
    3769 => 22,
    3770 => 22,
    3771 => 22,
    3772 => 22,
    3773 => 22,
    3774 => 22,
    3775 => 22,
    3776 => 22,
    3777 => 22,
    3778 => 22,
    3779 => 22,
    3780 => 22,
    3781 => 22,
    3782 => 22,
    3783 => 22,
    3784 => 22,
    3785 => 22,
    3786 => 22,
    3787 => 22,
    3788 => 22,
    3789 => 22,
    3790 => 22,
    3791 => 22,
    3792 => 22,
    3793 => 22,
    3794 => 22,
    3795 => 22,
    3796 => 22,
    3797 => 22,
    3798 => 22,
    3799 => 22,
    3800 => 22,
    3801 => 22,
    3802 => 22,
    3803 => 22,
    3804 => 22,
    3805 => 22,
    3806 => 22,
    3807 => 22,
    3808 => 22,
    3809 => 22,
    3810 => 23,
    3811 => 23,
    3812 => 23,
    3813 => 23,
    3814 => 23,
    3815 => 23,
    3816 => 23,
    3817 => 23,
    3818 => 23,
    3819 => 23,
    3820 => 23,
    3821 => 23,
    3822 => 23,
    3823 => 23,
    3824 => 23,
    3825 => 23,
    3826 => 23,
    3827 => 23,
    3828 => 23,
    3829 => 23,
    3830 => 23,
    3831 => 23,
    3832 => 23,
    3833 => 23,
    3834 => 23,
    3835 => 23,
    3836 => 23,
    3837 => 23,
    3838 => 23,
    3839 => 23,
    3840 => 23,
    3841 => 23,
    3842 => 23,
    3843 => 23,
    3844 => 23,
    3845 => 23,
    3846 => 23,
    3847 => 23,
    3848 => 23,
    3849 => 23,
    3850 => 23,
    3851 => 23,
    3852 => 23,
    3853 => 23,
    3854 => 23,
    3855 => 23,
    3856 => 23,
    3857 => 23,
    3858 => 23,
    3859 => 23,
    3860 => 23,
    3861 => 23,
    3862 => 23,
    3863 => 23,
    3864 => 23,
    3865 => 23,
    3866 => 23,
    3867 => 23,
    3868 => 23,
    3869 => 23,
    3870 => 23,
    3871 => 23,
    3872 => 23,
    3873 => 23,
    3874 => 23,
    3875 => 23,
    3876 => 23,
    3877 => 23,
    3878 => 23,
    3879 => 23,
    3880 => 23,
    3881 => 23,
    3882 => 23,
    3883 => 23,
    3884 => 23,
    3885 => 23,
    3886 => 23,
    3887 => 23,
    3888 => 23,
    3889 => 23,
    3890 => 23,
    3891 => 23,
    3892 => 23,
    3893 => 23,
    3894 => 23,
    3895 => 23,
    3896 => 23,
    3897 => 23,
    3898 => 23,
    3899 => 23,
    3900 => 23,
    3901 => 23,
    3902 => 23,
    3903 => 23,
    3904 => 23,
    3905 => 23,
    3906 => 23,
    3907 => 23,
    3908 => 23,
    3909 => 23,
    3910 => 23,
    3911 => 23,
    3912 => 23,
    3913 => 23,
    3914 => 23,
    3915 => 23,
    3916 => 23,
    3917 => 23,
    3918 => 23,
    3919 => 23,
    3920 => 23,
    3921 => 23,
    3922 => 23,
    3923 => 23,
    3924 => 23,
    3925 => 23,
    3926 => 23,
    3927 => 23,
    3928 => 23,
    3929 => 23,
    3930 => 23,
    3931 => 23,
    3932 => 23,
    3933 => 23,
    3934 => 23,
    3935 => 23,
    3936 => 23,
    3937 => 23,
    3938 => 23,
    3939 => 23,
    3940 => 23,
    3941 => 23,
    3942 => 23,
    3943 => 23,
    3944 => 23,
    3945 => 23,
    3946 => 23,
    3947 => 23,
    3948 => 23,
    3949 => 23,
    3950 => 23,
    3951 => 23,
    3952 => 23,
    3953 => 23,
    3954 => 23,
    3955 => 23,
    3956 => 23,
    3957 => 23,
    3958 => 23,
    3959 => 23,
    3960 => 23,
    3961 => 23,
    3962 => 23,
    3963 => 23,
    3964 => 23,
    3965 => 23,
    3966 => 23,
    3967 => 23,
    3968 => 23,
    3969 => 23,
    3970 => 23,
    3971 => 23,
    3972 => 23,
    3973 => 23,
    3974 => 23,
    3975 => 23,
    3976 => 23,
    3977 => 23,
    3978 => 23,
    3979 => 23,
    3980 => 23,
    3981 => 23,
    3982 => 23,
    3983 => 23,
    3984 => 23,
    3985 => 23,
    3986 => 23,
    3987 => 23,
    3988 => 24,
    3989 => 24,
    3990 => 24,
    3991 => 24,
    3992 => 24,
    3993 => 24,
    3994 => 24,
    3995 => 24,
    3996 => 24,
    3997 => 24,
    3998 => 24,
    3999 => 24,
    4000 => 24,
    4001 => 24,
    4002 => 24,
    4003 => 24,
    4004 => 24,
    4005 => 24,
    4006 => 24,
    4007 => 24,
    4008 => 24,
    4009 => 24,
    4010 => 24,
    4011 => 24,
    4012 => 24,
    4013 => 24,
    4014 => 24,
    4015 => 24,
    4016 => 24,
    4017 => 24,
    4018 => 24,
    4019 => 24,
    4020 => 24,
    4021 => 24,
    4022 => 24,
    4023 => 24,
    4024 => 24,
    4025 => 24,
    4026 => 24,
    4027 => 24,
    4028 => 24,
    4029 => 24,
    4030 => 24,
    4031 => 24,
    4032 => 24,
    4033 => 24,
    4034 => 24,
    4035 => 24,
    4036 => 24,
    4037 => 24,
    4038 => 24,
    4039 => 24,
    4040 => 24,
    4041 => 24,
    4042 => 24,
    4043 => 24,
    4044 => 24,
    4045 => 24,
    4046 => 24,
    4047 => 24,
    4048 => 24,
    4049 => 24,
    4050 => 24,
    4051 => 24,
    4052 => 24,
    4053 => 24,
    4054 => 24,
    4055 => 24,
    4056 => 24,
    4057 => 24,
    4058 => 24,
    4059 => 24,
    4060 => 24,
    4061 => 24,
    4062 => 24,
    4063 => 24,
    4064 => 24,
    4065 => 24,
    4066 => 24,
    4067 => 24,
    4068 => 24,
    4069 => 24,
    4070 => 24,
    4071 => 24,
    4072 => 24,
    4073 => 24,
    4074 => 24,
    4075 => 24,
    4076 => 24,
    4077 => 24,
    4078 => 24,
    4079 => 24,
    4080 => 24,
    4081 => 24,
    4082 => 24,
    4083 => 24,
    4084 => 24,
    4085 => 24,
    4086 => 24,
    4087 => 24,
    4088 => 24,
    4089 => 24,
    4090 => 24,
    4091 => 24,
    4092 => 24,
    4093 => 24,
    4094 => 24,
    4095 => 24,
    4096 => 24,
    4097 => 24,
    4098 => 24,
    4099 => 24,
    4100 => 24,
    4101 => 24,
    4102 => 24,
    4103 => 24,
    4104 => 24,
    4105 => 24,
    4106 => 24,
    4107 => 24,
    4108 => 24,
    4109 => 24,
    4110 => 24,
    4111 => 24,
    4112 => 24,
    4113 => 24,
    4114 => 24,
    4115 => 24,
    4116 => 24,
    4117 => 24,
    4118 => 24,
    4119 => 24,
    4120 => 24,
    4121 => 24,
    4122 => 24,
    4123 => 24,
    4124 => 24,
    4125 => 24,
    4126 => 24,
    4127 => 24,
    4128 => 24,
    4129 => 24,
    4130 => 24,
    4131 => 24,
    4132 => 24,
    4133 => 24,
    4134 => 24,
    4135 => 24,
    4136 => 24,
    4137 => 24,
    4138 => 24,
    4139 => 24,
    4140 => 24,
    4141 => 24,
    4142 => 24,
    4143 => 24,
    4144 => 24,
    4145 => 24,
    4146 => 24,
    4147 => 24,
    4148 => 24,
    4149 => 24,
    4150 => 24,
    4151 => 24,
    4152 => 24,
    4153 => 24,
    4154 => 24,
    4155 => 24,
    4156 => 24,
    4157 => 24,
    4158 => 24,
    4159 => 24,
    4160 => 24,
    4161 => 24,
    4162 => 24,
    4163 => 24,
    4164 => 24,
    4165 => 24,
    4166 => 24,
    4167 => 25,
    4168 => 25,
    4169 => 25,
    4170 => 25,
    4171 => 25,
    4172 => 25,
    4173 => 25,
    4174 => 25,
    4175 => 25,
    4176 => 25,
    4177 => 25,
    4178 => 25,
    4179 => 25,
    4180 => 25,
    4181 => 25,
    4182 => 25,
    4183 => 25,
    4184 => 25,
    4185 => 25,
    4186 => 25,
    4187 => 25,
    4188 => 25,
    4189 => 25,
    4190 => 25,
    4191 => 25,
    4192 => 25,
    4193 => 25,
    4194 => 25,
    4195 => 25,
    4196 => 25,
    4197 => 25,
    4198 => 25,
    4199 => 25,
    4200 => 25,
    4201 => 25,
    4202 => 25,
    4203 => 25,
    4204 => 25,
    4205 => 25,
    4206 => 25,
    4207 => 25,
    4208 => 25,
    4209 => 25,
    4210 => 25,
    4211 => 25,
    4212 => 25,
    4213 => 25,
    4214 => 25,
    4215 => 25,
    4216 => 25,
    4217 => 25,
    4218 => 25,
    4219 => 25,
    4220 => 25,
    4221 => 25,
    4222 => 25,
    4223 => 25,
    4224 => 25,
    4225 => 25,
    4226 => 25,
    4227 => 25,
    4228 => 25,
    4229 => 25,
    4230 => 25,
    4231 => 25,
    4232 => 25,
    4233 => 25,
    4234 => 25,
    4235 => 25,
    4236 => 25,
    4237 => 25,
    4238 => 25,
    4239 => 25,
    4240 => 25,
    4241 => 25,
    4242 => 25,
    4243 => 25,
    4244 => 25,
    4245 => 25,
    4246 => 25,
    4247 => 25,
    4248 => 25,
    4249 => 25,
    4250 => 25,
    4251 => 25,
    4252 => 25,
    4253 => 25,
    4254 => 25,
    4255 => 25,
    4256 => 25,
    4257 => 25,
    4258 => 25,
    4259 => 25,
    4260 => 25,
    4261 => 25,
    4262 => 25,
    4263 => 25,
    4264 => 25,
    4265 => 25,
    4266 => 25,
    4267 => 25,
    4268 => 25,
    4269 => 25,
    4270 => 25,
    4271 => 25,
    4272 => 25,
    4273 => 25,
    4274 => 25,
    4275 => 25,
    4276 => 25,
    4277 => 25,
    4278 => 25,
    4279 => 25,
    4280 => 25,
    4281 => 25,
    4282 => 25,
    4283 => 25,
    4284 => 25,
    4285 => 25,
    4286 => 25,
    4287 => 25,
    4288 => 25,
    4289 => 25,
    4290 => 25,
    4291 => 25,
    4292 => 25,
    4293 => 25,
    4294 => 25,
    4295 => 25,
    4296 => 25,
    4297 => 25,
    4298 => 25,
    4299 => 25,
    4300 => 25,
    4301 => 25,
    4302 => 25,
    4303 => 25,
    4304 => 25,
    4305 => 25,
    4306 => 25,
    4307 => 25,
    4308 => 25,
    4309 => 25,
    4310 => 25,
    4311 => 25,
    4312 => 25,
    4313 => 25,
    4314 => 25,
    4315 => 25,
    4316 => 25,
    4317 => 25,
    4318 => 25,
    4319 => 25,
    4320 => 25,
    4321 => 25,
    4322 => 25,
    4323 => 25,
    4324 => 25,
    4325 => 25,
    4326 => 25,
    4327 => 25,
    4328 => 25,
    4329 => 25,
    4330 => 25,
    4331 => 25,
    4332 => 25,
    4333 => 25,
    4334 => 25,
    4335 => 25,
    4336 => 25,
    4337 => 25,
    4338 => 25,
    4339 => 25,
    4340 => 25,
    4341 => 25,
    4342 => 25,
    4343 => 25,
    4344 => 25,
    4345 => 25,
    4346 => 25,
    4347 => 26,
    4348 => 26,
    4349 => 26,
    4350 => 26,
    4351 => 26,
    4352 => 26,
    4353 => 26,
    4354 => 26,
    4355 => 26,
    4356 => 26,
    4357 => 26,
    4358 => 26,
    4359 => 26,
    4360 => 26,
    4361 => 26,
    4362 => 26,
    4363 => 26,
    4364 => 26,
    4365 => 26,
    4366 => 26,
    4367 => 26,
    4368 => 26,
    4369 => 26,
    4370 => 26,
    4371 => 26,
    4372 => 26,
    4373 => 26,
    4374 => 26,
    4375 => 26,
    4376 => 26,
    4377 => 26,
    4378 => 26,
    4379 => 26,
    4380 => 26,
    4381 => 26,
    4382 => 26,
    4383 => 26,
    4384 => 26,
    4385 => 26,
    4386 => 26,
    4387 => 26,
    4388 => 26,
    4389 => 26,
    4390 => 26,
    4391 => 26,
    4392 => 26,
    4393 => 26,
    4394 => 26,
    4395 => 26,
    4396 => 26,
    4397 => 26,
    4398 => 26,
    4399 => 26,
    4400 => 26,
    4401 => 26,
    4402 => 26,
    4403 => 26,
    4404 => 26,
    4405 => 26,
    4406 => 26,
    4407 => 26,
    4408 => 26,
    4409 => 26,
    4410 => 26,
    4411 => 26,
    4412 => 26,
    4413 => 26,
    4414 => 26,
    4415 => 26,
    4416 => 26,
    4417 => 26,
    4418 => 26,
    4419 => 26,
    4420 => 26,
    4421 => 26,
    4422 => 26,
    4423 => 26,
    4424 => 26,
    4425 => 26,
    4426 => 26,
    4427 => 26,
    4428 => 26,
    4429 => 26,
    4430 => 26,
    4431 => 26,
    4432 => 26,
    4433 => 26,
    4434 => 26,
    4435 => 26,
    4436 => 26,
    4437 => 26,
    4438 => 26,
    4439 => 26,
    4440 => 26,
    4441 => 26,
    4442 => 26,
    4443 => 26,
    4444 => 26,
    4445 => 26,
    4446 => 26,
    4447 => 26,
    4448 => 26,
    4449 => 26,
    4450 => 26,
    4451 => 26,
    4452 => 26,
    4453 => 26,
    4454 => 26,
    4455 => 26,
    4456 => 26,
    4457 => 26,
    4458 => 26,
    4459 => 26,
    4460 => 26,
    4461 => 26,
    4462 => 26,
    4463 => 26,
    4464 => 26,
    4465 => 26,
    4466 => 26,
    4467 => 26,
    4468 => 26,
    4469 => 26,
    4470 => 26,
    4471 => 26,
    4472 => 26,
    4473 => 26,
    4474 => 26,
    4475 => 26,
    4476 => 26,
    4477 => 26,
    4478 => 26,
    4479 => 26,
    4480 => 26,
    4481 => 26,
    4482 => 26,
    4483 => 26,
    4484 => 26,
    4485 => 26,
    4486 => 26,
    4487 => 26,
    4488 => 26,
    4489 => 26,
    4490 => 26,
    4491 => 26,
    4492 => 26,
    4493 => 26,
    4494 => 26,
    4495 => 26,
    4496 => 26,
    4497 => 26,
    4498 => 26,
    4499 => 26,
    4500 => 26,
    4501 => 26,
    4502 => 26,
    4503 => 26,
    4504 => 26,
    4505 => 26,
    4506 => 26,
    4507 => 26,
    4508 => 26,
    4509 => 26,
    4510 => 26,
    4511 => 26,
    4512 => 26,
    4513 => 26,
    4514 => 26,
    4515 => 26,
    4516 => 26,
    4517 => 26,
    4518 => 26,
    4519 => 26,
    4520 => 26,
    4521 => 26,
    4522 => 26,
    4523 => 26,
    4524 => 26,
    4525 => 26,
    4526 => 26,
    4527 => 26,
    4528 => 26,
    4529 => 27,
    4530 => 27,
    4531 => 27,
    4532 => 27,
    4533 => 27,
    4534 => 27,
    4535 => 27,
    4536 => 27,
    4537 => 27,
    4538 => 27,
    4539 => 27,
    4540 => 27,
    4541 => 27,
    4542 => 27,
    4543 => 27,
    4544 => 27,
    4545 => 27,
    4546 => 27,
    4547 => 27,
    4548 => 27,
    4549 => 27,
    4550 => 27,
    4551 => 27,
    4552 => 27,
    4553 => 27,
    4554 => 27,
    4555 => 27,
    4556 => 27,
    4557 => 27,
    4558 => 27,
    4559 => 27,
    4560 => 27,
    4561 => 27,
    4562 => 27,
    4563 => 27,
    4564 => 27,
    4565 => 27,
    4566 => 27,
    4567 => 27,
    4568 => 27,
    4569 => 27,
    4570 => 27,
    4571 => 27,
    4572 => 27,
    4573 => 27,
    4574 => 27,
    4575 => 27,
    4576 => 27,
    4577 => 27,
    4578 => 27,
    4579 => 27,
    4580 => 27,
    4581 => 27,
    4582 => 27,
    4583 => 27,
    4584 => 27,
    4585 => 27,
    4586 => 27,
    4587 => 27,
    4588 => 27,
    4589 => 27,
    4590 => 27,
    4591 => 27,
    4592 => 27,
    4593 => 27,
    4594 => 27,
    4595 => 27,
    4596 => 27,
    4597 => 27,
    4598 => 27,
    4599 => 27,
    4600 => 27,
    4601 => 27,
    4602 => 27,
    4603 => 27,
    4604 => 27,
    4605 => 27,
    4606 => 27,
    4607 => 27,
    4608 => 27,
    4609 => 27,
    4610 => 27,
    4611 => 27,
    4612 => 27,
    4613 => 27,
    4614 => 27,
    4615 => 27,
    4616 => 27,
    4617 => 27,
    4618 => 27,
    4619 => 27,
    4620 => 27,
    4621 => 27,
    4622 => 27,
    4623 => 27,
    4624 => 27,
    4625 => 27,
    4626 => 27,
    4627 => 27,
    4628 => 27,
    4629 => 27,
    4630 => 27,
    4631 => 27,
    4632 => 27,
    4633 => 27,
    4634 => 27,
    4635 => 27,
    4636 => 27,
    4637 => 27,
    4638 => 27,
    4639 => 27,
    4640 => 27,
    4641 => 27,
    4642 => 27,
    4643 => 27,
    4644 => 27,
    4645 => 27,
    4646 => 27,
    4647 => 27,
    4648 => 27,
    4649 => 27,
    4650 => 27,
    4651 => 27,
    4652 => 27,
    4653 => 27,
    4654 => 27,
    4655 => 27,
    4656 => 27,
    4657 => 27,
    4658 => 27,
    4659 => 27,
    4660 => 27,
    4661 => 27,
    4662 => 27,
    4663 => 27,
    4664 => 27,
    4665 => 27,
    4666 => 27,
    4667 => 27,
    4668 => 27,
    4669 => 27,
    4670 => 27,
    4671 => 27,
    4672 => 27,
    4673 => 27,
    4674 => 27,
    4675 => 27,
    4676 => 27,
    4677 => 27,
    4678 => 27,
    4679 => 27,
    4680 => 27,
    4681 => 27,
    4682 => 27,
    4683 => 27,
    4684 => 27,
    4685 => 27,
    4686 => 27,
    4687 => 27,
    4688 => 27,
    4689 => 27,
    4690 => 27,
    4691 => 27,
    4692 => 27,
    4693 => 27,
    4694 => 27,
    4695 => 27,
    4696 => 27,
    4697 => 27,
    4698 => 27,
    4699 => 27,
    4700 => 27,
    4701 => 27,
    4702 => 27,
    4703 => 27,
    4704 => 27,
    4705 => 27,
    4706 => 27,
    4707 => 27,
    4708 => 27,
    4709 => 27,
    4710 => 27,
    4711 => 27,
    4712 => 28,
    4713 => 28,
    4714 => 28,
    4715 => 28,
    4716 => 28,
    4717 => 28,
    4718 => 28,
    4719 => 28,
    4720 => 28,
    4721 => 28,
    4722 => 28,
    4723 => 28,
    4724 => 28,
    4725 => 28,
    4726 => 28,
    4727 => 28,
    4728 => 28,
    4729 => 28,
    4730 => 28,
    4731 => 28,
    4732 => 28,
    4733 => 28,
    4734 => 28,
    4735 => 28,
    4736 => 28,
    4737 => 28,
    4738 => 28,
    4739 => 28,
    4740 => 28,
    4741 => 28,
    4742 => 28,
    4743 => 28,
    4744 => 28,
    4745 => 28,
    4746 => 28,
    4747 => 28,
    4748 => 28,
    4749 => 28,
    4750 => 28,
    4751 => 28,
    4752 => 28,
    4753 => 28,
    4754 => 28,
    4755 => 28,
    4756 => 28,
    4757 => 28,
    4758 => 28,
    4759 => 28,
    4760 => 28,
    4761 => 28,
    4762 => 28,
    4763 => 28,
    4764 => 28,
    4765 => 28,
    4766 => 28,
    4767 => 28,
    4768 => 28,
    4769 => 28,
    4770 => 28,
    4771 => 28,
    4772 => 28,
    4773 => 28,
    4774 => 28,
    4775 => 28,
    4776 => 28,
    4777 => 28,
    4778 => 28,
    4779 => 28,
    4780 => 28,
    4781 => 28,
    4782 => 28,
    4783 => 28,
    4784 => 28,
    4785 => 28,
    4786 => 28,
    4787 => 28,
    4788 => 28,
    4789 => 28,
    4790 => 28,
    4791 => 28,
    4792 => 28,
    4793 => 28,
    4794 => 28,
    4795 => 28,
    4796 => 28,
    4797 => 28,
    4798 => 28,
    4799 => 28,
    4800 => 28,
    4801 => 28,
    4802 => 28,
    4803 => 28,
    4804 => 28,
    4805 => 28,
    4806 => 28,
    4807 => 28,
    4808 => 28,
    4809 => 28,
    4810 => 28,
    4811 => 28,
    4812 => 28,
    4813 => 28,
    4814 => 28,
    4815 => 28,
    4816 => 28,
    4817 => 28,
    4818 => 28,
    4819 => 28,
    4820 => 28,
    4821 => 28,
    4822 => 28,
    4823 => 28,
    4824 => 28,
    4825 => 28,
    4826 => 28,
    4827 => 28,
    4828 => 28,
    4829 => 28,
    4830 => 28,
    4831 => 28,
    4832 => 28,
    4833 => 28,
    4834 => 28,
    4835 => 28,
    4836 => 28,
    4837 => 28,
    4838 => 28,
    4839 => 28,
    4840 => 28,
    4841 => 28,
    4842 => 28,
    4843 => 28,
    4844 => 28,
    4845 => 28,
    4846 => 28,
    4847 => 28,
    4848 => 28,
    4849 => 28,
    4850 => 28,
    4851 => 28,
    4852 => 28,
    4853 => 28,
    4854 => 28,
    4855 => 28,
    4856 => 28,
    4857 => 28,
    4858 => 28,
    4859 => 28,
    4860 => 28,
    4861 => 28,
    4862 => 28,
    4863 => 28,
    4864 => 28,
    4865 => 28,
    4866 => 28,
    4867 => 28,
    4868 => 28,
    4869 => 28,
    4870 => 28,
    4871 => 28,
    4872 => 28,
    4873 => 28,
    4874 => 28,
    4875 => 28,
    4876 => 28,
    4877 => 28,
    4878 => 28,
    4879 => 28,
    4880 => 28,
    4881 => 28,
    4882 => 28,
    4883 => 28,
    4884 => 28,
    4885 => 28,
    4886 => 28,
    4887 => 28,
    4888 => 28,
    4889 => 28,
    4890 => 28,
    4891 => 28,
    4892 => 28,
    4893 => 28,
    4894 => 28,
    4895 => 28,
    4896 => 28,
    4897 => 29,
    4898 => 29,
    4899 => 29,
    4900 => 29,
    4901 => 29,
    4902 => 29,
    4903 => 29,
    4904 => 29,
    4905 => 29,
    4906 => 29,
    4907 => 29,
    4908 => 29,
    4909 => 29,
    4910 => 29,
    4911 => 29,
    4912 => 29,
    4913 => 29,
    4914 => 29,
    4915 => 29,
    4916 => 29,
    4917 => 29,
    4918 => 29,
    4919 => 29,
    4920 => 29,
    4921 => 29,
    4922 => 29,
    4923 => 29,
    4924 => 29,
    4925 => 29,
    4926 => 29,
    4927 => 29,
    4928 => 29,
    4929 => 29,
    4930 => 29,
    4931 => 29,
    4932 => 29,
    4933 => 29,
    4934 => 29,
    4935 => 29,
    4936 => 29,
    4937 => 29,
    4938 => 29,
    4939 => 29,
    4940 => 29,
    4941 => 29,
    4942 => 29,
    4943 => 29,
    4944 => 29,
    4945 => 29,
    4946 => 29,
    4947 => 29,
    4948 => 29,
    4949 => 29,
    4950 => 29,
    4951 => 29,
    4952 => 29,
    4953 => 29,
    4954 => 29,
    4955 => 29,
    4956 => 29,
    4957 => 29,
    4958 => 29,
    4959 => 29,
    4960 => 29,
    4961 => 29,
    4962 => 29,
    4963 => 29,
    4964 => 29,
    4965 => 29,
    4966 => 29,
    4967 => 29,
    4968 => 29,
    4969 => 29,
    4970 => 29,
    4971 => 29,
    4972 => 29,
    4973 => 29,
    4974 => 29,
    4975 => 29,
    4976 => 29,
    4977 => 29,
    4978 => 29,
    4979 => 29,
    4980 => 29,
    4981 => 29,
    4982 => 29,
    4983 => 29,
    4984 => 29,
    4985 => 29,
    4986 => 29,
    4987 => 29,
    4988 => 29,
    4989 => 29,
    4990 => 29,
    4991 => 29,
    4992 => 29,
    4993 => 29,
    4994 => 29,
    4995 => 29,
    4996 => 29,
    4997 => 29,
    4998 => 29,
    4999 => 29,
    5000 => 29,
    5001 => 29,
    5002 => 29,
    5003 => 29,
    5004 => 29,
    5005 => 29,
    5006 => 29,
    5007 => 29,
    5008 => 29,
    5009 => 29,
    5010 => 29,
    5011 => 29,
    5012 => 29,
    5013 => 29,
    5014 => 29,
    5015 => 29,
    5016 => 29,
    5017 => 29,
    5018 => 29,
    5019 => 29,
    5020 => 29,
    5021 => 29,
    5022 => 29,
    5023 => 29,
    5024 => 29,
    5025 => 29,
    5026 => 29,
    5027 => 29,
    5028 => 29,
    5029 => 29,
    5030 => 29,
    5031 => 29,
    5032 => 29,
    5033 => 29,
    5034 => 29,
    5035 => 29,
    5036 => 29,
    5037 => 29,
    5038 => 29,
    5039 => 29,
    5040 => 29,
    5041 => 29,
    5042 => 29,
    5043 => 29,
    5044 => 29,
    5045 => 29,
    5046 => 29,
    5047 => 29,
    5048 => 29,
    5049 => 29,
    5050 => 29,
    5051 => 29,
    5052 => 29,
    5053 => 29,
    5054 => 29,
    5055 => 29,
    5056 => 29,
    5057 => 29,
    5058 => 29,
    5059 => 29,
    5060 => 29,
    5061 => 29,
    5062 => 29,
    5063 => 29,
    5064 => 29,
    5065 => 29,
    5066 => 29,
    5067 => 29,
    5068 => 29,
    5069 => 29,
    5070 => 29,
    5071 => 29,
    5072 => 29,
    5073 => 29,
    5074 => 29,
    5075 => 29,
    5076 => 29,
    5077 => 29,
    5078 => 29,
    5079 => 29,
    5080 => 29,
    5081 => 29,
    5082 => 29,
    5083 => 30,
    5084 => 30,
    5085 => 30,
    5086 => 30,
    5087 => 30,
    5088 => 30,
    5089 => 30,
    5090 => 30,
    5091 => 30,
    5092 => 30,
    5093 => 30,
    5094 => 30,
    5095 => 30,
    5096 => 30,
    5097 => 30,
    5098 => 30,
    5099 => 30,
    5100 => 30,
    5101 => 30,
    5102 => 30,
    5103 => 30,
    5104 => 30,
    5105 => 30,
    5106 => 30,
    5107 => 30,
    5108 => 30,
    5109 => 30,
    5110 => 30,
    5111 => 30,
    5112 => 30,
    5113 => 30,
    5114 => 30,
    5115 => 30,
    5116 => 30,
    5117 => 30,
    5118 => 30,
    5119 => 30,
    5120 => 30,
    5121 => 30,
    5122 => 30,
    5123 => 30,
    5124 => 30,
    5125 => 30,
    5126 => 30,
    5127 => 30,
    5128 => 30,
    5129 => 30,
    5130 => 30,
    5131 => 30,
    5132 => 30,
    5133 => 30,
    5134 => 30,
    5135 => 30,
    5136 => 30,
    5137 => 30,
    5138 => 30,
    5139 => 30,
    5140 => 30,
    5141 => 30,
    5142 => 30,
    5143 => 30,
    5144 => 30,
    5145 => 30,
    5146 => 30,
    5147 => 30,
    5148 => 30,
    5149 => 30,
    5150 => 30,
    5151 => 30,
    5152 => 30,
    5153 => 30,
    5154 => 30,
    5155 => 30,
    5156 => 30,
    5157 => 30,
    5158 => 30,
    5159 => 30,
    5160 => 30,
    5161 => 30,
    5162 => 30,
    5163 => 30,
    5164 => 30,
    5165 => 30,
    5166 => 30,
    5167 => 30,
    5168 => 30,
    5169 => 30,
    5170 => 30,
    5171 => 30,
    5172 => 30,
    5173 => 30,
    5174 => 30,
    5175 => 30,
    5176 => 30,
    5177 => 30,
    5178 => 30,
    5179 => 30,
    5180 => 30,
    5181 => 30,
    5182 => 30,
    5183 => 30,
    5184 => 30,
    5185 => 30,
    5186 => 30,
    5187 => 30,
    5188 => 30,
    5189 => 30,
    5190 => 30,
    5191 => 30,
    5192 => 30,
    5193 => 30,
    5194 => 30,
    5195 => 30,
    5196 => 30,
    5197 => 30,
    5198 => 30,
    5199 => 30,
    5200 => 30,
    5201 => 30,
    5202 => 30,
    5203 => 30,
    5204 => 30,
    5205 => 30,
    5206 => 30,
    5207 => 30,
    5208 => 30,
    5209 => 30,
    5210 => 30,
    5211 => 30,
    5212 => 30,
    5213 => 30,
    5214 => 30,
    5215 => 30,
    5216 => 30,
    5217 => 30,
    5218 => 30,
    5219 => 30,
    5220 => 30,
    5221 => 30,
    5222 => 30,
    5223 => 30,
    5224 => 30,
    5225 => 30,
    5226 => 30,
    5227 => 30,
    5228 => 30,
    5229 => 30,
    5230 => 30,
    5231 => 30,
    5232 => 30,
    5233 => 30,
    5234 => 30,
    5235 => 30,
    5236 => 30,
    5237 => 30,
    5238 => 30,
    5239 => 30,
    5240 => 30,
    5241 => 30,
    5242 => 30,
    5243 => 30,
    5244 => 30,
    5245 => 30,
    5246 => 30,
    5247 => 30,
    5248 => 30,
    5249 => 30,
    5250 => 30,
    5251 => 30,
    5252 => 30,
    5253 => 30,
    5254 => 30,
    5255 => 30,
    5256 => 30,
    5257 => 30,
    5258 => 30,
    5259 => 30,
    5260 => 30,
    5261 => 30,
    5262 => 30,
    5263 => 30,
    5264 => 30,
    5265 => 30,
    5266 => 30,
    5267 => 30,
    5268 => 30,
    5269 => 30,
    5270 => 30,
    5271 => 30,
    5272 => 31,
    5273 => 31,
    5274 => 31,
    5275 => 31,
    5276 => 31,
    5277 => 31,
    5278 => 31,
    5279 => 31,
    5280 => 31,
    5281 => 31,
    5282 => 31,
    5283 => 31,
    5284 => 31,
    5285 => 31,
    5286 => 31,
    5287 => 31,
    5288 => 31,
    5289 => 31,
    5290 => 31,
    5291 => 31,
    5292 => 31,
    5293 => 31,
    5294 => 31,
    5295 => 31,
    5296 => 31,
    5297 => 31,
    5298 => 31,
    5299 => 31,
    5300 => 31,
    5301 => 31,
    5302 => 31,
    5303 => 31,
    5304 => 31,
    5305 => 31,
    5306 => 31,
    5307 => 31,
    5308 => 31,
    5309 => 31,
    5310 => 31,
    5311 => 31,
    5312 => 31,
    5313 => 31,
    5314 => 31,
    5315 => 31,
    5316 => 31,
    5317 => 31,
    5318 => 31,
    5319 => 31,
    5320 => 31,
    5321 => 31,
    5322 => 31,
    5323 => 31,
    5324 => 31,
    5325 => 31,
    5326 => 31,
    5327 => 31,
    5328 => 31,
    5329 => 31,
    5330 => 31,
    5331 => 31,
    5332 => 31,
    5333 => 31,
    5334 => 31,
    5335 => 31,
    5336 => 31,
    5337 => 31,
    5338 => 31,
    5339 => 31,
    5340 => 31,
    5341 => 31,
    5342 => 31,
    5343 => 31,
    5344 => 31,
    5345 => 31,
    5346 => 31,
    5347 => 31,
    5348 => 31,
    5349 => 31,
    5350 => 31,
    5351 => 31,
    5352 => 31,
    5353 => 31,
    5354 => 31,
    5355 => 31,
    5356 => 31,
    5357 => 31,
    5358 => 31,
    5359 => 31,
    5360 => 31,
    5361 => 31,
    5362 => 31,
    5363 => 31,
    5364 => 31,
    5365 => 31,
    5366 => 31,
    5367 => 31,
    5368 => 31,
    5369 => 31,
    5370 => 31,
    5371 => 31,
    5372 => 31,
    5373 => 31,
    5374 => 31,
    5375 => 31,
    5376 => 31,
    5377 => 31,
    5378 => 31,
    5379 => 31,
    5380 => 31,
    5381 => 31,
    5382 => 31,
    5383 => 31,
    5384 => 31,
    5385 => 31,
    5386 => 31,
    5387 => 31,
    5388 => 31,
    5389 => 31,
    5390 => 31,
    5391 => 31,
    5392 => 31,
    5393 => 31,
    5394 => 31,
    5395 => 31,
    5396 => 31,
    5397 => 31,
    5398 => 31,
    5399 => 31,
    5400 => 31,
    5401 => 31,
    5402 => 31,
    5403 => 31,
    5404 => 31,
    5405 => 31,
    5406 => 31,
    5407 => 31,
    5408 => 31,
    5409 => 31,
    5410 => 31,
    5411 => 31,
    5412 => 31,
    5413 => 31,
    5414 => 31,
    5415 => 31,
    5416 => 31,
    5417 => 31,
    5418 => 31,
    5419 => 31,
    5420 => 31,
    5421 => 31,
    5422 => 31,
    5423 => 31,
    5424 => 31,
    5425 => 31,
    5426 => 31,
    5427 => 31,
    5428 => 31,
    5429 => 31,
    5430 => 31,
    5431 => 31,
    5432 => 31,
    5433 => 31,
    5434 => 31,
    5435 => 31,
    5436 => 31,
    5437 => 31,
    5438 => 31,
    5439 => 31,
    5440 => 31,
    5441 => 31,
    5442 => 31,
    5443 => 31,
    5444 => 31,
    5445 => 31,
    5446 => 31,
    5447 => 31,
    5448 => 31,
    5449 => 31,
    5450 => 31,
    5451 => 31,
    5452 => 31,
    5453 => 31,
    5454 => 31,
    5455 => 31,
    5456 => 31,
    5457 => 31,
    5458 => 31,
    5459 => 31,
    5460 => 31,
    5461 => 31,
    5462 => 32,
    5463 => 32,
    5464 => 32,
    5465 => 32,
    5466 => 32,
    5467 => 32,
    5468 => 32,
    5469 => 32,
    5470 => 32,
    5471 => 32,
    5472 => 32,
    5473 => 32,
    5474 => 32,
    5475 => 32,
    5476 => 32,
    5477 => 32,
    5478 => 32,
    5479 => 32,
    5480 => 32,
    5481 => 32,
    5482 => 32,
    5483 => 32,
    5484 => 32,
    5485 => 32,
    5486 => 32,
    5487 => 32,
    5488 => 32,
    5489 => 32,
    5490 => 32,
    5491 => 32,
    5492 => 32,
    5493 => 32,
    5494 => 32,
    5495 => 32,
    5496 => 32,
    5497 => 32,
    5498 => 32,
    5499 => 32,
    5500 => 32,
    5501 => 32,
    5502 => 32,
    5503 => 32,
    5504 => 32,
    5505 => 32,
    5506 => 32,
    5507 => 32,
    5508 => 32,
    5509 => 32,
    5510 => 32,
    5511 => 32,
    5512 => 32,
    5513 => 32,
    5514 => 32,
    5515 => 32,
    5516 => 32,
    5517 => 32,
    5518 => 32,
    5519 => 32,
    5520 => 32,
    5521 => 32,
    5522 => 32,
    5523 => 32,
    5524 => 32,
    5525 => 32,
    5526 => 32,
    5527 => 32,
    5528 => 32,
    5529 => 32,
    5530 => 32,
    5531 => 32,
    5532 => 32,
    5533 => 32,
    5534 => 32,
    5535 => 32,
    5536 => 32,
    5537 => 32,
    5538 => 32,
    5539 => 32,
    5540 => 32,
    5541 => 32,
    5542 => 32,
    5543 => 32,
    5544 => 32,
    5545 => 32,
    5546 => 32,
    5547 => 32,
    5548 => 32,
    5549 => 32,
    5550 => 32,
    5551 => 32,
    5552 => 32,
    5553 => 32,
    5554 => 32,
    5555 => 32,
    5556 => 32,
    5557 => 32,
    5558 => 32,
    5559 => 32,
    5560 => 32,
    5561 => 32,
    5562 => 32,
    5563 => 32,
    5564 => 32,
    5565 => 32,
    5566 => 32,
    5567 => 32,
    5568 => 32,
    5569 => 32,
    5570 => 32,
    5571 => 32,
    5572 => 32,
    5573 => 32,
    5574 => 32,
    5575 => 32,
    5576 => 32,
    5577 => 32,
    5578 => 32,
    5579 => 32,
    5580 => 32,
    5581 => 32,
    5582 => 32,
    5583 => 32,
    5584 => 32,
    5585 => 32,
    5586 => 32,
    5587 => 32,
    5588 => 32,
    5589 => 32,
    5590 => 32,
    5591 => 32,
    5592 => 32,
    5593 => 32,
    5594 => 32,
    5595 => 32,
    5596 => 32,
    5597 => 32,
    5598 => 32,
    5599 => 32,
    5600 => 32,
    5601 => 32,
    5602 => 32,
    5603 => 32,
    5604 => 32,
    5605 => 32,
    5606 => 32,
    5607 => 32,
    5608 => 32,
    5609 => 32,
    5610 => 32,
    5611 => 32,
    5612 => 32,
    5613 => 32,
    5614 => 32,
    5615 => 32,
    5616 => 32,
    5617 => 32,
    5618 => 32,
    5619 => 32,
    5620 => 32,
    5621 => 32,
    5622 => 32,
    5623 => 32,
    5624 => 32,
    5625 => 32,
    5626 => 32,
    5627 => 32,
    5628 => 32,
    5629 => 32,
    5630 => 32,
    5631 => 32,
    5632 => 32,
    5633 => 32,
    5634 => 32,
    5635 => 32,
    5636 => 32,
    5637 => 32,
    5638 => 32,
    5639 => 32,
    5640 => 32,
    5641 => 32,
    5642 => 32,
    5643 => 32,
    5644 => 32,
    5645 => 32,
    5646 => 32,
    5647 => 32,
    5648 => 32,
    5649 => 32,
    5650 => 32,
    5651 => 32,
    5652 => 32,
    5653 => 32,
    5654 => 33,
    5655 => 33,
    5656 => 33,
    5657 => 33,
    5658 => 33,
    5659 => 33,
    5660 => 33,
    5661 => 33,
    5662 => 33,
    5663 => 33,
    5664 => 33,
    5665 => 33,
    5666 => 33,
    5667 => 33,
    5668 => 33,
    5669 => 33,
    5670 => 33,
    5671 => 33,
    5672 => 33,
    5673 => 33,
    5674 => 33,
    5675 => 33,
    5676 => 33,
    5677 => 33,
    5678 => 33,
    5679 => 33,
    5680 => 33,
    5681 => 33,
    5682 => 33,
    5683 => 33,
    5684 => 33,
    5685 => 33,
    5686 => 33,
    5687 => 33,
    5688 => 33,
    5689 => 33,
    5690 => 33,
    5691 => 33,
    5692 => 33,
    5693 => 33,
    5694 => 33,
    5695 => 33,
    5696 => 33,
    5697 => 33,
    5698 => 33,
    5699 => 33,
    5700 => 33,
    5701 => 33,
    5702 => 33,
    5703 => 33,
    5704 => 33,
    5705 => 33,
    5706 => 33,
    5707 => 33,
    5708 => 33,
    5709 => 33,
    5710 => 33,
    5711 => 33,
    5712 => 33,
    5713 => 33,
    5714 => 33,
    5715 => 33,
    5716 => 33,
    5717 => 33,
    5718 => 33,
    5719 => 33,
    5720 => 33,
    5721 => 33,
    5722 => 33,
    5723 => 33,
    5724 => 33,
    5725 => 33,
    5726 => 33,
    5727 => 33,
    5728 => 33,
    5729 => 33,
    5730 => 33,
    5731 => 33,
    5732 => 33,
    5733 => 33,
    5734 => 33,
    5735 => 33,
    5736 => 33,
    5737 => 33,
    5738 => 33,
    5739 => 33,
    5740 => 33,
    5741 => 33,
    5742 => 33,
    5743 => 33,
    5744 => 33,
    5745 => 33,
    5746 => 33,
    5747 => 33,
    5748 => 33,
    5749 => 33,
    5750 => 33,
    5751 => 33,
    5752 => 33,
    5753 => 33,
    5754 => 33,
    5755 => 33,
    5756 => 33,
    5757 => 33,
    5758 => 33,
    5759 => 33,
    5760 => 33,
    5761 => 33,
    5762 => 33,
    5763 => 33,
    5764 => 33,
    5765 => 33,
    5766 => 33,
    5767 => 33,
    5768 => 33,
    5769 => 33,
    5770 => 33,
    5771 => 33,
    5772 => 33,
    5773 => 33,
    5774 => 33,
    5775 => 33,
    5776 => 33,
    5777 => 33,
    5778 => 33,
    5779 => 33,
    5780 => 33,
    5781 => 33,
    5782 => 33,
    5783 => 33,
    5784 => 33,
    5785 => 33,
    5786 => 33,
    5787 => 33,
    5788 => 33,
    5789 => 33,
    5790 => 33,
    5791 => 33,
    5792 => 33,
    5793 => 33,
    5794 => 33,
    5795 => 33,
    5796 => 33,
    5797 => 33,
    5798 => 33,
    5799 => 33,
    5800 => 33,
    5801 => 33,
    5802 => 33,
    5803 => 33,
    5804 => 33,
    5805 => 33,
    5806 => 33,
    5807 => 33,
    5808 => 33,
    5809 => 33,
    5810 => 33,
    5811 => 33,
    5812 => 33,
    5813 => 33,
    5814 => 33,
    5815 => 33,
    5816 => 33,
    5817 => 33,
    5818 => 33,
    5819 => 33,
    5820 => 33,
    5821 => 33,
    5822 => 33,
    5823 => 33,
    5824 => 33,
    5825 => 33,
    5826 => 33,
    5827 => 33,
    5828 => 33,
    5829 => 33,
    5830 => 33,
    5831 => 33,
    5832 => 33,
    5833 => 33,
    5834 => 33,
    5835 => 33,
    5836 => 33,
    5837 => 33,
    5838 => 33,
    5839 => 33,
    5840 => 33,
    5841 => 33,
    5842 => 33,
    5843 => 33,
    5844 => 33,
    5845 => 33,
    5846 => 33,
    5847 => 33,
    5848 => 34,
    5849 => 34,
    5850 => 34,
    5851 => 34,
    5852 => 34,
    5853 => 34,
    5854 => 34,
    5855 => 34,
    5856 => 34,
    5857 => 34,
    5858 => 34,
    5859 => 34,
    5860 => 34,
    5861 => 34,
    5862 => 34,
    5863 => 34,
    5864 => 34,
    5865 => 34,
    5866 => 34,
    5867 => 34,
    5868 => 34,
    5869 => 34,
    5870 => 34,
    5871 => 34,
    5872 => 34,
    5873 => 34,
    5874 => 34,
    5875 => 34,
    5876 => 34,
    5877 => 34,
    5878 => 34,
    5879 => 34,
    5880 => 34,
    5881 => 34,
    5882 => 34,
    5883 => 34,
    5884 => 34,
    5885 => 34,
    5886 => 34,
    5887 => 34,
    5888 => 34,
    5889 => 34,
    5890 => 34,
    5891 => 34,
    5892 => 34,
    5893 => 34,
    5894 => 34,
    5895 => 34,
    5896 => 34,
    5897 => 34,
    5898 => 34,
    5899 => 34,
    5900 => 34,
    5901 => 34,
    5902 => 34,
    5903 => 34,
    5904 => 34,
    5905 => 34,
    5906 => 34,
    5907 => 34,
    5908 => 34,
    5909 => 34,
    5910 => 34,
    5911 => 34,
    5912 => 34,
    5913 => 34,
    5914 => 34,
    5915 => 34,
    5916 => 34,
    5917 => 34,
    5918 => 34,
    5919 => 34,
    5920 => 34,
    5921 => 34,
    5922 => 34,
    5923 => 34,
    5924 => 34,
    5925 => 34,
    5926 => 34,
    5927 => 34,
    5928 => 34,
    5929 => 34,
    5930 => 34,
    5931 => 34,
    5932 => 34,
    5933 => 34,
    5934 => 34,
    5935 => 34,
    5936 => 34,
    5937 => 34,
    5938 => 34,
    5939 => 34,
    5940 => 34,
    5941 => 34,
    5942 => 34,
    5943 => 34,
    5944 => 34,
    5945 => 34,
    5946 => 34,
    5947 => 34,
    5948 => 34,
    5949 => 34,
    5950 => 34,
    5951 => 34,
    5952 => 34,
    5953 => 34,
    5954 => 34,
    5955 => 34,
    5956 => 34,
    5957 => 34,
    5958 => 34,
    5959 => 34,
    5960 => 34,
    5961 => 34,
    5962 => 34,
    5963 => 34,
    5964 => 34,
    5965 => 34,
    5966 => 34,
    5967 => 34,
    5968 => 34,
    5969 => 34,
    5970 => 34,
    5971 => 34,
    5972 => 34,
    5973 => 34,
    5974 => 34,
    5975 => 34,
    5976 => 34,
    5977 => 34,
    5978 => 34,
    5979 => 34,
    5980 => 34,
    5981 => 34,
    5982 => 34,
    5983 => 34,
    5984 => 34,
    5985 => 34,
    5986 => 34,
    5987 => 34,
    5988 => 34,
    5989 => 34,
    5990 => 34,
    5991 => 34,
    5992 => 34,
    5993 => 34,
    5994 => 34,
    5995 => 34,
    5996 => 34,
    5997 => 34,
    5998 => 34,
    5999 => 34,
    6000 => 34,
    6001 => 34,
    6002 => 34,
    6003 => 34,
    6004 => 34,
    6005 => 34,
    6006 => 34,
    6007 => 34,
    6008 => 34,
    6009 => 34,
    6010 => 34,
    6011 => 34,
    6012 => 34,
    6013 => 34,
    6014 => 34,
    6015 => 34,
    6016 => 34,
    6017 => 34,
    6018 => 34,
    6019 => 34,
    6020 => 34,
    6021 => 34,
    6022 => 34,
    6023 => 34,
    6024 => 34,
    6025 => 34,
    6026 => 34,
    6027 => 34,
    6028 => 34,
    6029 => 34,
    6030 => 34,
    6031 => 34,
    6032 => 34,
    6033 => 34,
    6034 => 34,
    6035 => 34,
    6036 => 34,
    6037 => 34,
    6038 => 34,
    6039 => 34,
    6040 => 34,
    6041 => 34,
    6042 => 34,
    6043 => 34,
    6044 => 34,
    6045 => 35,
    6046 => 35,
    6047 => 35,
    6048 => 35,
    6049 => 35,
    6050 => 35,
    6051 => 35,
    6052 => 35,
    6053 => 35,
    6054 => 35,
    6055 => 35,
    6056 => 35,
    6057 => 35,
    6058 => 35,
    6059 => 35,
    6060 => 35,
    6061 => 35,
    6062 => 35,
    6063 => 35,
    6064 => 35,
    6065 => 35,
    6066 => 35,
    6067 => 35,
    6068 => 35,
    6069 => 35,
    6070 => 35,
    6071 => 35,
    6072 => 35,
    6073 => 35,
    6074 => 35,
    6075 => 35,
    6076 => 35,
    6077 => 35,
    6078 => 35,
    6079 => 35,
    6080 => 35,
    6081 => 35,
    6082 => 35,
    6083 => 35,
    6084 => 35,
    6085 => 35,
    6086 => 35,
    6087 => 35,
    6088 => 35,
    6089 => 35,
    6090 => 35,
    6091 => 35,
    6092 => 35,
    6093 => 35,
    6094 => 35,
    6095 => 35,
    6096 => 35,
    6097 => 35,
    6098 => 35,
    6099 => 35,
    6100 => 35,
    6101 => 35,
    6102 => 35,
    6103 => 35,
    6104 => 35,
    6105 => 35,
    6106 => 35,
    6107 => 35,
    6108 => 35,
    6109 => 35,
    6110 => 35,
    6111 => 35,
    6112 => 35,
    6113 => 35,
    6114 => 35,
    6115 => 35,
    6116 => 35,
    6117 => 35,
    6118 => 35,
    6119 => 35,
    6120 => 35,
    6121 => 35,
    6122 => 35,
    6123 => 35,
    6124 => 35,
    6125 => 35,
    6126 => 35,
    6127 => 35,
    6128 => 35,
    6129 => 35,
    6130 => 35,
    6131 => 35,
    6132 => 35,
    6133 => 35,
    6134 => 35,
    6135 => 35,
    6136 => 35,
    6137 => 35,
    6138 => 35,
    6139 => 35,
    6140 => 35,
    6141 => 35,
    6142 => 35,
    6143 => 35,
    6144 => 35,
    6145 => 35,
    6146 => 35,
    6147 => 35,
    6148 => 35,
    6149 => 35,
    6150 => 35,
    6151 => 35,
    6152 => 35,
    6153 => 35,
    6154 => 35,
    6155 => 35,
    6156 => 35,
    6157 => 35,
    6158 => 35,
    6159 => 35,
    6160 => 35,
    6161 => 35,
    6162 => 35,
    6163 => 35,
    6164 => 35,
    6165 => 35,
    6166 => 35,
    6167 => 35,
    6168 => 35,
    6169 => 35,
    6170 => 35,
    6171 => 35,
    6172 => 35,
    6173 => 35,
    6174 => 35,
    6175 => 35,
    6176 => 35,
    6177 => 35,
    6178 => 35,
    6179 => 35,
    6180 => 35,
    6181 => 35,
    6182 => 35,
    6183 => 35,
    6184 => 35,
    6185 => 35,
    6186 => 35,
    6187 => 35,
    6188 => 35,
    6189 => 35,
    6190 => 35,
    6191 => 35,
    6192 => 35,
    6193 => 35,
    6194 => 35,
    6195 => 35,
    6196 => 35,
    6197 => 35,
    6198 => 35,
    6199 => 35,
    6200 => 35,
    6201 => 35,
    6202 => 35,
    6203 => 35,
    6204 => 35,
    6205 => 35,
    6206 => 35,
    6207 => 35,
    6208 => 35,
    6209 => 35,
    6210 => 35,
    6211 => 35,
    6212 => 35,
    6213 => 35,
    6214 => 35,
    6215 => 35,
    6216 => 35,
    6217 => 35,
    6218 => 35,
    6219 => 35,
    6220 => 35,
    6221 => 35,
    6222 => 35,
    6223 => 35,
    6224 => 35,
    6225 => 35,
    6226 => 35,
    6227 => 35,
    6228 => 35,
    6229 => 35,
    6230 => 35,
    6231 => 35,
    6232 => 35,
    6233 => 35,
    6234 => 35,
    6235 => 35,
    6236 => 35,
    6237 => 35,
    6238 => 35,
    6239 => 35,
    6240 => 35,
    6241 => 35,
    6242 => 35,
    6243 => 35,
    6244 => 36,
    6245 => 36,
    6246 => 36,
    6247 => 36,
    6248 => 36,
    6249 => 36,
    6250 => 36,
    6251 => 36,
    6252 => 36,
    6253 => 36,
    6254 => 36,
    6255 => 36,
    6256 => 36,
    6257 => 36,
    6258 => 36,
    6259 => 36,
    6260 => 36,
    6261 => 36,
    6262 => 36,
    6263 => 36,
    6264 => 36,
    6265 => 36,
    6266 => 36,
    6267 => 36,
    6268 => 36,
    6269 => 36,
    6270 => 36,
    6271 => 36,
    6272 => 36,
    6273 => 36,
    6274 => 36,
    6275 => 36,
    6276 => 36,
    6277 => 36,
    6278 => 36,
    6279 => 36,
    6280 => 36,
    6281 => 36,
    6282 => 36,
    6283 => 36,
    6284 => 36,
    6285 => 36,
    6286 => 36,
    6287 => 36,
    6288 => 36,
    6289 => 36,
    6290 => 36,
    6291 => 36,
    6292 => 36,
    6293 => 36,
    6294 => 36,
    6295 => 36,
    6296 => 36,
    6297 => 36,
    6298 => 36,
    6299 => 36,
    6300 => 36,
    6301 => 36,
    6302 => 36,
    6303 => 36,
    6304 => 36,
    6305 => 36,
    6306 => 36,
    6307 => 36,
    6308 => 36,
    6309 => 36,
    6310 => 36,
    6311 => 36,
    6312 => 36,
    6313 => 36,
    6314 => 36,
    6315 => 36,
    6316 => 36,
    6317 => 36,
    6318 => 36,
    6319 => 36,
    6320 => 36,
    6321 => 36,
    6322 => 36,
    6323 => 36,
    6324 => 36,
    6325 => 36,
    6326 => 36,
    6327 => 36,
    6328 => 36,
    6329 => 36,
    6330 => 36,
    6331 => 36,
    6332 => 36,
    6333 => 36,
    6334 => 36,
    6335 => 36,
    6336 => 36,
    6337 => 36,
    6338 => 36,
    6339 => 36,
    6340 => 36,
    6341 => 36,
    6342 => 36,
    6343 => 36,
    6344 => 36,
    6345 => 36,
    6346 => 36,
    6347 => 36,
    6348 => 36,
    6349 => 36,
    6350 => 36,
    6351 => 36,
    6352 => 36,
    6353 => 36,
    6354 => 36,
    6355 => 36,
    6356 => 36,
    6357 => 36,
    6358 => 36,
    6359 => 36,
    6360 => 36,
    6361 => 36,
    6362 => 36,
    6363 => 36,
    6364 => 36,
    6365 => 36,
    6366 => 36,
    6367 => 36,
    6368 => 36,
    6369 => 36,
    6370 => 36,
    6371 => 36,
    6372 => 36,
    6373 => 36,
    6374 => 36,
    6375 => 36,
    6376 => 36,
    6377 => 36,
    6378 => 36,
    6379 => 36,
    6380 => 36,
    6381 => 36,
    6382 => 36,
    6383 => 36,
    6384 => 36,
    6385 => 36,
    6386 => 36,
    6387 => 36,
    6388 => 36,
    6389 => 36,
    6390 => 36,
    6391 => 36,
    6392 => 36,
    6393 => 36,
    6394 => 36,
    6395 => 36,
    6396 => 36,
    6397 => 36,
    6398 => 36,
    6399 => 36,
    6400 => 36,
    6401 => 36,
    6402 => 36,
    6403 => 36,
    6404 => 36,
    6405 => 36,
    6406 => 36,
    6407 => 36,
    6408 => 36,
    6409 => 36,
    6410 => 36,
    6411 => 36,
    6412 => 36,
    6413 => 36,
    6414 => 36,
    6415 => 36,
    6416 => 36,
    6417 => 36,
    6418 => 36,
    6419 => 36,
    6420 => 36,
    6421 => 36,
    6422 => 36,
    6423 => 36,
    6424 => 36,
    6425 => 36,
    6426 => 36,
    6427 => 36,
    6428 => 36,
    6429 => 36,
    6430 => 36,
    6431 => 36,
    6432 => 36,
    6433 => 36,
    6434 => 36,
    6435 => 36,
    6436 => 36,
    6437 => 36,
    6438 => 36,
    6439 => 36,
    6440 => 36,
    6441 => 36,
    6442 => 36,
    6443 => 36,
    6444 => 36,
    6445 => 36,
    6446 => 37,
    6447 => 37,
    6448 => 37,
    6449 => 37,
    6450 => 37,
    6451 => 37,
    6452 => 37,
    6453 => 37,
    6454 => 37,
    6455 => 37,
    6456 => 37,
    6457 => 37,
    6458 => 37,
    6459 => 37,
    6460 => 37,
    6461 => 37,
    6462 => 37,
    6463 => 37,
    6464 => 37,
    6465 => 37,
    6466 => 37,
    6467 => 37,
    6468 => 37,
    6469 => 37,
    6470 => 37,
    6471 => 37,
    6472 => 37,
    6473 => 37,
    6474 => 37,
    6475 => 37,
    6476 => 37,
    6477 => 37,
    6478 => 37,
    6479 => 37,
    6480 => 37,
    6481 => 37,
    6482 => 37,
    6483 => 37,
    6484 => 37,
    6485 => 37,
    6486 => 37,
    6487 => 37,
    6488 => 37,
    6489 => 37,
    6490 => 37,
    6491 => 37,
    6492 => 37,
    6493 => 37,
    6494 => 37,
    6495 => 37,
    6496 => 37,
    6497 => 37,
    6498 => 37,
    6499 => 37,
    6500 => 37,
    6501 => 37,
    6502 => 37,
    6503 => 37,
    6504 => 37,
    6505 => 37,
    6506 => 37,
    6507 => 37,
    6508 => 37,
    6509 => 37,
    6510 => 37,
    6511 => 37,
    6512 => 37,
    6513 => 37,
    6514 => 37,
    6515 => 37,
    6516 => 37,
    6517 => 37,
    6518 => 37,
    6519 => 37,
    6520 => 37,
    6521 => 37,
    6522 => 37,
    6523 => 37,
    6524 => 37,
    6525 => 37,
    6526 => 37,
    6527 => 37,
    6528 => 37,
    6529 => 37,
    6530 => 37,
    6531 => 37,
    6532 => 37,
    6533 => 37,
    6534 => 37,
    6535 => 37,
    6536 => 37,
    6537 => 37,
    6538 => 37,
    6539 => 37,
    6540 => 37,
    6541 => 37,
    6542 => 37,
    6543 => 37,
    6544 => 37,
    6545 => 37,
    6546 => 37,
    6547 => 37,
    6548 => 37,
    6549 => 37,
    6550 => 37,
    6551 => 37,
    6552 => 37,
    6553 => 37,
    6554 => 37,
    6555 => 37,
    6556 => 37,
    6557 => 37,
    6558 => 37,
    6559 => 37,
    6560 => 37,
    6561 => 37,
    6562 => 37,
    6563 => 37,
    6564 => 37,
    6565 => 37,
    6566 => 37,
    6567 => 37,
    6568 => 37,
    6569 => 37,
    6570 => 37,
    6571 => 37,
    6572 => 37,
    6573 => 37,
    6574 => 37,
    6575 => 37,
    6576 => 37,
    6577 => 37,
    6578 => 37,
    6579 => 37,
    6580 => 37,
    6581 => 37,
    6582 => 37,
    6583 => 37,
    6584 => 37,
    6585 => 37,
    6586 => 37,
    6587 => 37,
    6588 => 37,
    6589 => 37,
    6590 => 37,
    6591 => 37,
    6592 => 37,
    6593 => 37,
    6594 => 37,
    6595 => 37,
    6596 => 37,
    6597 => 37,
    6598 => 37,
    6599 => 37,
    6600 => 37,
    6601 => 37,
    6602 => 37,
    6603 => 37,
    6604 => 37,
    6605 => 37,
    6606 => 37,
    6607 => 37,
    6608 => 37,
    6609 => 37,
    6610 => 37,
    6611 => 37,
    6612 => 37,
    6613 => 37,
    6614 => 37,
    6615 => 37,
    6616 => 37,
    6617 => 37,
    6618 => 37,
    6619 => 37,
    6620 => 37,
    6621 => 37,
    6622 => 37,
    6623 => 37,
    6624 => 37,
    6625 => 37,
    6626 => 37,
    6627 => 37,
    6628 => 37,
    6629 => 37,
    6630 => 37,
    6631 => 37,
    6632 => 37,
    6633 => 37,
    6634 => 37,
    6635 => 37,
    6636 => 37,
    6637 => 37,
    6638 => 37,
    6639 => 37,
    6640 => 37,
    6641 => 37,
    6642 => 37,
    6643 => 37,
    6644 => 37,
    6645 => 37,
    6646 => 37,
    6647 => 37,
    6648 => 37,
    6649 => 37,
    6650 => 37,
    6651 => 38,
    6652 => 38,
    6653 => 38,
    6654 => 38,
    6655 => 38,
    6656 => 38,
    6657 => 38,
    6658 => 38,
    6659 => 38,
    6660 => 38,
    6661 => 38,
    6662 => 38,
    6663 => 38,
    6664 => 38,
    6665 => 38,
    6666 => 38,
    6667 => 38,
    6668 => 38,
    6669 => 38,
    6670 => 38,
    6671 => 38,
    6672 => 38,
    6673 => 38,
    6674 => 38,
    6675 => 38,
    6676 => 38,
    6677 => 38,
    6678 => 38,
    6679 => 38,
    6680 => 38,
    6681 => 38,
    6682 => 38,
    6683 => 38,
    6684 => 38,
    6685 => 38,
    6686 => 38,
    6687 => 38,
    6688 => 38,
    6689 => 38,
    6690 => 38,
    6691 => 38,
    6692 => 38,
    6693 => 38,
    6694 => 38,
    6695 => 38,
    6696 => 38,
    6697 => 38,
    6698 => 38,
    6699 => 38,
    6700 => 38,
    6701 => 38,
    6702 => 38,
    6703 => 38,
    6704 => 38,
    6705 => 38,
    6706 => 38,
    6707 => 38,
    6708 => 38,
    6709 => 38,
    6710 => 38,
    6711 => 38,
    6712 => 38,
    6713 => 38,
    6714 => 38,
    6715 => 38,
    6716 => 38,
    6717 => 38,
    6718 => 38,
    6719 => 38,
    6720 => 38,
    6721 => 38,
    6722 => 38,
    6723 => 38,
    6724 => 38,
    6725 => 38,
    6726 => 38,
    6727 => 38,
    6728 => 38,
    6729 => 38,
    6730 => 38,
    6731 => 38,
    6732 => 38,
    6733 => 38,
    6734 => 38,
    6735 => 38,
    6736 => 38,
    6737 => 38,
    6738 => 38,
    6739 => 38,
    6740 => 38,
    6741 => 38,
    6742 => 38,
    6743 => 38,
    6744 => 38,
    6745 => 38,
    6746 => 38,
    6747 => 38,
    6748 => 38,
    6749 => 38,
    6750 => 38,
    6751 => 38,
    6752 => 38,
    6753 => 38,
    6754 => 38,
    6755 => 38,
    6756 => 38,
    6757 => 38,
    6758 => 38,
    6759 => 38,
    6760 => 38,
    6761 => 38,
    6762 => 38,
    6763 => 38,
    6764 => 38,
    6765 => 38,
    6766 => 38,
    6767 => 38,
    6768 => 38,
    6769 => 38,
    6770 => 38,
    6771 => 38,
    6772 => 38,
    6773 => 38,
    6774 => 38,
    6775 => 38,
    6776 => 38,
    6777 => 38,
    6778 => 38,
    6779 => 38,
    6780 => 38,
    6781 => 38,
    6782 => 38,
    6783 => 38,
    6784 => 38,
    6785 => 38,
    6786 => 38,
    6787 => 38,
    6788 => 38,
    6789 => 38,
    6790 => 38,
    6791 => 38,
    6792 => 38,
    6793 => 38,
    6794 => 38,
    6795 => 38,
    6796 => 38,
    6797 => 38,
    6798 => 38,
    6799 => 38,
    6800 => 38,
    6801 => 38,
    6802 => 38,
    6803 => 38,
    6804 => 38,
    6805 => 38,
    6806 => 38,
    6807 => 38,
    6808 => 38,
    6809 => 38,
    6810 => 38,
    6811 => 38,
    6812 => 38,
    6813 => 38,
    6814 => 38,
    6815 => 38,
    6816 => 38,
    6817 => 38,
    6818 => 38,
    6819 => 38,
    6820 => 38,
    6821 => 38,
    6822 => 38,
    6823 => 38,
    6824 => 38,
    6825 => 38,
    6826 => 38,
    6827 => 38,
    6828 => 38,
    6829 => 38,
    6830 => 38,
    6831 => 38,
    6832 => 38,
    6833 => 38,
    6834 => 38,
    6835 => 38,
    6836 => 38,
    6837 => 38,
    6838 => 38,
    6839 => 38,
    6840 => 38,
    6841 => 38,
    6842 => 38,
    6843 => 38,
    6844 => 38,
    6845 => 38,
    6846 => 38,
    6847 => 38,
    6848 => 38,
    6849 => 38,
    6850 => 38,
    6851 => 38,
    6852 => 38,
    6853 => 38,
    6854 => 38,
    6855 => 38,
    6856 => 38,
    6857 => 38,
    6858 => 39,
    6859 => 39,
    6860 => 39,
    6861 => 39,
    6862 => 39,
    6863 => 39,
    6864 => 39,
    6865 => 39,
    6866 => 39,
    6867 => 39,
    6868 => 39,
    6869 => 39,
    6870 => 39,
    6871 => 39,
    6872 => 39,
    6873 => 39,
    6874 => 39,
    6875 => 39,
    6876 => 39,
    6877 => 39,
    6878 => 39,
    6879 => 39,
    6880 => 39,
    6881 => 39,
    6882 => 39,
    6883 => 39,
    6884 => 39,
    6885 => 39,
    6886 => 39,
    6887 => 39,
    6888 => 39,
    6889 => 39,
    6890 => 39,
    6891 => 39,
    6892 => 39,
    6893 => 39,
    6894 => 39,
    6895 => 39,
    6896 => 39,
    6897 => 39,
    6898 => 39,
    6899 => 39,
    6900 => 39,
    6901 => 39,
    6902 => 39,
    6903 => 39,
    6904 => 39,
    6905 => 39,
    6906 => 39,
    6907 => 39,
    6908 => 39,
    6909 => 39,
    6910 => 39,
    6911 => 39,
    6912 => 39,
    6913 => 39,
    6914 => 39,
    6915 => 39,
    6916 => 39,
    6917 => 39,
    6918 => 39,
    6919 => 39,
    6920 => 39,
    6921 => 39,
    6922 => 39,
    6923 => 39,
    6924 => 39,
    6925 => 39,
    6926 => 39,
    6927 => 39,
    6928 => 39,
    6929 => 39,
    6930 => 39,
    6931 => 39,
    6932 => 39,
    6933 => 39,
    6934 => 39,
    6935 => 39,
    6936 => 39,
    6937 => 39,
    6938 => 39,
    6939 => 39,
    6940 => 39,
    6941 => 39,
    6942 => 39,
    6943 => 39,
    6944 => 39,
    6945 => 39,
    6946 => 39,
    6947 => 39,
    6948 => 39,
    6949 => 39,
    6950 => 39,
    6951 => 39,
    6952 => 39,
    6953 => 39,
    6954 => 39,
    6955 => 39,
    6956 => 39,
    6957 => 39,
    6958 => 39,
    6959 => 39,
    6960 => 39,
    6961 => 39,
    6962 => 39,
    6963 => 39,
    6964 => 39,
    6965 => 39,
    6966 => 39,
    6967 => 39,
    6968 => 39,
    6969 => 39,
    6970 => 39,
    6971 => 39,
    6972 => 39,
    6973 => 39,
    6974 => 39,
    6975 => 39,
    6976 => 39,
    6977 => 39,
    6978 => 39,
    6979 => 39,
    6980 => 39,
    6981 => 39,
    6982 => 39,
    6983 => 39,
    6984 => 39,
    6985 => 39,
    6986 => 39,
    6987 => 39,
    6988 => 39,
    6989 => 39,
    6990 => 39,
    6991 => 39,
    6992 => 39,
    6993 => 39,
    6994 => 39,
    6995 => 39,
    6996 => 39,
    6997 => 39,
    6998 => 39,
    6999 => 39,
    7000 => 39,
    7001 => 39,
    7002 => 39,
    7003 => 39,
    7004 => 39,
    7005 => 39,
    7006 => 39,
    7007 => 39,
    7008 => 39,
    7009 => 39,
    7010 => 39,
    7011 => 39,
    7012 => 39,
    7013 => 39,
    7014 => 39,
    7015 => 39,
    7016 => 39,
    7017 => 39,
    7018 => 39,
    7019 => 39,
    7020 => 39,
    7021 => 39,
    7022 => 39,
    7023 => 39,
    7024 => 39,
    7025 => 39,
    7026 => 39,
    7027 => 39,
    7028 => 39,
    7029 => 39,
    7030 => 39,
    7031 => 39,
    7032 => 39,
    7033 => 39,
    7034 => 39,
    7035 => 39,
    7036 => 39,
    7037 => 39,
    7038 => 39,
    7039 => 39,
    7040 => 39,
    7041 => 39,
    7042 => 39,
    7043 => 39,
    7044 => 39,
    7045 => 39,
    7046 => 39,
    7047 => 39,
    7048 => 39,
    7049 => 39,
    7050 => 39,
    7051 => 39,
    7052 => 39,
    7053 => 39,
    7054 => 39,
    7055 => 39,
    7056 => 39,
    7057 => 39,
    7058 => 39,
    7059 => 39,
    7060 => 39,
    7061 => 39,
    7062 => 39,
    7063 => 39,
    7064 => 39,
    7065 => 39,
    7066 => 39,
    7067 => 39,
    7068 => 39,
    7069 => 40,
    7070 => 40,
    7071 => 40,
    7072 => 40,
    7073 => 40,
    7074 => 40,
    7075 => 40,
    7076 => 40,
    7077 => 40,
    7078 => 40,
    7079 => 40,
    7080 => 40,
    7081 => 40,
    7082 => 40,
    7083 => 40,
    7084 => 40,
    7085 => 40,
    7086 => 40,
    7087 => 40,
    7088 => 40,
    7089 => 40,
    7090 => 40,
    7091 => 40,
    7092 => 40,
    7093 => 40,
    7094 => 40,
    7095 => 40,
    7096 => 40,
    7097 => 40,
    7098 => 40,
    7099 => 40,
    7100 => 40,
    7101 => 40,
    7102 => 40,
    7103 => 40,
    7104 => 40,
    7105 => 40,
    7106 => 40,
    7107 => 40,
    7108 => 40,
    7109 => 40,
    7110 => 40,
    7111 => 40,
    7112 => 40,
    7113 => 40,
    7114 => 40,
    7115 => 40,
    7116 => 40,
    7117 => 40,
    7118 => 40,
    7119 => 40,
    7120 => 40,
    7121 => 40,
    7122 => 40,
    7123 => 40,
    7124 => 40,
    7125 => 40,
    7126 => 40,
    7127 => 40,
    7128 => 40,
    7129 => 40,
    7130 => 40,
    7131 => 40,
    7132 => 40,
    7133 => 40,
    7134 => 40,
    7135 => 40,
    7136 => 40,
    7137 => 40,
    7138 => 40,
    7139 => 40,
    7140 => 40,
    7141 => 40,
    7142 => 40,
    7143 => 40,
    7144 => 40,
    7145 => 40,
    7146 => 40,
    7147 => 40,
    7148 => 40,
    7149 => 40,
    7150 => 40,
    7151 => 40,
    7152 => 40,
    7153 => 40,
    7154 => 40,
    7155 => 40,
    7156 => 40,
    7157 => 40,
    7158 => 40,
    7159 => 40,
    7160 => 40,
    7161 => 40,
    7162 => 40,
    7163 => 40,
    7164 => 40,
    7165 => 40,
    7166 => 40,
    7167 => 40,
    7168 => 40,
    7169 => 40,
    7170 => 40,
    7171 => 40,
    7172 => 40,
    7173 => 40,
    7174 => 40,
    7175 => 40,
    7176 => 40,
    7177 => 40,
    7178 => 40,
    7179 => 40,
    7180 => 40,
    7181 => 40,
    7182 => 40,
    7183 => 40,
    7184 => 40,
    7185 => 40,
    7186 => 40,
    7187 => 40,
    7188 => 40,
    7189 => 40,
    7190 => 40,
    7191 => 40,
    7192 => 40,
    7193 => 40,
    7194 => 40,
    7195 => 40,
    7196 => 40,
    7197 => 40,
    7198 => 40,
    7199 => 40,
    7200 => 40,
    7201 => 40,
    7202 => 40,
    7203 => 40,
    7204 => 40,
    7205 => 40,
    7206 => 40,
    7207 => 40,
    7208 => 40,
    7209 => 40,
    7210 => 40,
    7211 => 40,
    7212 => 40,
    7213 => 40,
    7214 => 40,
    7215 => 40,
    7216 => 40,
    7217 => 40,
    7218 => 40,
    7219 => 40,
    7220 => 40,
    7221 => 40,
    7222 => 40,
    7223 => 40,
    7224 => 40,
    7225 => 40,
    7226 => 40,
    7227 => 40,
    7228 => 40,
    7229 => 40,
    7230 => 40,
    7231 => 40,
    7232 => 40,
    7233 => 40,
    7234 => 40,
    7235 => 40,
    7236 => 40,
    7237 => 40,
    7238 => 40,
    7239 => 40,
    7240 => 40,
    7241 => 40,
    7242 => 40,
    7243 => 40,
    7244 => 40,
    7245 => 40,
    7246 => 40,
    7247 => 40,
    7248 => 40,
    7249 => 40,
    7250 => 40,
    7251 => 40,
    7252 => 40,
    7253 => 40,
    7254 => 40,
    7255 => 40,
    7256 => 40,
    7257 => 40,
    7258 => 40,
    7259 => 40,
    7260 => 40,
    7261 => 40,
    7262 => 40,
    7263 => 40,
    7264 => 40,
    7265 => 40,
    7266 => 40,
    7267 => 40,
    7268 => 40,
    7269 => 40,
    7270 => 40,
    7271 => 40,
    7272 => 40,
    7273 => 40,
    7274 => 40,
    7275 => 40,
    7276 => 40,
    7277 => 40,
    7278 => 40,
    7279 => 40,
    7280 => 40,
    7281 => 40,
    7282 => 40,
    7283 => 41,
    7284 => 41,
    7285 => 41,
    7286 => 41,
    7287 => 41,
    7288 => 41,
    7289 => 41,
    7290 => 41,
    7291 => 41,
    7292 => 41,
    7293 => 41,
    7294 => 41,
    7295 => 41,
    7296 => 41,
    7297 => 41,
    7298 => 41,
    7299 => 41,
    7300 => 41,
    7301 => 41,
    7302 => 41,
    7303 => 41,
    7304 => 41,
    7305 => 41,
    7306 => 41,
    7307 => 41,
    7308 => 41,
    7309 => 41,
    7310 => 41,
    7311 => 41,
    7312 => 41,
    7313 => 41,
    7314 => 41,
    7315 => 41,
    7316 => 41,
    7317 => 41,
    7318 => 41,
    7319 => 41,
    7320 => 41,
    7321 => 41,
    7322 => 41,
    7323 => 41,
    7324 => 41,
    7325 => 41,
    7326 => 41,
    7327 => 41,
    7328 => 41,
    7329 => 41,
    7330 => 41,
    7331 => 41,
    7332 => 41,
    7333 => 41,
    7334 => 41,
    7335 => 41,
    7336 => 41,
    7337 => 41,
    7338 => 41,
    7339 => 41,
    7340 => 41,
    7341 => 41,
    7342 => 41,
    7343 => 41,
    7344 => 41,
    7345 => 41,
    7346 => 41,
    7347 => 41,
    7348 => 41,
    7349 => 41,
    7350 => 41,
    7351 => 41,
    7352 => 41,
    7353 => 41,
    7354 => 41,
    7355 => 41,
    7356 => 41,
    7357 => 41,
    7358 => 41,
    7359 => 41,
    7360 => 41,
    7361 => 41,
    7362 => 41,
    7363 => 41,
    7364 => 41,
    7365 => 41,
    7366 => 41,
    7367 => 41,
    7368 => 41,
    7369 => 41,
    7370 => 41,
    7371 => 41,
    7372 => 41,
    7373 => 41,
    7374 => 41,
    7375 => 41,
    7376 => 41,
    7377 => 41,
    7378 => 41,
    7379 => 41,
    7380 => 41,
    7381 => 41,
    7382 => 41,
    7383 => 41,
    7384 => 41,
    7385 => 41,
    7386 => 41,
    7387 => 41,
    7388 => 41,
    7389 => 41,
    7390 => 41,
    7391 => 41,
    7392 => 41,
    7393 => 41,
    7394 => 41,
    7395 => 41,
    7396 => 41,
    7397 => 41,
    7398 => 41,
    7399 => 41,
    7400 => 41,
    7401 => 41,
    7402 => 41,
    7403 => 41,
    7404 => 41,
    7405 => 41,
    7406 => 41,
    7407 => 41,
    7408 => 41,
    7409 => 41,
    7410 => 41,
    7411 => 41,
    7412 => 41,
    7413 => 41,
    7414 => 41,
    7415 => 41,
    7416 => 41,
    7417 => 41,
    7418 => 41,
    7419 => 41,
    7420 => 41,
    7421 => 41,
    7422 => 41,
    7423 => 41,
    7424 => 41,
    7425 => 41,
    7426 => 41,
    7427 => 41,
    7428 => 41,
    7429 => 41,
    7430 => 41,
    7431 => 41,
    7432 => 41,
    7433 => 41,
    7434 => 41,
    7435 => 41,
    7436 => 41,
    7437 => 41,
    7438 => 41,
    7439 => 41,
    7440 => 41,
    7441 => 41,
    7442 => 41,
    7443 => 41,
    7444 => 41,
    7445 => 41,
    7446 => 41,
    7447 => 41,
    7448 => 41,
    7449 => 41,
    7450 => 41,
    7451 => 41,
    7452 => 41,
    7453 => 41,
    7454 => 41,
    7455 => 41,
    7456 => 41,
    7457 => 41,
    7458 => 41,
    7459 => 41,
    7460 => 41,
    7461 => 41,
    7462 => 41,
    7463 => 41,
    7464 => 41,
    7465 => 41,
    7466 => 41,
    7467 => 41,
    7468 => 41,
    7469 => 41,
    7470 => 41,
    7471 => 41,
    7472 => 41,
    7473 => 41,
    7474 => 41,
    7475 => 41,
    7476 => 41,
    7477 => 41,
    7478 => 41,
    7479 => 41,
    7480 => 41,
    7481 => 41,
    7482 => 41,
    7483 => 41,
    7484 => 41,
    7485 => 41,
    7486 => 41,
    7487 => 41,
    7488 => 41,
    7489 => 41,
    7490 => 41,
    7491 => 41,
    7492 => 41,
    7493 => 41,
    7494 => 41,
    7495 => 41,
    7496 => 41,
    7497 => 41,
    7498 => 41,
    7499 => 41,
    7500 => 41,
    7501 => 42,
    7502 => 42,
    7503 => 42,
    7504 => 42,
    7505 => 42,
    7506 => 42,
    7507 => 42,
    7508 => 42,
    7509 => 42,
    7510 => 42,
    7511 => 42,
    7512 => 42,
    7513 => 42,
    7514 => 42,
    7515 => 42,
    7516 => 42,
    7517 => 42,
    7518 => 42,
    7519 => 42,
    7520 => 42,
    7521 => 42,
    7522 => 42,
    7523 => 42,
    7524 => 42,
    7525 => 42,
    7526 => 42,
    7527 => 42,
    7528 => 42,
    7529 => 42,
    7530 => 42,
    7531 => 42,
    7532 => 42,
    7533 => 42,
    7534 => 42,
    7535 => 42,
    7536 => 42,
    7537 => 42,
    7538 => 42,
    7539 => 42,
    7540 => 42,
    7541 => 42,
    7542 => 42,
    7543 => 42,
    7544 => 42,
    7545 => 42,
    7546 => 42,
    7547 => 42,
    7548 => 42,
    7549 => 42,
    7550 => 42,
    7551 => 42,
    7552 => 42,
    7553 => 42,
    7554 => 42,
    7555 => 42,
    7556 => 42,
    7557 => 42,
    7558 => 42,
    7559 => 42,
    7560 => 42,
    7561 => 42,
    7562 => 42,
    7563 => 42,
    7564 => 42,
    7565 => 42,
    7566 => 42,
    7567 => 42,
    7568 => 42,
    7569 => 42,
    7570 => 42,
    7571 => 42,
    7572 => 42,
    7573 => 42,
    7574 => 42,
    7575 => 42,
    7576 => 42,
    7577 => 42,
    7578 => 42,
    7579 => 42,
    7580 => 42,
    7581 => 42,
    7582 => 42,
    7583 => 42,
    7584 => 42,
    7585 => 42,
    7586 => 42,
    7587 => 42,
    7588 => 42,
    7589 => 42,
    7590 => 42,
    7591 => 42,
    7592 => 42,
    7593 => 42,
    7594 => 42,
    7595 => 42,
    7596 => 42,
    7597 => 42,
    7598 => 42,
    7599 => 42,
    7600 => 42,
    7601 => 42,
    7602 => 42,
    7603 => 42,
    7604 => 42,
    7605 => 42,
    7606 => 42,
    7607 => 42,
    7608 => 42,
    7609 => 42,
    7610 => 42,
    7611 => 42,
    7612 => 42,
    7613 => 42,
    7614 => 42,
    7615 => 42,
    7616 => 42,
    7617 => 42,
    7618 => 42,
    7619 => 42,
    7620 => 42,
    7621 => 42,
    7622 => 42,
    7623 => 42,
    7624 => 42,
    7625 => 42,
    7626 => 42,
    7627 => 42,
    7628 => 42,
    7629 => 42,
    7630 => 42,
    7631 => 42,
    7632 => 42,
    7633 => 42,
    7634 => 42,
    7635 => 42,
    7636 => 42,
    7637 => 42,
    7638 => 42,
    7639 => 42,
    7640 => 42,
    7641 => 42,
    7642 => 42,
    7643 => 42,
    7644 => 42,
    7645 => 42,
    7646 => 42,
    7647 => 42,
    7648 => 42,
    7649 => 42,
    7650 => 42,
    7651 => 42,
    7652 => 42,
    7653 => 42,
    7654 => 42,
    7655 => 42,
    7656 => 42,
    7657 => 42,
    7658 => 42,
    7659 => 42,
    7660 => 42,
    7661 => 42,
    7662 => 42,
    7663 => 42,
    7664 => 42,
    7665 => 42,
    7666 => 42,
    7667 => 42,
    7668 => 42,
    7669 => 42,
    7670 => 42,
    7671 => 42,
    7672 => 42,
    7673 => 42,
    7674 => 42,
    7675 => 42,
    7676 => 42,
    7677 => 42,
    7678 => 42,
    7679 => 42,
    7680 => 42,
    7681 => 42,
    7682 => 42,
    7683 => 42,
    7684 => 42,
    7685 => 42,
    7686 => 42,
    7687 => 42,
    7688 => 42,
    7689 => 42,
    7690 => 42,
    7691 => 42,
    7692 => 42,
    7693 => 42,
    7694 => 42,
    7695 => 42,
    7696 => 42,
    7697 => 42,
    7698 => 42,
    7699 => 42,
    7700 => 42,
    7701 => 42,
    7702 => 42,
    7703 => 42,
    7704 => 42,
    7705 => 42,
    7706 => 42,
    7707 => 42,
    7708 => 42,
    7709 => 42,
    7710 => 42,
    7711 => 42,
    7712 => 42,
    7713 => 42,
    7714 => 42,
    7715 => 42,
    7716 => 42,
    7717 => 42,
    7718 => 42,
    7719 => 42,
    7720 => 42,
    7721 => 42,
    7722 => 42,
    7723 => 43,
    7724 => 43,
    7725 => 43,
    7726 => 43,
    7727 => 43,
    7728 => 43,
    7729 => 43,
    7730 => 43,
    7731 => 43,
    7732 => 43,
    7733 => 43,
    7734 => 43,
    7735 => 43,
    7736 => 43,
    7737 => 43,
    7738 => 43,
    7739 => 43,
    7740 => 43,
    7741 => 43,
    7742 => 43,
    7743 => 43,
    7744 => 43,
    7745 => 43,
    7746 => 43,
    7747 => 43,
    7748 => 43,
    7749 => 43,
    7750 => 43,
    7751 => 43,
    7752 => 43,
    7753 => 43,
    7754 => 43,
    7755 => 43,
    7756 => 43,
    7757 => 43,
    7758 => 43,
    7759 => 43,
    7760 => 43,
    7761 => 43,
    7762 => 43,
    7763 => 43,
    7764 => 43,
    7765 => 43,
    7766 => 43,
    7767 => 43,
    7768 => 43,
    7769 => 43,
    7770 => 43,
    7771 => 43,
    7772 => 43,
    7773 => 43,
    7774 => 43,
    7775 => 43,
    7776 => 43,
    7777 => 43,
    7778 => 43,
    7779 => 43,
    7780 => 43,
    7781 => 43,
    7782 => 43,
    7783 => 43,
    7784 => 43,
    7785 => 43,
    7786 => 43,
    7787 => 43,
    7788 => 43,
    7789 => 43,
    7790 => 43,
    7791 => 43,
    7792 => 43,
    7793 => 43,
    7794 => 43,
    7795 => 43,
    7796 => 43,
    7797 => 43,
    7798 => 43,
    7799 => 43,
    7800 => 43,
    7801 => 43,
    7802 => 43,
    7803 => 43,
    7804 => 43,
    7805 => 43,
    7806 => 43,
    7807 => 43,
    7808 => 43,
    7809 => 43,
    7810 => 43,
    7811 => 43,
    7812 => 43,
    7813 => 43,
    7814 => 43,
    7815 => 43,
    7816 => 43,
    7817 => 43,
    7818 => 43,
    7819 => 43,
    7820 => 43,
    7821 => 43,
    7822 => 43,
    7823 => 43,
    7824 => 43,
    7825 => 43,
    7826 => 43,
    7827 => 43,
    7828 => 43,
    7829 => 43,
    7830 => 43,
    7831 => 43,
    7832 => 43,
    7833 => 43,
    7834 => 43,
    7835 => 43,
    7836 => 43,
    7837 => 43,
    7838 => 43,
    7839 => 43,
    7840 => 43,
    7841 => 43,
    7842 => 43,
    7843 => 43,
    7844 => 43,
    7845 => 43,
    7846 => 43,
    7847 => 43,
    7848 => 43,
    7849 => 43,
    7850 => 43,
    7851 => 43,
    7852 => 43,
    7853 => 43,
    7854 => 43,
    7855 => 43,
    7856 => 43,
    7857 => 43,
    7858 => 43,
    7859 => 43,
    7860 => 43,
    7861 => 43,
    7862 => 43,
    7863 => 43,
    7864 => 43,
    7865 => 43,
    7866 => 43,
    7867 => 43,
    7868 => 43,
    7869 => 43,
    7870 => 43,
    7871 => 43,
    7872 => 43,
    7873 => 43,
    7874 => 43,
    7875 => 43,
    7876 => 43,
    7877 => 43,
    7878 => 43,
    7879 => 43,
    7880 => 43,
    7881 => 43,
    7882 => 43,
    7883 => 43,
    7884 => 43,
    7885 => 43,
    7886 => 43,
    7887 => 43,
    7888 => 43,
    7889 => 43,
    7890 => 43,
    7891 => 43,
    7892 => 43,
    7893 => 43,
    7894 => 43,
    7895 => 43,
    7896 => 43,
    7897 => 43,
    7898 => 43,
    7899 => 43,
    7900 => 43,
    7901 => 43,
    7902 => 43,
    7903 => 43,
    7904 => 43,
    7905 => 43,
    7906 => 43,
    7907 => 43,
    7908 => 43,
    7909 => 43,
    7910 => 43,
    7911 => 43,
    7912 => 43,
    7913 => 43,
    7914 => 43,
    7915 => 43,
    7916 => 43,
    7917 => 43,
    7918 => 43,
    7919 => 43,
    7920 => 43,
    7921 => 43,
    7922 => 43,
    7923 => 43,
    7924 => 43,
    7925 => 43,
    7926 => 43,
    7927 => 43,
    7928 => 43,
    7929 => 43,
    7930 => 43,
    7931 => 43,
    7932 => 43,
    7933 => 43,
    7934 => 43,
    7935 => 43,
    7936 => 43,
    7937 => 43,
    7938 => 43,
    7939 => 43,
    7940 => 43,
    7941 => 43,
    7942 => 43,
    7943 => 43,
    7944 => 43,
    7945 => 43,
    7946 => 43,
    7947 => 43,
    7948 => 43,
    7949 => 43,
    7950 => 44,
    7951 => 44,
    7952 => 44,
    7953 => 44,
    7954 => 44,
    7955 => 44,
    7956 => 44,
    7957 => 44,
    7958 => 44,
    7959 => 44,
    7960 => 44,
    7961 => 44,
    7962 => 44,
    7963 => 44,
    7964 => 44,
    7965 => 44,
    7966 => 44,
    7967 => 44,
    7968 => 44,
    7969 => 44,
    7970 => 44,
    7971 => 44,
    7972 => 44,
    7973 => 44,
    7974 => 44,
    7975 => 44,
    7976 => 44,
    7977 => 44,
    7978 => 44,
    7979 => 44,
    7980 => 44,
    7981 => 44,
    7982 => 44,
    7983 => 44,
    7984 => 44,
    7985 => 44,
    7986 => 44,
    7987 => 44,
    7988 => 44,
    7989 => 44,
    7990 => 44,
    7991 => 44,
    7992 => 44,
    7993 => 44,
    7994 => 44,
    7995 => 44,
    7996 => 44,
    7997 => 44,
    7998 => 44,
    7999 => 44,
    8000 => 44,
    8001 => 44,
    8002 => 44,
    8003 => 44,
    8004 => 44,
    8005 => 44,
    8006 => 44,
    8007 => 44,
    8008 => 44,
    8009 => 44,
    8010 => 44,
    8011 => 44,
    8012 => 44,
    8013 => 44,
    8014 => 44,
    8015 => 44,
    8016 => 44,
    8017 => 44,
    8018 => 44,
    8019 => 44,
    8020 => 44,
    8021 => 44,
    8022 => 44,
    8023 => 44,
    8024 => 44,
    8025 => 44,
    8026 => 44,
    8027 => 44,
    8028 => 44,
    8029 => 44,
    8030 => 44,
    8031 => 44,
    8032 => 44,
    8033 => 44,
    8034 => 44,
    8035 => 44,
    8036 => 44,
    8037 => 44,
    8038 => 44,
    8039 => 44,
    8040 => 44,
    8041 => 44,
    8042 => 44,
    8043 => 44,
    8044 => 44,
    8045 => 44,
    8046 => 44,
    8047 => 44,
    8048 => 44,
    8049 => 44,
    8050 => 44,
    8051 => 44,
    8052 => 44,
    8053 => 44,
    8054 => 44,
    8055 => 44,
    8056 => 44,
    8057 => 44,
    8058 => 44,
    8059 => 44,
    8060 => 44,
    8061 => 44,
    8062 => 44,
    8063 => 44,
    8064 => 44,
    8065 => 44,
    8066 => 44,
    8067 => 44,
    8068 => 44,
    8069 => 44,
    8070 => 44,
    8071 => 44,
    8072 => 44,
    8073 => 44,
    8074 => 44,
    8075 => 44,
    8076 => 44,
    8077 => 44,
    8078 => 44,
    8079 => 44,
    8080 => 44,
    8081 => 44,
    8082 => 44,
    8083 => 44,
    8084 => 44,
    8085 => 44,
    8086 => 44,
    8087 => 44,
    8088 => 44,
    8089 => 44,
    8090 => 44,
    8091 => 44,
    8092 => 44,
    8093 => 44,
    8094 => 44,
    8095 => 44,
    8096 => 44,
    8097 => 44,
    8098 => 44,
    8099 => 44,
    8100 => 44,
    8101 => 44,
    8102 => 44,
    8103 => 44,
    8104 => 44,
    8105 => 44,
    8106 => 44,
    8107 => 44,
    8108 => 44,
    8109 => 44,
    8110 => 44,
    8111 => 44,
    8112 => 44,
    8113 => 44,
    8114 => 44,
    8115 => 44,
    8116 => 44,
    8117 => 44,
    8118 => 44,
    8119 => 44,
    8120 => 44,
    8121 => 44,
    8122 => 44,
    8123 => 44,
    8124 => 44,
    8125 => 44,
    8126 => 44,
    8127 => 44,
    8128 => 44,
    8129 => 44,
    8130 => 44,
    8131 => 44,
    8132 => 44,
    8133 => 44,
    8134 => 44,
    8135 => 44,
    8136 => 44,
    8137 => 44,
    8138 => 44,
    8139 => 44,
    8140 => 44,
    8141 => 44,
    8142 => 44,
    8143 => 44,
    8144 => 44,
    8145 => 44,
    8146 => 44,
    8147 => 44,
    8148 => 44,
    8149 => 44,
    8150 => 44,
    8151 => 44,
    8152 => 44,
    8153 => 44,
    8154 => 44,
    8155 => 44,
    8156 => 44,
    8157 => 44,
    8158 => 44,
    8159 => 44,
    8160 => 44,
    8161 => 44,
    8162 => 44,
    8163 => 44,
    8164 => 44,
    8165 => 44,
    8166 => 44,
    8167 => 44,
    8168 => 44,
    8169 => 44,
    8170 => 44,
    8171 => 44,
    8172 => 44,
    8173 => 44,
    8174 => 44,
    8175 => 44,
    8176 => 44,
    8177 => 44,
    8178 => 44,
    8179 => 44,
    8180 => 44,
    8181 => 45,
    8182 => 45,
    8183 => 45,
    8184 => 45,
    8185 => 45,
    8186 => 45,
    8187 => 45,
    8188 => 45,
    8189 => 45,
    8190 => 45,
    8191 => 45,
    8192 => 45,
    8193 => 45,
    8194 => 45,
    8195 => 45,
    8196 => 45,
    8197 => 45,
    8198 => 45,
    8199 => 45,
    8200 => 45,
    8201 => 45,
    8202 => 45,
    8203 => 45,
    8204 => 45,
    8205 => 45,
    8206 => 45,
    8207 => 45,
    8208 => 45,
    8209 => 45,
    8210 => 45,
    8211 => 45,
    8212 => 45,
    8213 => 45,
    8214 => 45,
    8215 => 45,
    8216 => 45,
    8217 => 45,
    8218 => 45,
    8219 => 45,
    8220 => 45,
    8221 => 45,
    8222 => 45,
    8223 => 45,
    8224 => 45,
    8225 => 45,
    8226 => 45,
    8227 => 45,
    8228 => 45,
    8229 => 45,
    8230 => 45,
    8231 => 45,
    8232 => 45,
    8233 => 45,
    8234 => 45,
    8235 => 45,
    8236 => 45,
    8237 => 45,
    8238 => 45,
    8239 => 45,
    8240 => 45,
    8241 => 45,
    8242 => 45,
    8243 => 45,
    8244 => 45,
    8245 => 45,
    8246 => 45,
    8247 => 45,
    8248 => 45,
    8249 => 45,
    8250 => 45,
    8251 => 45,
    8252 => 45,
    8253 => 45,
    8254 => 45,
    8255 => 45,
    8256 => 45,
    8257 => 45,
    8258 => 45,
    8259 => 45,
    8260 => 45,
    8261 => 45,
    8262 => 45,
    8263 => 45,
    8264 => 45,
    8265 => 45,
    8266 => 45,
    8267 => 45,
    8268 => 45,
    8269 => 45,
    8270 => 45,
    8271 => 45,
    8272 => 45,
    8273 => 45,
    8274 => 45,
    8275 => 45,
    8276 => 45,
    8277 => 45,
    8278 => 45,
    8279 => 45,
    8280 => 45,
    8281 => 45,
    8282 => 45,
    8283 => 45,
    8284 => 45,
    8285 => 45,
    8286 => 45,
    8287 => 45,
    8288 => 45,
    8289 => 45,
    8290 => 45,
    8291 => 45,
    8292 => 45,
    8293 => 45,
    8294 => 45,
    8295 => 45,
    8296 => 45,
    8297 => 45,
    8298 => 45,
    8299 => 45,
    8300 => 45,
    8301 => 45,
    8302 => 45,
    8303 => 45,
    8304 => 45,
    8305 => 45,
    8306 => 45,
    8307 => 45,
    8308 => 45,
    8309 => 45,
    8310 => 45,
    8311 => 45,
    8312 => 45,
    8313 => 45,
    8314 => 45,
    8315 => 45,
    8316 => 45,
    8317 => 45,
    8318 => 45,
    8319 => 45,
    8320 => 45,
    8321 => 45,
    8322 => 45,
    8323 => 45,
    8324 => 45,
    8325 => 45,
    8326 => 45,
    8327 => 45,
    8328 => 45,
    8329 => 45,
    8330 => 45,
    8331 => 45,
    8332 => 45,
    8333 => 45,
    8334 => 45,
    8335 => 45,
    8336 => 45,
    8337 => 45,
    8338 => 45,
    8339 => 45,
    8340 => 45,
    8341 => 45,
    8342 => 45,
    8343 => 45,
    8344 => 45,
    8345 => 45,
    8346 => 45,
    8347 => 45,
    8348 => 45,
    8349 => 45,
    8350 => 45,
    8351 => 45,
    8352 => 45,
    8353 => 45,
    8354 => 45,
    8355 => 45,
    8356 => 45,
    8357 => 45,
    8358 => 45,
    8359 => 45,
    8360 => 45,
    8361 => 45,
    8362 => 45,
    8363 => 45,
    8364 => 45,
    8365 => 45,
    8366 => 45,
    8367 => 45,
    8368 => 45,
    8369 => 45,
    8370 => 45,
    8371 => 45,
    8372 => 45,
    8373 => 45,
    8374 => 45,
    8375 => 45,
    8376 => 45,
    8377 => 45,
    8378 => 45,
    8379 => 45,
    8380 => 45,
    8381 => 45,
    8382 => 45,
    8383 => 45,
    8384 => 45,
    8385 => 45,
    8386 => 45,
    8387 => 45,
    8388 => 45,
    8389 => 45,
    8390 => 45,
    8391 => 45,
    8392 => 45,
    8393 => 45,
    8394 => 45,
    8395 => 45,
    8396 => 45,
    8397 => 45,
    8398 => 45,
    8399 => 45,
    8400 => 45,
    8401 => 45,
    8402 => 45,
    8403 => 45,
    8404 => 45,
    8405 => 45,
    8406 => 45,
    8407 => 45,
    8408 => 45,
    8409 => 45,
    8410 => 45,
    8411 => 45,
    8412 => 45,
    8413 => 45,
    8414 => 45,
    8415 => 45,
    8416 => 45,
    8417 => 45,
    8418 => 46,
    8419 => 46,
    8420 => 46,
    8421 => 46,
    8422 => 46,
    8423 => 46,
    8424 => 46,
    8425 => 46,
    8426 => 46,
    8427 => 46,
    8428 => 46,
    8429 => 46,
    8430 => 46,
    8431 => 46,
    8432 => 46,
    8433 => 46,
    8434 => 46,
    8435 => 46,
    8436 => 46,
    8437 => 46,
    8438 => 46,
    8439 => 46,
    8440 => 46,
    8441 => 46,
    8442 => 46,
    8443 => 46,
    8444 => 46,
    8445 => 46,
    8446 => 46,
    8447 => 46,
    8448 => 46,
    8449 => 46,
    8450 => 46,
    8451 => 46,
    8452 => 46,
    8453 => 46,
    8454 => 46,
    8455 => 46,
    8456 => 46,
    8457 => 46,
    8458 => 46,
    8459 => 46,
    8460 => 46,
    8461 => 46,
    8462 => 46,
    8463 => 46,
    8464 => 46,
    8465 => 46,
    8466 => 46,
    8467 => 46,
    8468 => 46,
    8469 => 46,
    8470 => 46,
    8471 => 46,
    8472 => 46,
    8473 => 46,
    8474 => 46,
    8475 => 46,
    8476 => 46,
    8477 => 46,
    8478 => 46,
    8479 => 46,
    8480 => 46,
    8481 => 46,
    8482 => 46,
    8483 => 46,
    8484 => 46,
    8485 => 46,
    8486 => 46,
    8487 => 46,
    8488 => 46,
    8489 => 46,
    8490 => 46,
    8491 => 46,
    8492 => 46,
    8493 => 46,
    8494 => 46,
    8495 => 46,
    8496 => 46,
    8497 => 46,
    8498 => 46,
    8499 => 46,
    8500 => 46,
    8501 => 46,
    8502 => 46,
    8503 => 46,
    8504 => 46,
    8505 => 46,
    8506 => 46,
    8507 => 46,
    8508 => 46,
    8509 => 46,
    8510 => 46,
    8511 => 46,
    8512 => 46,
    8513 => 46,
    8514 => 46,
    8515 => 46,
    8516 => 46,
    8517 => 46,
    8518 => 46,
    8519 => 46,
    8520 => 46,
    8521 => 46,
    8522 => 46,
    8523 => 46,
    8524 => 46,
    8525 => 46,
    8526 => 46,
    8527 => 46,
    8528 => 46,
    8529 => 46,
    8530 => 46,
    8531 => 46,
    8532 => 46,
    8533 => 46,
    8534 => 46,
    8535 => 46,
    8536 => 46,
    8537 => 46,
    8538 => 46,
    8539 => 46,
    8540 => 46,
    8541 => 46,
    8542 => 46,
    8543 => 46,
    8544 => 46,
    8545 => 46,
    8546 => 46,
    8547 => 46,
    8548 => 46,
    8549 => 46,
    8550 => 46,
    8551 => 46,
    8552 => 46,
    8553 => 46,
    8554 => 46,
    8555 => 46,
    8556 => 46,
    8557 => 46,
    8558 => 46,
    8559 => 46,
    8560 => 46,
    8561 => 46,
    8562 => 46,
    8563 => 46,
    8564 => 46,
    8565 => 46,
    8566 => 46,
    8567 => 46,
    8568 => 46,
    8569 => 46,
    8570 => 46,
    8571 => 46,
    8572 => 46,
    8573 => 46,
    8574 => 46,
    8575 => 46,
    8576 => 46,
    8577 => 46,
    8578 => 46,
    8579 => 46,
    8580 => 46,
    8581 => 46,
    8582 => 46,
    8583 => 46,
    8584 => 46,
    8585 => 46,
    8586 => 46,
    8587 => 46,
    8588 => 46,
    8589 => 46,
    8590 => 46,
    8591 => 46,
    8592 => 46,
    8593 => 46,
    8594 => 46,
    8595 => 46,
    8596 => 46,
    8597 => 46,
    8598 => 46,
    8599 => 46,
    8600 => 46,
    8601 => 46,
    8602 => 46,
    8603 => 46,
    8604 => 46,
    8605 => 46,
    8606 => 46,
    8607 => 46,
    8608 => 46,
    8609 => 46,
    8610 => 46,
    8611 => 46,
    8612 => 46,
    8613 => 46,
    8614 => 46,
    8615 => 46,
    8616 => 46,
    8617 => 46,
    8618 => 46,
    8619 => 46,
    8620 => 46,
    8621 => 46,
    8622 => 46,
    8623 => 46,
    8624 => 46,
    8625 => 46,
    8626 => 46,
    8627 => 46,
    8628 => 46,
    8629 => 46,
    8630 => 46,
    8631 => 46,
    8632 => 46,
    8633 => 46,
    8634 => 46,
    8635 => 46,
    8636 => 46,
    8637 => 46,
    8638 => 46,
    8639 => 46,
    8640 => 46,
    8641 => 46,
    8642 => 46,
    8643 => 46,
    8644 => 46,
    8645 => 46,
    8646 => 46,
    8647 => 46,
    8648 => 46,
    8649 => 46,
    8650 => 46,
    8651 => 46,
    8652 => 46,
    8653 => 46,
    8654 => 46,
    8655 => 46,
    8656 => 46,
    8657 => 46,
    8658 => 46,
    8659 => 46,
    8660 => 47,
    8661 => 47,
    8662 => 47,
    8663 => 47,
    8664 => 47,
    8665 => 47,
    8666 => 47,
    8667 => 47,
    8668 => 47,
    8669 => 47,
    8670 => 47,
    8671 => 47,
    8672 => 47,
    8673 => 47,
    8674 => 47,
    8675 => 47,
    8676 => 47,
    8677 => 47,
    8678 => 47,
    8679 => 47,
    8680 => 47,
    8681 => 47,
    8682 => 47,
    8683 => 47,
    8684 => 47,
    8685 => 47,
    8686 => 47,
    8687 => 47,
    8688 => 47,
    8689 => 47,
    8690 => 47,
    8691 => 47,
    8692 => 47,
    8693 => 47,
    8694 => 47,
    8695 => 47,
    8696 => 47,
    8697 => 47,
    8698 => 47,
    8699 => 47,
    8700 => 47,
    8701 => 47,
    8702 => 47,
    8703 => 47,
    8704 => 47,
    8705 => 47,
    8706 => 47,
    8707 => 47,
    8708 => 47,
    8709 => 47,
    8710 => 47,
    8711 => 47,
    8712 => 47,
    8713 => 47,
    8714 => 47,
    8715 => 47,
    8716 => 47,
    8717 => 47,
    8718 => 47,
    8719 => 47,
    8720 => 47,
    8721 => 47,
    8722 => 47,
    8723 => 47,
    8724 => 47,
    8725 => 47,
    8726 => 47,
    8727 => 47,
    8728 => 47,
    8729 => 47,
    8730 => 47,
    8731 => 47,
    8732 => 47,
    8733 => 47,
    8734 => 47,
    8735 => 47,
    8736 => 47,
    8737 => 47,
    8738 => 47,
    8739 => 47,
    8740 => 47,
    8741 => 47,
    8742 => 47,
    8743 => 47,
    8744 => 47,
    8745 => 47,
    8746 => 47,
    8747 => 47,
    8748 => 47,
    8749 => 47,
    8750 => 47,
    8751 => 47,
    8752 => 47,
    8753 => 47,
    8754 => 47,
    8755 => 47,
    8756 => 47,
    8757 => 47,
    8758 => 47,
    8759 => 47,
    8760 => 47,
    8761 => 47,
    8762 => 47,
    8763 => 47,
    8764 => 47,
    8765 => 47,
    8766 => 47,
    8767 => 47,
    8768 => 47,
    8769 => 47,
    8770 => 47,
    8771 => 47,
    8772 => 47,
    8773 => 47,
    8774 => 47,
    8775 => 47,
    8776 => 47,
    8777 => 47,
    8778 => 47,
    8779 => 47,
    8780 => 47,
    8781 => 47,
    8782 => 47,
    8783 => 47,
    8784 => 47,
    8785 => 47,
    8786 => 47,
    8787 => 47,
    8788 => 47,
    8789 => 47,
    8790 => 47,
    8791 => 47,
    8792 => 47,
    8793 => 47,
    8794 => 47,
    8795 => 47,
    8796 => 47,
    8797 => 47,
    8798 => 47,
    8799 => 47,
    8800 => 47,
    8801 => 47,
    8802 => 47,
    8803 => 47,
    8804 => 47,
    8805 => 47,
    8806 => 47,
    8807 => 47,
    8808 => 47,
    8809 => 47,
    8810 => 47,
    8811 => 47,
    8812 => 47,
    8813 => 47,
    8814 => 47,
    8815 => 47,
    8816 => 47,
    8817 => 47,
    8818 => 47,
    8819 => 47,
    8820 => 47,
    8821 => 47,
    8822 => 47,
    8823 => 47,
    8824 => 47,
    8825 => 47,
    8826 => 47,
    8827 => 47,
    8828 => 47,
    8829 => 47,
    8830 => 47,
    8831 => 47,
    8832 => 47,
    8833 => 47,
    8834 => 47,
    8835 => 47,
    8836 => 47,
    8837 => 47,
    8838 => 47,
    8839 => 47,
    8840 => 47,
    8841 => 47,
    8842 => 47,
    8843 => 47,
    8844 => 47,
    8845 => 47,
    8846 => 47,
    8847 => 47,
    8848 => 47,
    8849 => 47,
    8850 => 47,
    8851 => 47,
    8852 => 47,
    8853 => 47,
    8854 => 47,
    8855 => 47,
    8856 => 47,
    8857 => 47,
    8858 => 47,
    8859 => 47,
    8860 => 47,
    8861 => 47,
    8862 => 47,
    8863 => 47,
    8864 => 47,
    8865 => 47,
    8866 => 47,
    8867 => 47,
    8868 => 47,
    8869 => 47,
    8870 => 47,
    8871 => 47,
    8872 => 47,
    8873 => 47,
    8874 => 47,
    8875 => 47,
    8876 => 47,
    8877 => 47,
    8878 => 47,
    8879 => 47,
    8880 => 47,
    8881 => 47,
    8882 => 47,
    8883 => 47,
    8884 => 47,
    8885 => 47,
    8886 => 47,
    8887 => 47,
    8888 => 47,
    8889 => 47,
    8890 => 47,
    8891 => 47,
    8892 => 47,
    8893 => 47,
    8894 => 47,
    8895 => 47,
    8896 => 47,
    8897 => 47,
    8898 => 47,
    8899 => 47,
    8900 => 47,
    8901 => 47,
    8902 => 47,
    8903 => 47,
    8904 => 47,
    8905 => 47,
    8906 => 47,
    8907 => 47,
    8908 => 47,
    8909 => 48,
    8910 => 48,
    8911 => 48,
    8912 => 48,
    8913 => 48,
    8914 => 48,
    8915 => 48,
    8916 => 48,
    8917 => 48,
    8918 => 48,
    8919 => 48,
    8920 => 48,
    8921 => 48,
    8922 => 48,
    8923 => 48,
    8924 => 48,
    8925 => 48,
    8926 => 48,
    8927 => 48,
    8928 => 48,
    8929 => 48,
    8930 => 48,
    8931 => 48,
    8932 => 48,
    8933 => 48,
    8934 => 48,
    8935 => 48,
    8936 => 48,
    8937 => 48,
    8938 => 48,
    8939 => 48,
    8940 => 48,
    8941 => 48,
    8942 => 48,
    8943 => 48,
    8944 => 48,
    8945 => 48,
    8946 => 48,
    8947 => 48,
    8948 => 48,
    8949 => 48,
    8950 => 48,
    8951 => 48,
    8952 => 48,
    8953 => 48,
    8954 => 48,
    8955 => 48,
    8956 => 48,
    8957 => 48,
    8958 => 48,
    8959 => 48,
    8960 => 48,
    8961 => 48,
    8962 => 48,
    8963 => 48,
    8964 => 48,
    8965 => 48,
    8966 => 48,
    8967 => 48,
    8968 => 48,
    8969 => 48,
    8970 => 48,
    8971 => 48,
    8972 => 48,
    8973 => 48,
    8974 => 48,
    8975 => 48,
    8976 => 48,
    8977 => 48,
    8978 => 48,
    8979 => 48,
    8980 => 48,
    8981 => 48,
    8982 => 48,
    8983 => 48,
    8984 => 48,
    8985 => 48,
    8986 => 48,
    8987 => 48,
    8988 => 48,
    8989 => 48,
    8990 => 48,
    8991 => 48,
    8992 => 48,
    8993 => 48,
    8994 => 48,
    8995 => 48,
    8996 => 48,
    8997 => 48,
    8998 => 48,
    8999 => 48,
    9000 => 48,
    9001 => 48,
    9002 => 48,
    9003 => 48,
    9004 => 48,
    9005 => 48,
    9006 => 48,
    9007 => 48,
    9008 => 48,
    9009 => 48,
    9010 => 48,
    9011 => 48,
    9012 => 48,
    9013 => 48,
    9014 => 48,
    9015 => 48,
    9016 => 48,
    9017 => 48,
    9018 => 48,
    9019 => 48,
    9020 => 48,
    9021 => 48,
    9022 => 48,
    9023 => 48,
    9024 => 48,
    9025 => 48,
    9026 => 48,
    9027 => 48,
    9028 => 48,
    9029 => 48,
    9030 => 48,
    9031 => 48,
    9032 => 48,
    9033 => 48,
    9034 => 48,
    9035 => 48,
    9036 => 48,
    9037 => 48,
    9038 => 48,
    9039 => 48,
    9040 => 48,
    9041 => 48,
    9042 => 48,
    9043 => 48,
    9044 => 48,
    9045 => 48,
    9046 => 48,
    9047 => 48,
    9048 => 48,
    9049 => 48,
    9050 => 48,
    9051 => 48,
    9052 => 48,
    9053 => 48,
    9054 => 48,
    9055 => 48,
    9056 => 48,
    9057 => 48,
    9058 => 48,
    9059 => 48,
    9060 => 48,
    9061 => 48,
    9062 => 48,
    9063 => 48,
    9064 => 48,
    9065 => 48,
    9066 => 48,
    9067 => 48,
    9068 => 48,
    9069 => 48,
    9070 => 48,
    9071 => 48,
    9072 => 48,
    9073 => 48,
    9074 => 48,
    9075 => 48,
    9076 => 48,
    9077 => 48,
    9078 => 48,
    9079 => 48,
    9080 => 48,
    9081 => 48,
    9082 => 48,
    9083 => 48,
    9084 => 48,
    9085 => 48,
    9086 => 48,
    9087 => 48,
    9088 => 48,
    9089 => 48,
    9090 => 48,
    9091 => 48,
    9092 => 48,
    9093 => 48,
    9094 => 48,
    9095 => 48,
    9096 => 48,
    9097 => 48,
    9098 => 48,
    9099 => 48,
    9100 => 48,
    9101 => 48,
    9102 => 48,
    9103 => 48,
    9104 => 48,
    9105 => 48,
    9106 => 48,
    9107 => 48,
    9108 => 48,
    9109 => 48,
    9110 => 48,
    9111 => 48,
    9112 => 48,
    9113 => 48,
    9114 => 48,
    9115 => 48,
    9116 => 48,
    9117 => 48,
    9118 => 48,
    9119 => 48,
    9120 => 48,
    9121 => 48,
    9122 => 48,
    9123 => 48,
    9124 => 48,
    9125 => 48,
    9126 => 48,
    9127 => 48,
    9128 => 48,
    9129 => 48,
    9130 => 48,
    9131 => 48,
    9132 => 48,
    9133 => 48,
    9134 => 48,
    9135 => 48,
    9136 => 48,
    9137 => 48,
    9138 => 48,
    9139 => 48,
    9140 => 48,
    9141 => 48,
    9142 => 48,
    9143 => 48,
    9144 => 48,
    9145 => 48,
    9146 => 48,
    9147 => 48,
    9148 => 48,
    9149 => 48,
    9150 => 48,
    9151 => 48,
    9152 => 48,
    9153 => 48,
    9154 => 48,
    9155 => 48,
    9156 => 48,
    9157 => 48,
    9158 => 48,
    9159 => 48,
    9160 => 48,
    9161 => 48,
    9162 => 48,
    9163 => 48,
    9164 => 48,
    9165 => 49,
    9166 => 49,
    9167 => 49,
    9168 => 49,
    9169 => 49,
    9170 => 49,
    9171 => 49,
    9172 => 49,
    9173 => 49,
    9174 => 49,
    9175 => 49,
    9176 => 49,
    9177 => 49,
    9178 => 49,
    9179 => 49,
    9180 => 49,
    9181 => 49,
    9182 => 49,
    9183 => 49,
    9184 => 49,
    9185 => 49,
    9186 => 49,
    9187 => 49,
    9188 => 49,
    9189 => 49,
    9190 => 49,
    9191 => 49,
    9192 => 49,
    9193 => 49,
    9194 => 49,
    9195 => 49,
    9196 => 49,
    9197 => 49,
    9198 => 49,
    9199 => 49,
    9200 => 49,
    9201 => 49,
    9202 => 49,
    9203 => 49,
    9204 => 49,
    9205 => 49,
    9206 => 49,
    9207 => 49,
    9208 => 49,
    9209 => 49,
    9210 => 49,
    9211 => 49,
    9212 => 49,
    9213 => 49,
    9214 => 49,
    9215 => 49,
    9216 => 49,
    9217 => 49,
    9218 => 49,
    9219 => 49,
    9220 => 49,
    9221 => 49,
    9222 => 49,
    9223 => 49,
    9224 => 49,
    9225 => 49,
    9226 => 49,
    9227 => 49,
    9228 => 49,
    9229 => 49,
    9230 => 49,
    9231 => 49,
    9232 => 49,
    9233 => 49,
    9234 => 49,
    9235 => 49,
    9236 => 49,
    9237 => 49,
    9238 => 49,
    9239 => 49,
    9240 => 49,
    9241 => 49,
    9242 => 49,
    9243 => 49,
    9244 => 49,
    9245 => 49,
    9246 => 49,
    9247 => 49,
    9248 => 49,
    9249 => 49,
    9250 => 49,
    9251 => 49,
    9252 => 49,
    9253 => 49,
    9254 => 49,
    9255 => 49,
    9256 => 49,
    9257 => 49,
    9258 => 49,
    9259 => 49,
    9260 => 49,
    9261 => 49,
    9262 => 49,
    9263 => 49,
    9264 => 49,
    9265 => 49,
    9266 => 49,
    9267 => 49,
    9268 => 49,
    9269 => 49,
    9270 => 49,
    9271 => 49,
    9272 => 49,
    9273 => 49,
    9274 => 49,
    9275 => 49,
    9276 => 49,
    9277 => 49,
    9278 => 49,
    9279 => 49,
    9280 => 49,
    9281 => 49,
    9282 => 49,
    9283 => 49,
    9284 => 49,
    9285 => 49,
    9286 => 49,
    9287 => 49,
    9288 => 49,
    9289 => 49,
    9290 => 49,
    9291 => 49,
    9292 => 49,
    9293 => 49,
    9294 => 49,
    9295 => 49,
    9296 => 49,
    9297 => 49,
    9298 => 49,
    9299 => 49,
    9300 => 49,
    9301 => 49,
    9302 => 49,
    9303 => 49,
    9304 => 49,
    9305 => 49,
    9306 => 49,
    9307 => 49,
    9308 => 49,
    9309 => 49,
    9310 => 49,
    9311 => 49,
    9312 => 49,
    9313 => 49,
    9314 => 49,
    9315 => 49,
    9316 => 49,
    9317 => 49,
    9318 => 49,
    9319 => 49,
    9320 => 49,
    9321 => 49,
    9322 => 49,
    9323 => 49,
    9324 => 49,
    9325 => 49,
    9326 => 49,
    9327 => 49,
    9328 => 49,
    9329 => 49,
    9330 => 49,
    9331 => 49,
    9332 => 49,
    9333 => 49,
    9334 => 49,
    9335 => 49,
    9336 => 49,
    9337 => 49,
    9338 => 49,
    9339 => 49,
    9340 => 49,
    9341 => 49,
    9342 => 49,
    9343 => 49,
    9344 => 49,
    9345 => 49,
    9346 => 49,
    9347 => 49,
    9348 => 49,
    9349 => 49,
    9350 => 49,
    9351 => 49,
    9352 => 49,
    9353 => 49,
    9354 => 49,
    9355 => 49,
    9356 => 49,
    9357 => 49,
    9358 => 49,
    9359 => 49,
    9360 => 49,
    9361 => 49,
    9362 => 49,
    9363 => 49,
    9364 => 49,
    9365 => 49,
    9366 => 49,
    9367 => 49,
    9368 => 49,
    9369 => 49,
    9370 => 49,
    9371 => 49,
    9372 => 49,
    9373 => 49,
    9374 => 49,
    9375 => 49,
    9376 => 49,
    9377 => 49,
    9378 => 49,
    9379 => 49,
    9380 => 49,
    9381 => 49,
    9382 => 49,
    9383 => 49,
    9384 => 49,
    9385 => 49,
    9386 => 49,
    9387 => 49,
    9388 => 49,
    9389 => 49,
    9390 => 49,
    9391 => 49,
    9392 => 49,
    9393 => 49,
    9394 => 49,
    9395 => 49,
    9396 => 49,
    9397 => 49,
    9398 => 49,
    9399 => 49,
    9400 => 49,
    9401 => 49,
    9402 => 49,
    9403 => 49,
    9404 => 49,
    9405 => 49,
    9406 => 49,
    9407 => 49,
    9408 => 49,
    9409 => 49,
    9410 => 49,
    9411 => 49,
    9412 => 49,
    9413 => 49,
    9414 => 49,
    9415 => 49,
    9416 => 49,
    9417 => 49,
    9418 => 49,
    9419 => 49,
    9420 => 49,
    9421 => 49,
    9422 => 49,
    9423 => 49,
    9424 => 49,
    9425 => 49,
    9426 => 49,
    9427 => 49,
    9428 => 50,
    9429 => 50,
    9430 => 50,
    9431 => 50,
    9432 => 50,
    9433 => 50,
    9434 => 50,
    9435 => 50,
    9436 => 50,
    9437 => 50,
    9438 => 50,
    9439 => 50,
    9440 => 50,
    9441 => 50,
    9442 => 50,
    9443 => 50,
    9444 => 50,
    9445 => 50,
    9446 => 50,
    9447 => 50,
    9448 => 50,
    9449 => 50,
    9450 => 50,
    9451 => 50,
    9452 => 50,
    9453 => 50,
    9454 => 50,
    9455 => 50,
    9456 => 50,
    9457 => 50,
    9458 => 50,
    9459 => 50,
    9460 => 50,
    9461 => 50,
    9462 => 50,
    9463 => 50,
    9464 => 50,
    9465 => 50,
    9466 => 50,
    9467 => 50,
    9468 => 50,
    9469 => 50,
    9470 => 50,
    9471 => 50,
    9472 => 50,
    9473 => 50,
    9474 => 50,
    9475 => 50,
    9476 => 50,
    9477 => 50,
    9478 => 50,
    9479 => 50,
    9480 => 50,
    9481 => 50,
    9482 => 50,
    9483 => 50,
    9484 => 50,
    9485 => 50,
    9486 => 50,
    9487 => 50,
    9488 => 50,
    9489 => 50,
    9490 => 50,
    9491 => 50,
    9492 => 50,
    9493 => 50,
    9494 => 50,
    9495 => 50,
    9496 => 50,
    9497 => 50,
    9498 => 50,
    9499 => 50,
    9500 => 50,
    9501 => 50,
    9502 => 50,
    9503 => 50,
    9504 => 50,
    9505 => 50,
    9506 => 50,
    9507 => 50,
    9508 => 50,
    9509 => 50,
    9510 => 50,
    9511 => 50,
    9512 => 50,
    9513 => 50,
    9514 => 50,
    9515 => 50,
    9516 => 50,
    9517 => 50,
    9518 => 50,
    9519 => 50,
    9520 => 50,
    9521 => 50,
    9522 => 50,
    9523 => 50,
    9524 => 50,
    9525 => 50,
    9526 => 50,
    9527 => 50,
    9528 => 50,
    9529 => 50,
    9530 => 50,
    9531 => 50,
    9532 => 50,
    9533 => 50,
    9534 => 50,
    9535 => 50,
    9536 => 50,
    9537 => 50,
    9538 => 50,
    9539 => 50,
    9540 => 50,
    9541 => 50,
    9542 => 50,
    9543 => 50,
    9544 => 50,
    9545 => 50,
    9546 => 50,
    9547 => 50,
    9548 => 50,
    9549 => 50,
    9550 => 50,
    9551 => 50,
    9552 => 50,
    9553 => 50,
    9554 => 50,
    9555 => 50,
    9556 => 50,
    9557 => 50,
    9558 => 50,
    9559 => 50,
    9560 => 50,
    9561 => 50,
    9562 => 50,
    9563 => 50,
    9564 => 50,
    9565 => 50,
    9566 => 50,
    9567 => 50,
    9568 => 50,
    9569 => 50,
    9570 => 50,
    9571 => 50,
    9572 => 50,
    9573 => 50,
    9574 => 50,
    9575 => 50,
    9576 => 50,
    9577 => 50,
    9578 => 50,
    9579 => 50,
    9580 => 50,
    9581 => 50,
    9582 => 50,
    9583 => 50,
    9584 => 50,
    9585 => 50,
    9586 => 50,
    9587 => 50,
    9588 => 50,
    9589 => 50,
    9590 => 50,
    9591 => 50,
    9592 => 50,
    9593 => 50,
    9594 => 50,
    9595 => 50,
    9596 => 50,
    9597 => 50,
    9598 => 50,
    9599 => 50,
    9600 => 50,
    9601 => 50,
    9602 => 50,
    9603 => 50,
    9604 => 50,
    9605 => 50,
    9606 => 50,
    9607 => 50,
    9608 => 50,
    9609 => 50,
    9610 => 50,
    9611 => 50,
    9612 => 50,
    9613 => 50,
    9614 => 50,
    9615 => 50,
    9616 => 50,
    9617 => 50,
    9618 => 50,
    9619 => 50,
    9620 => 50,
    9621 => 50,
    9622 => 50,
    9623 => 50,
    9624 => 50,
    9625 => 50,
    9626 => 50,
    9627 => 50,
    9628 => 50,
    9629 => 50,
    9630 => 50,
    9631 => 50,
    9632 => 50,
    9633 => 50,
    9634 => 50,
    9635 => 50,
    9636 => 50,
    9637 => 50,
    9638 => 50,
    9639 => 50,
    9640 => 50,
    9641 => 50,
    9642 => 50,
    9643 => 50,
    9644 => 50,
    9645 => 50,
    9646 => 50,
    9647 => 50,
    9648 => 50,
    9649 => 50,
    9650 => 50,
    9651 => 50,
    9652 => 50,
    9653 => 50,
    9654 => 50,
    9655 => 50,
    9656 => 50,
    9657 => 50,
    9658 => 50,
    9659 => 50,
    9660 => 50,
    9661 => 50,
    9662 => 50,
    9663 => 50,
    9664 => 50,
    9665 => 50,
    9666 => 50,
    9667 => 50,
    9668 => 50,
    9669 => 50,
    9670 => 50,
    9671 => 50,
    9672 => 50,
    9673 => 50,
    9674 => 50,
    9675 => 50,
    9676 => 50,
    9677 => 50,
    9678 => 50,
    9679 => 50,
    9680 => 50,
    9681 => 50,
    9682 => 50,
    9683 => 50,
    9684 => 50,
    9685 => 50,
    9686 => 50,
    9687 => 50,
    9688 => 50,
    9689 => 50,
    9690 => 50,
    9691 => 50,
    9692 => 50,
    9693 => 50,
    9694 => 50,
    9695 => 50,
    9696 => 50,
    9697 => 50,
    9698 => 50,
    9699 => 50,
    9700 => 51,
    9701 => 51,
    9702 => 51,
    9703 => 51,
    9704 => 51,
    9705 => 51,
    9706 => 51,
    9707 => 51,
    9708 => 51,
    9709 => 51,
    9710 => 51,
    9711 => 51,
    9712 => 51,
    9713 => 51,
    9714 => 51,
    9715 => 51,
    9716 => 51,
    9717 => 51,
    9718 => 51,
    9719 => 51,
    9720 => 51,
    9721 => 51,
    9722 => 51,
    9723 => 51,
    9724 => 51,
    9725 => 51,
    9726 => 51,
    9727 => 51,
    9728 => 51,
    9729 => 51,
    9730 => 51,
    9731 => 51,
    9732 => 51,
    9733 => 51,
    9734 => 51,
    9735 => 51,
    9736 => 51,
    9737 => 51,
    9738 => 51,
    9739 => 51,
    9740 => 51,
    9741 => 51,
    9742 => 51,
    9743 => 51,
    9744 => 51,
    9745 => 51,
    9746 => 51,
    9747 => 51,
    9748 => 51,
    9749 => 51,
    9750 => 51,
    9751 => 51,
    9752 => 51,
    9753 => 51,
    9754 => 51,
    9755 => 51,
    9756 => 51,
    9757 => 51,
    9758 => 51,
    9759 => 51,
    9760 => 51,
    9761 => 51,
    9762 => 51,
    9763 => 51,
    9764 => 51,
    9765 => 51,
    9766 => 51,
    9767 => 51,
    9768 => 51,
    9769 => 51,
    9770 => 51,
    9771 => 51,
    9772 => 51,
    9773 => 51,
    9774 => 51,
    9775 => 51,
    9776 => 51,
    9777 => 51,
    9778 => 51,
    9779 => 51,
    9780 => 51,
    9781 => 51,
    9782 => 51,
    9783 => 51,
    9784 => 51,
    9785 => 51,
    9786 => 51,
    9787 => 51,
    9788 => 51,
    9789 => 51,
    9790 => 51,
    9791 => 51,
    9792 => 51,
    9793 => 51,
    9794 => 51,
    9795 => 51,
    9796 => 51,
    9797 => 51,
    9798 => 51,
    9799 => 51,
    9800 => 51,
    9801 => 51,
    9802 => 51,
    9803 => 51,
    9804 => 51,
    9805 => 51,
    9806 => 51,
    9807 => 51,
    9808 => 51,
    9809 => 51,
    9810 => 51,
    9811 => 51,
    9812 => 51,
    9813 => 51,
    9814 => 51,
    9815 => 51,
    9816 => 51,
    9817 => 51,
    9818 => 51,
    9819 => 51,
    9820 => 51,
    9821 => 51,
    9822 => 51,
    9823 => 51,
    9824 => 51,
    9825 => 51,
    9826 => 51,
    9827 => 51,
    9828 => 51,
    9829 => 51,
    9830 => 51,
    9831 => 51,
    9832 => 51,
    9833 => 51,
    9834 => 51,
    9835 => 51,
    9836 => 51,
    9837 => 51,
    9838 => 51,
    9839 => 51,
    9840 => 51,
    9841 => 51,
    9842 => 51,
    9843 => 51,
    9844 => 51,
    9845 => 51,
    9846 => 51,
    9847 => 51,
    9848 => 51,
    9849 => 51,
    9850 => 51,
    9851 => 51,
    9852 => 51,
    9853 => 51,
    9854 => 51,
    9855 => 51,
    9856 => 51,
    9857 => 51,
    9858 => 51,
    9859 => 51,
    9860 => 51,
    9861 => 51,
    9862 => 51,
    9863 => 51,
    9864 => 51,
    9865 => 51,
    9866 => 51,
    9867 => 51,
    9868 => 51,
    9869 => 51,
    9870 => 51,
    9871 => 51,
    9872 => 51,
    9873 => 51,
    9874 => 51,
    9875 => 51,
    9876 => 51,
    9877 => 51,
    9878 => 51,
    9879 => 51,
    9880 => 51,
    9881 => 51,
    9882 => 51,
    9883 => 51,
    9884 => 51,
    9885 => 51,
    9886 => 51,
    9887 => 51,
    9888 => 51,
    9889 => 51,
    9890 => 51,
    9891 => 51,
    9892 => 51,
    9893 => 51,
    9894 => 51,
    9895 => 51,
    9896 => 51,
    9897 => 51,
    9898 => 51,
    9899 => 51,
    9900 => 51,
    9901 => 51,
    9902 => 51,
    9903 => 51,
    9904 => 51,
    9905 => 51,
    9906 => 51,
    9907 => 51,
    9908 => 51,
    9909 => 51,
    9910 => 51,
    9911 => 51,
    9912 => 51,
    9913 => 51,
    9914 => 51,
    9915 => 51,
    9916 => 51,
    9917 => 51,
    9918 => 51,
    9919 => 51,
    9920 => 51,
    9921 => 51,
    9922 => 51,
    9923 => 51,
    9924 => 51,
    9925 => 51,
    9926 => 51,
    9927 => 51,
    9928 => 51,
    9929 => 51,
    9930 => 51,
    9931 => 51,
    9932 => 51,
    9933 => 51,
    9934 => 51,
    9935 => 51,
    9936 => 51,
    9937 => 51,
    9938 => 51,
    9939 => 51,
    9940 => 51,
    9941 => 51,
    9942 => 51,
    9943 => 51,
    9944 => 51,
    9945 => 51,
    9946 => 51,
    9947 => 51,
    9948 => 51,
    9949 => 51,
    9950 => 51,
    9951 => 51,
    9952 => 51,
    9953 => 51,
    9954 => 51,
    9955 => 51,
    9956 => 51,
    9957 => 51,
    9958 => 51,
    9959 => 51,
    9960 => 51,
    9961 => 51,
    9962 => 51,
    9963 => 51,
    9964 => 51,
    9965 => 51,
    9966 => 51,
    9967 => 51,
    9968 => 51,
    9969 => 51,
    9970 => 51,
    9971 => 51,
    9972 => 51,
    9973 => 51,
    9974 => 51,
    9975 => 51,
    9976 => 51,
    9977 => 51,
    9978 => 51,
    9979 => 51,
    9980 => 51,
    9981 => 51,
    9982 => 52,
    9983 => 52,
    9984 => 52,
    9985 => 52,
    9986 => 52,
    9987 => 52,
    9988 => 52,
    9989 => 52,
    9990 => 52,
    9991 => 52,
    9992 => 52,
    9993 => 52,
    9994 => 52,
    9995 => 52,
    9996 => 52,
    9997 => 52,
    9998 => 52,
    9999 => 52,
    10000 => 52,
    10001 => 52,
    10002 => 52,
    10003 => 52,
    10004 => 52,
    10005 => 52,
    10006 => 52,
    10007 => 52,
    10008 => 52,
    10009 => 52,
    10010 => 52,
    10011 => 52,
    10012 => 52,
    10013 => 52,
    10014 => 52,
    10015 => 52,
    10016 => 52,
    10017 => 52,
    10018 => 52,
    10019 => 52,
    10020 => 52,
    10021 => 52,
    10022 => 52,
    10023 => 52,
    10024 => 52,
    10025 => 52,
    10026 => 52,
    10027 => 52,
    10028 => 52,
    10029 => 52,
    10030 => 52,
    10031 => 52,
    10032 => 52,
    10033 => 52,
    10034 => 52,
    10035 => 52,
    10036 => 52,
    10037 => 52,
    10038 => 52,
    10039 => 52,
    10040 => 52,
    10041 => 52,
    10042 => 52,
    10043 => 52,
    10044 => 52,
    10045 => 52,
    10046 => 52,
    10047 => 52,
    10048 => 52,
    10049 => 52,
    10050 => 52,
    10051 => 52,
    10052 => 52,
    10053 => 52,
    10054 => 52,
    10055 => 52,
    10056 => 52,
    10057 => 52,
    10058 => 52,
    10059 => 52,
    10060 => 52,
    10061 => 52,
    10062 => 52,
    10063 => 52,
    10064 => 52,
    10065 => 52,
    10066 => 52,
    10067 => 52,
    10068 => 52,
    10069 => 52,
    10070 => 52,
    10071 => 52,
    10072 => 52,
    10073 => 52,
    10074 => 52,
    10075 => 52,
    10076 => 52,
    10077 => 52,
    10078 => 52,
    10079 => 52,
    10080 => 52,
    10081 => 52,
    10082 => 52,
    10083 => 52,
    10084 => 52,
    10085 => 52,
    10086 => 52,
    10087 => 52,
    10088 => 52,
    10089 => 52,
    10090 => 52,
    10091 => 52,
    10092 => 52,
    10093 => 52,
    10094 => 52,
    10095 => 52,
    10096 => 52,
    10097 => 52,
    10098 => 52,
    10099 => 52,
    10100 => 52,
    10101 => 52,
    10102 => 52,
    10103 => 52,
    10104 => 52,
    10105 => 52,
    10106 => 52,
    10107 => 52,
    10108 => 52,
    10109 => 52,
    10110 => 52,
    10111 => 52,
    10112 => 52,
    10113 => 52,
    10114 => 52,
    10115 => 52,
    10116 => 52,
    10117 => 52,
    10118 => 52,
    10119 => 52,
    10120 => 52,
    10121 => 52,
    10122 => 52,
    10123 => 52,
    10124 => 52,
    10125 => 52,
    10126 => 52,
    10127 => 52,
    10128 => 52,
    10129 => 52,
    10130 => 52,
    10131 => 52,
    10132 => 52,
    10133 => 52,
    10134 => 52,
    10135 => 52,
    10136 => 52,
    10137 => 52,
    10138 => 52,
    10139 => 52,
    10140 => 52,
    10141 => 52,
    10142 => 52,
    10143 => 52,
    10144 => 52,
    10145 => 52,
    10146 => 52,
    10147 => 52,
    10148 => 52,
    10149 => 52,
    10150 => 52,
    10151 => 52,
    10152 => 52,
    10153 => 52,
    10154 => 52,
    10155 => 52,
    10156 => 52,
    10157 => 52,
    10158 => 52,
    10159 => 52,
    10160 => 52,
    10161 => 52,
    10162 => 52,
    10163 => 52,
    10164 => 52,
    10165 => 52,
    10166 => 52,
    10167 => 52,
    10168 => 52,
    10169 => 52,
    10170 => 52,
    10171 => 52,
    10172 => 52,
    10173 => 52,
    10174 => 52,
    10175 => 52,
    10176 => 52,
    10177 => 52,
    10178 => 52,
    10179 => 52,
    10180 => 52,
    10181 => 52,
    10182 => 52,
    10183 => 52,
    10184 => 52,
    10185 => 52,
    10186 => 52,
    10187 => 52,
    10188 => 52,
    10189 => 52,
    10190 => 52,
    10191 => 52,
    10192 => 52,
    10193 => 52,
    10194 => 52,
    10195 => 52,
    10196 => 52,
    10197 => 52,
    10198 => 52,
    10199 => 52,
    10200 => 52,
    10201 => 52,
    10202 => 52,
    10203 => 52,
    10204 => 52,
    10205 => 52,
    10206 => 52,
    10207 => 52,
    10208 => 52,
    10209 => 52,
    10210 => 52,
    10211 => 52,
    10212 => 52,
    10213 => 52,
    10214 => 52,
    10215 => 52,
    10216 => 52,
    10217 => 52,
    10218 => 52,
    10219 => 52,
    10220 => 52,
    10221 => 52,
    10222 => 52,
    10223 => 52,
    10224 => 52,
    10225 => 52,
    10226 => 52,
    10227 => 52,
    10228 => 52,
    10229 => 52,
    10230 => 52,
    10231 => 52,
    10232 => 52,
    10233 => 52,
    10234 => 52,
    10235 => 52,
    10236 => 52,
    10237 => 52,
    10238 => 52,
    10239 => 52,
    10240 => 52,
    10241 => 52,
    10242 => 52,
    10243 => 52,
    10244 => 52,
    10245 => 52,
    10246 => 52,
    10247 => 52,
    10248 => 52,
    10249 => 52,
    10250 => 52,
    10251 => 52,
    10252 => 52,
    10253 => 52,
    10254 => 52,
    10255 => 52,
    10256 => 52,
    10257 => 52,
    10258 => 52,
    10259 => 52,
    10260 => 52,
    10261 => 52,
    10262 => 52,
    10263 => 52,
    10264 => 52,
    10265 => 52,
    10266 => 52,
    10267 => 52,
    10268 => 52,
    10269 => 52,
    10270 => 52,
    10271 => 52,
    10272 => 52,
    10273 => 52,
    10274 => 52,
    10275 => 52,
    10276 => 53,
    10277 => 53,
    10278 => 53,
    10279 => 53,
    10280 => 53,
    10281 => 53,
    10282 => 53,
    10283 => 53,
    10284 => 53,
    10285 => 53,
    10286 => 53,
    10287 => 53,
    10288 => 53,
    10289 => 53,
    10290 => 53,
    10291 => 53,
    10292 => 53,
    10293 => 53,
    10294 => 53,
    10295 => 53,
    10296 => 53,
    10297 => 53,
    10298 => 53,
    10299 => 53,
    10300 => 53,
    10301 => 53,
    10302 => 53,
    10303 => 53,
    10304 => 53,
    10305 => 53,
    10306 => 53,
    10307 => 53,
    10308 => 53,
    10309 => 53,
    10310 => 53,
    10311 => 53,
    10312 => 53,
    10313 => 53,
    10314 => 53,
    10315 => 53,
    10316 => 53,
    10317 => 53,
    10318 => 53,
    10319 => 53,
    10320 => 53,
    10321 => 53,
    10322 => 53,
    10323 => 53,
    10324 => 53,
    10325 => 53,
    10326 => 53,
    10327 => 53,
    10328 => 53,
    10329 => 53,
    10330 => 53,
    10331 => 53,
    10332 => 53,
    10333 => 53,
    10334 => 53,
    10335 => 53,
    10336 => 53,
    10337 => 53,
    10338 => 53,
    10339 => 53,
    10340 => 53,
    10341 => 53,
    10342 => 53,
    10343 => 53,
    10344 => 53,
    10345 => 53,
    10346 => 53,
    10347 => 53,
    10348 => 53,
    10349 => 53,
    10350 => 53,
    10351 => 53,
    10352 => 53,
    10353 => 53,
    10354 => 53,
    10355 => 53,
    10356 => 53,
    10357 => 53,
    10358 => 53,
    10359 => 53,
    10360 => 53,
    10361 => 53,
    10362 => 53,
    10363 => 53,
    10364 => 53,
    10365 => 53,
    10366 => 53,
    10367 => 53,
    10368 => 53,
    10369 => 53,
    10370 => 53,
    10371 => 53,
    10372 => 53,
    10373 => 53,
    10374 => 53,
    10375 => 53,
    10376 => 53,
    10377 => 53,
    10378 => 53,
    10379 => 53,
    10380 => 53,
    10381 => 53,
    10382 => 53,
    10383 => 53,
    10384 => 53,
    10385 => 53,
    10386 => 53,
    10387 => 53,
    10388 => 53,
    10389 => 53,
    10390 => 53,
    10391 => 53,
    10392 => 53,
    10393 => 53,
    10394 => 53,
    10395 => 53,
    10396 => 53,
    10397 => 53,
    10398 => 53,
    10399 => 53,
    10400 => 53,
    10401 => 53,
    10402 => 53,
    10403 => 53,
    10404 => 53,
    10405 => 53,
    10406 => 53,
    10407 => 53,
    10408 => 53,
    10409 => 53,
    10410 => 53,
    10411 => 53,
    10412 => 53,
    10413 => 53,
    10414 => 53,
    10415 => 53,
    10416 => 53,
    10417 => 53,
    10418 => 53,
    10419 => 53,
    10420 => 53,
    10421 => 53,
    10422 => 53,
    10423 => 53,
    10424 => 53,
    10425 => 53,
    10426 => 53,
    10427 => 53,
    10428 => 53,
    10429 => 53,
    10430 => 53,
    10431 => 53,
    10432 => 53,
    10433 => 53,
    10434 => 53,
    10435 => 53,
    10436 => 53,
    10437 => 53,
    10438 => 53,
    10439 => 53,
    10440 => 53,
    10441 => 53,
    10442 => 53,
    10443 => 53,
    10444 => 53,
    10445 => 53,
    10446 => 53,
    10447 => 53,
    10448 => 53,
    10449 => 53,
    10450 => 53,
    10451 => 53,
    10452 => 53,
    10453 => 53,
    10454 => 53,
    10455 => 53,
    10456 => 53,
    10457 => 53,
    10458 => 53,
    10459 => 53,
    10460 => 53,
    10461 => 53,
    10462 => 53,
    10463 => 53,
    10464 => 53,
    10465 => 53,
    10466 => 53,
    10467 => 53,
    10468 => 53,
    10469 => 53,
    10470 => 53,
    10471 => 53,
    10472 => 53,
    10473 => 53,
    10474 => 53,
    10475 => 53,
    10476 => 53,
    10477 => 53,
    10478 => 53,
    10479 => 53,
    10480 => 53,
    10481 => 53,
    10482 => 53,
    10483 => 53,
    10484 => 53,
    10485 => 53,
    10486 => 53,
    10487 => 53,
    10488 => 53,
    10489 => 53,
    10490 => 53,
    10491 => 53,
    10492 => 53,
    10493 => 53,
    10494 => 53,
    10495 => 53,
    10496 => 53,
    10497 => 53,
    10498 => 53,
    10499 => 53,
    10500 => 53,
    10501 => 53,
    10502 => 53,
    10503 => 53,
    10504 => 53,
    10505 => 53,
    10506 => 53,
    10507 => 53,
    10508 => 53,
    10509 => 53,
    10510 => 53,
    10511 => 53,
    10512 => 53,
    10513 => 53,
    10514 => 53,
    10515 => 53,
    10516 => 53,
    10517 => 53,
    10518 => 53,
    10519 => 53,
    10520 => 53,
    10521 => 53,
    10522 => 53,
    10523 => 53,
    10524 => 53,
    10525 => 53,
    10526 => 53,
    10527 => 53,
    10528 => 53,
    10529 => 53,
    10530 => 53,
    10531 => 53,
    10532 => 53,
    10533 => 53,
    10534 => 53,
    10535 => 53,
    10536 => 53,
    10537 => 53,
    10538 => 53,
    10539 => 53,
    10540 => 53,
    10541 => 53,
    10542 => 53,
    10543 => 53,
    10544 => 53,
    10545 => 53,
    10546 => 53,
    10547 => 53,
    10548 => 53,
    10549 => 53,
    10550 => 53,
    10551 => 53,
    10552 => 53,
    10553 => 53,
    10554 => 53,
    10555 => 53,
    10556 => 53,
    10557 => 53,
    10558 => 53,
    10559 => 53,
    10560 => 53,
    10561 => 53,
    10562 => 53,
    10563 => 53,
    10564 => 53,
    10565 => 53,
    10566 => 53,
    10567 => 53,
    10568 => 53,
    10569 => 53,
    10570 => 53,
    10571 => 53,
    10572 => 53,
    10573 => 53,
    10574 => 53,
    10575 => 53,
    10576 => 53,
    10577 => 53,
    10578 => 53,
    10579 => 53,
    10580 => 53,
    10581 => 53,
    10582 => 54,
    10583 => 54,
    10584 => 54,
    10585 => 54,
    10586 => 54,
    10587 => 54,
    10588 => 54,
    10589 => 54,
    10590 => 54,
    10591 => 54,
    10592 => 54,
    10593 => 54,
    10594 => 54,
    10595 => 54,
    10596 => 54,
    10597 => 54,
    10598 => 54,
    10599 => 54,
    10600 => 54,
    10601 => 54,
    10602 => 54,
    10603 => 54,
    10604 => 54,
    10605 => 54,
    10606 => 54,
    10607 => 54,
    10608 => 54,
    10609 => 54,
    10610 => 54,
    10611 => 54,
    10612 => 54,
    10613 => 54,
    10614 => 54,
    10615 => 54,
    10616 => 54,
    10617 => 54,
    10618 => 54,
    10619 => 54,
    10620 => 54,
    10621 => 54,
    10622 => 54,
    10623 => 54,
    10624 => 54,
    10625 => 54,
    10626 => 54,
    10627 => 54,
    10628 => 54,
    10629 => 54,
    10630 => 54,
    10631 => 54,
    10632 => 54,
    10633 => 54,
    10634 => 54,
    10635 => 54,
    10636 => 54,
    10637 => 54,
    10638 => 54,
    10639 => 54,
    10640 => 54,
    10641 => 54,
    10642 => 54,
    10643 => 54,
    10644 => 54,
    10645 => 54,
    10646 => 54,
    10647 => 54,
    10648 => 54,
    10649 => 54,
    10650 => 54,
    10651 => 54,
    10652 => 54,
    10653 => 54,
    10654 => 54,
    10655 => 54,
    10656 => 54,
    10657 => 54,
    10658 => 54,
    10659 => 54,
    10660 => 54,
    10661 => 54,
    10662 => 54,
    10663 => 54,
    10664 => 54,
    10665 => 54,
    10666 => 54,
    10667 => 54,
    10668 => 54,
    10669 => 54,
    10670 => 54,
    10671 => 54,
    10672 => 54,
    10673 => 54,
    10674 => 54,
    10675 => 54,
    10676 => 54,
    10677 => 54,
    10678 => 54,
    10679 => 54,
    10680 => 54,
    10681 => 54,
    10682 => 54,
    10683 => 54,
    10684 => 54,
    10685 => 54,
    10686 => 54,
    10687 => 54,
    10688 => 54,
    10689 => 54,
    10690 => 54,
    10691 => 54,
    10692 => 54,
    10693 => 54,
    10694 => 54,
    10695 => 54,
    10696 => 54,
    10697 => 54,
    10698 => 54,
    10699 => 54,
    10700 => 54,
    10701 => 54,
    10702 => 54,
    10703 => 54,
    10704 => 54,
    10705 => 54,
    10706 => 54,
    10707 => 54,
    10708 => 54,
    10709 => 54,
    10710 => 54,
    10711 => 54,
    10712 => 54,
    10713 => 54,
    10714 => 54,
    10715 => 54,
    10716 => 54,
    10717 => 54,
    10718 => 54,
    10719 => 54,
    10720 => 54,
    10721 => 54,
    10722 => 54,
    10723 => 54,
    10724 => 54,
    10725 => 54,
    10726 => 54,
    10727 => 54,
    10728 => 54,
    10729 => 54,
    10730 => 54,
    10731 => 54,
    10732 => 54,
    10733 => 54,
    10734 => 54,
    10735 => 54,
    10736 => 54,
    10737 => 54,
    10738 => 54,
    10739 => 54,
    10740 => 54,
    10741 => 54,
    10742 => 54,
    10743 => 54,
    10744 => 54,
    10745 => 54,
    10746 => 54,
    10747 => 54,
    10748 => 54,
    10749 => 54,
    10750 => 54,
    10751 => 54,
    10752 => 54,
    10753 => 54,
    10754 => 54,
    10755 => 54,
    10756 => 54,
    10757 => 54,
    10758 => 54,
    10759 => 54,
    10760 => 54,
    10761 => 54,
    10762 => 54,
    10763 => 54,
    10764 => 54,
    10765 => 54,
    10766 => 54,
    10767 => 54,
    10768 => 54,
    10769 => 54,
    10770 => 54,
    10771 => 54,
    10772 => 54,
    10773 => 54,
    10774 => 54,
    10775 => 54,
    10776 => 54,
    10777 => 54,
    10778 => 54,
    10779 => 54,
    10780 => 54,
    10781 => 54,
    10782 => 54,
    10783 => 54,
    10784 => 54,
    10785 => 54,
    10786 => 54,
    10787 => 54,
    10788 => 54,
    10789 => 54,
    10790 => 54,
    10791 => 54,
    10792 => 54,
    10793 => 54,
    10794 => 54,
    10795 => 54,
    10796 => 54,
    10797 => 54,
    10798 => 54,
    10799 => 54,
    10800 => 54,
    10801 => 54,
    10802 => 54,
    10803 => 54,
    10804 => 54,
    10805 => 54,
    10806 => 54,
    10807 => 54,
    10808 => 54,
    10809 => 54,
    10810 => 54,
    10811 => 54,
    10812 => 54,
    10813 => 54,
    10814 => 54,
    10815 => 54,
    10816 => 54,
    10817 => 54,
    10818 => 54,
    10819 => 54,
    10820 => 54,
    10821 => 54,
    10822 => 54,
    10823 => 54,
    10824 => 54,
    10825 => 54,
    10826 => 54,
    10827 => 54,
    10828 => 54,
    10829 => 54,
    10830 => 54,
    10831 => 54,
    10832 => 54,
    10833 => 54,
    10834 => 54,
    10835 => 54,
    10836 => 54,
    10837 => 54,
    10838 => 54,
    10839 => 54,
    10840 => 54,
    10841 => 54,
    10842 => 54,
    10843 => 54,
    10844 => 54,
    10845 => 54,
    10846 => 54,
    10847 => 54,
    10848 => 54,
    10849 => 54,
    10850 => 54,
    10851 => 54,
    10852 => 54,
    10853 => 54,
    10854 => 54,
    10855 => 54,
    10856 => 54,
    10857 => 54,
    10858 => 54,
    10859 => 54,
    10860 => 54,
    10861 => 54,
    10862 => 54,
    10863 => 54,
    10864 => 54,
    10865 => 54,
    10866 => 54,
    10867 => 54,
    10868 => 54,
    10869 => 54,
    10870 => 54,
    10871 => 54,
    10872 => 54,
    10873 => 54,
    10874 => 54,
    10875 => 54,
    10876 => 54,
    10877 => 54,
    10878 => 54,
    10879 => 54,
    10880 => 54,
    10881 => 54,
    10882 => 54,
    10883 => 54,
    10884 => 54,
    10885 => 54,
    10886 => 54,
    10887 => 54,
    10888 => 54,
    10889 => 54,
    10890 => 54,
    10891 => 54,
    10892 => 54,
    10893 => 54,
    10894 => 54,
    10895 => 54,
    10896 => 54,
    10897 => 54,
    10898 => 54,
    10899 => 54,
    10900 => 54,
    10901 => 54,
    10902 => 54,
    10903 => 55,
    10904 => 55,
    10905 => 55,
    10906 => 55,
    10907 => 55,
    10908 => 55,
    10909 => 55,
    10910 => 55,
    10911 => 55,
    10912 => 55,
    10913 => 55,
    10914 => 55,
    10915 => 55,
    10916 => 55,
    10917 => 55,
    10918 => 55,
    10919 => 55,
    10920 => 55,
    10921 => 55,
    10922 => 55,
    10923 => 55,
    10924 => 55,
    10925 => 55,
    10926 => 55,
    10927 => 55,
    10928 => 55,
    10929 => 55,
    10930 => 55,
    10931 => 55,
    10932 => 55,
    10933 => 55,
    10934 => 55,
    10935 => 55,
    10936 => 55,
    10937 => 55,
    10938 => 55,
    10939 => 55,
    10940 => 55,
    10941 => 55,
    10942 => 55,
    10943 => 55,
    10944 => 55,
    10945 => 55,
    10946 => 55,
    10947 => 55,
    10948 => 55,
    10949 => 55,
    10950 => 55,
    10951 => 55,
    10952 => 55,
    10953 => 55,
    10954 => 55,
    10955 => 55,
    10956 => 55,
    10957 => 55,
    10958 => 55,
    10959 => 55,
    10960 => 55,
    10961 => 55,
    10962 => 55,
    10963 => 55,
    10964 => 55,
    10965 => 55,
    10966 => 55,
    10967 => 55,
    10968 => 55,
    10969 => 55,
    10970 => 55,
    10971 => 55,
    10972 => 55,
    10973 => 55,
    10974 => 55,
    10975 => 55,
    10976 => 55,
    10977 => 55,
    10978 => 55,
    10979 => 55,
    10980 => 55,
    10981 => 55,
    10982 => 55,
    10983 => 55,
    10984 => 55,
    10985 => 55,
    10986 => 55,
    10987 => 55,
    10988 => 55,
    10989 => 55,
    10990 => 55,
    10991 => 55,
    10992 => 55,
    10993 => 55,
    10994 => 55,
    10995 => 55,
    10996 => 55,
    10997 => 55,
    10998 => 55,
    10999 => 55,
    11000 => 55,
    11001 => 55,
    11002 => 55,
    11003 => 55,
    11004 => 55,
    11005 => 55,
    11006 => 55,
    11007 => 55,
    11008 => 55,
    11009 => 55,
    11010 => 55,
    11011 => 55,
    11012 => 55,
    11013 => 55,
    11014 => 55,
    11015 => 55,
    11016 => 55,
    11017 => 55,
    11018 => 55,
    11019 => 55,
    11020 => 55,
    11021 => 55,
    11022 => 55,
    11023 => 55,
    11024 => 55,
    11025 => 55,
    11026 => 55,
    11027 => 55,
    11028 => 55,
    11029 => 55,
    11030 => 55,
    11031 => 55,
    11032 => 55,
    11033 => 55,
    11034 => 55,
    11035 => 55,
    11036 => 55,
    11037 => 55,
    11038 => 55,
    11039 => 55,
    11040 => 55,
    11041 => 55,
    11042 => 55,
    11043 => 55,
    11044 => 55,
    11045 => 55,
    11046 => 55,
    11047 => 55,
    11048 => 55,
    11049 => 55,
    11050 => 55,
    11051 => 55,
    11052 => 55,
    11053 => 55,
    11054 => 55,
    11055 => 55,
    11056 => 55,
    11057 => 55,
    11058 => 55,
    11059 => 55,
    11060 => 55,
    11061 => 55,
    11062 => 55,
    11063 => 55,
    11064 => 55,
    11065 => 55,
    11066 => 55,
    11067 => 55,
    11068 => 55,
    11069 => 55,
    11070 => 55,
    11071 => 55,
    11072 => 55,
    11073 => 55,
    11074 => 55,
    11075 => 55,
    11076 => 55,
    11077 => 55,
    11078 => 55,
    11079 => 55,
    11080 => 55,
    11081 => 55,
    11082 => 55,
    11083 => 55,
    11084 => 55,
    11085 => 55,
    11086 => 55,
    11087 => 55,
    11088 => 55,
    11089 => 55,
    11090 => 55,
    11091 => 55,
    11092 => 55,
    11093 => 55,
    11094 => 55,
    11095 => 55,
    11096 => 55,
    11097 => 55,
    11098 => 55,
    11099 => 55,
    11100 => 55,
    11101 => 55,
    11102 => 55,
    11103 => 55,
    11104 => 55,
    11105 => 55,
    11106 => 55,
    11107 => 55,
    11108 => 55,
    11109 => 55,
    11110 => 55,
    11111 => 55,
    11112 => 55,
    11113 => 55,
    11114 => 55,
    11115 => 55,
    11116 => 55,
    11117 => 55,
    11118 => 55,
    11119 => 55,
    11120 => 55,
    11121 => 55,
    11122 => 55,
    11123 => 55,
    11124 => 55,
    11125 => 55,
    11126 => 55,
    11127 => 55,
    11128 => 55,
    11129 => 55,
    11130 => 55,
    11131 => 55,
    11132 => 55,
    11133 => 55,
    11134 => 55,
    11135 => 55,
    11136 => 55,
    11137 => 55,
    11138 => 55,
    11139 => 55,
    11140 => 55,
    11141 => 55,
    11142 => 55,
    11143 => 55,
    11144 => 55,
    11145 => 55,
    11146 => 55,
    11147 => 55,
    11148 => 55,
    11149 => 55,
    11150 => 55,
    11151 => 55,
    11152 => 55,
    11153 => 55,
    11154 => 55,
    11155 => 55,
    11156 => 55,
    11157 => 55,
    11158 => 55,
    11159 => 55,
    11160 => 55,
    11161 => 55,
    11162 => 55,
    11163 => 55,
    11164 => 55,
    11165 => 55,
    11166 => 55,
    11167 => 55,
    11168 => 55,
    11169 => 55,
    11170 => 55,
    11171 => 55,
    11172 => 55,
    11173 => 55,
    11174 => 55,
    11175 => 55,
    11176 => 55,
    11177 => 55,
    11178 => 55,
    11179 => 55,
    11180 => 55,
    11181 => 55,
    11182 => 55,
    11183 => 55,
    11184 => 55,
    11185 => 55,
    11186 => 55,
    11187 => 55,
    11188 => 55,
    11189 => 55,
    11190 => 55,
    11191 => 55,
    11192 => 55,
    11193 => 55,
    11194 => 55,
    11195 => 55,
    11196 => 55,
    11197 => 55,
    11198 => 55,
    11199 => 55,
    11200 => 55,
    11201 => 55,
    11202 => 55,
    11203 => 55,
    11204 => 55,
    11205 => 55,
    11206 => 55,
    11207 => 55,
    11208 => 55,
    11209 => 55,
    11210 => 55,
    11211 => 55,
    11212 => 55,
    11213 => 55,
    11214 => 55,
    11215 => 55,
    11216 => 55,
    11217 => 55,
    11218 => 55,
    11219 => 55,
    11220 => 55,
    11221 => 55,
    11222 => 55,
    11223 => 55,
    11224 => 55,
    11225 => 55,
    11226 => 55,
    11227 => 55,
    11228 => 55,
    11229 => 55,
    11230 => 55,
    11231 => 55,
    11232 => 55,
    11233 => 55,
    11234 => 55,
    11235 => 55,
    11236 => 55,
    11237 => 55,
    11238 => 55,
    11239 => 55,
    11240 => 55,
    11241 => 55,
    11242 => 55,
    11243 => 56,
    11244 => 56,
    11245 => 56,
    11246 => 56,
    11247 => 56,
    11248 => 56,
    11249 => 56,
    11250 => 56,
    11251 => 56,
    11252 => 56,
    11253 => 56,
    11254 => 56,
    11255 => 56,
    11256 => 56,
    11257 => 56,
    11258 => 56,
    11259 => 56,
    11260 => 56,
    11261 => 56,
    11262 => 56,
    11263 => 56,
    11264 => 56,
    11265 => 56,
    11266 => 56,
    11267 => 56,
    11268 => 56,
    11269 => 56,
    11270 => 56,
    11271 => 56,
    11272 => 56,
    11273 => 56,
    11274 => 56,
    11275 => 56,
    11276 => 56,
    11277 => 56,
    11278 => 56,
    11279 => 56,
    11280 => 56,
    11281 => 56,
    11282 => 56,
    11283 => 56,
    11284 => 56,
    11285 => 56,
    11286 => 56,
    11287 => 56,
    11288 => 56,
    11289 => 56,
    11290 => 56,
    11291 => 56,
    11292 => 56,
    11293 => 56,
    11294 => 56,
    11295 => 56,
    11296 => 56,
    11297 => 56,
    11298 => 56,
    11299 => 56,
    11300 => 56,
    11301 => 56,
    11302 => 56,
    11303 => 56,
    11304 => 56,
    11305 => 56,
    11306 => 56,
    11307 => 56,
    11308 => 56,
    11309 => 56,
    11310 => 56,
    11311 => 56,
    11312 => 56,
    11313 => 56,
    11314 => 56,
    11315 => 56,
    11316 => 56,
    11317 => 56,
    11318 => 56,
    11319 => 56,
    11320 => 56,
    11321 => 56,
    11322 => 56,
    11323 => 56,
    11324 => 56,
    11325 => 56,
    11326 => 56,
    11327 => 56,
    11328 => 56,
    11329 => 56,
    11330 => 56,
    11331 => 56,
    11332 => 56,
    11333 => 56,
    11334 => 56,
    11335 => 56,
    11336 => 56,
    11337 => 56,
    11338 => 56,
    11339 => 56,
    11340 => 56,
    11341 => 56,
    11342 => 56,
    11343 => 56,
    11344 => 56,
    11345 => 56,
    11346 => 56,
    11347 => 56,
    11348 => 56,
    11349 => 56,
    11350 => 56,
    11351 => 56,
    11352 => 56,
    11353 => 56,
    11354 => 56,
    11355 => 56,
    11356 => 56,
    11357 => 56,
    11358 => 56,
    11359 => 56,
    11360 => 56,
    11361 => 56,
    11362 => 56,
    11363 => 56,
    11364 => 56,
    11365 => 56,
    11366 => 56,
    11367 => 56,
    11368 => 56,
    11369 => 56,
    11370 => 56,
    11371 => 56,
    11372 => 56,
    11373 => 56,
    11374 => 56,
    11375 => 56,
    11376 => 56,
    11377 => 56,
    11378 => 56,
    11379 => 56,
    11380 => 56,
    11381 => 56,
    11382 => 56,
    11383 => 56,
    11384 => 56,
    11385 => 56,
    11386 => 56,
    11387 => 56,
    11388 => 56,
    11389 => 56,
    11390 => 56,
    11391 => 56,
    11392 => 56,
    11393 => 56,
    11394 => 56,
    11395 => 56,
    11396 => 56,
    11397 => 56,
    11398 => 56,
    11399 => 56,
    11400 => 56,
    11401 => 56,
    11402 => 56,
    11403 => 56,
    11404 => 56,
    11405 => 56,
    11406 => 56,
    11407 => 56,
    11408 => 56,
    11409 => 56,
    11410 => 56,
    11411 => 56,
    11412 => 56,
    11413 => 56,
    11414 => 56,
    11415 => 56,
    11416 => 56,
    11417 => 56,
    11418 => 56,
    11419 => 56,
    11420 => 56,
    11421 => 56,
    11422 => 56,
    11423 => 56,
    11424 => 56,
    11425 => 56,
    11426 => 56,
    11427 => 56,
    11428 => 56,
    11429 => 56,
    11430 => 56,
    11431 => 56,
    11432 => 56,
    11433 => 56,
    11434 => 56,
    11435 => 56,
    11436 => 56,
    11437 => 56,
    11438 => 56,
    11439 => 56,
    11440 => 56,
    11441 => 56,
    11442 => 56,
    11443 => 56,
    11444 => 56,
    11445 => 56,
    11446 => 56,
    11447 => 56,
    11448 => 56,
    11449 => 56,
    11450 => 56,
    11451 => 56,
    11452 => 56,
    11453 => 56,
    11454 => 56,
    11455 => 56,
    11456 => 56,
    11457 => 56,
    11458 => 56,
    11459 => 56,
    11460 => 56,
    11461 => 56,
    11462 => 56,
    11463 => 56,
    11464 => 56,
    11465 => 56,
    11466 => 56,
    11467 => 56,
    11468 => 56,
    11469 => 56,
    11470 => 56,
    11471 => 56,
    11472 => 56,
    11473 => 56,
    11474 => 56,
    11475 => 56,
    11476 => 56,
    11477 => 56,
    11478 => 56,
    11479 => 56,
    11480 => 56,
    11481 => 56,
    11482 => 56,
    11483 => 56,
    11484 => 56,
    11485 => 56,
    11486 => 56,
    11487 => 56,
    11488 => 56,
    11489 => 56,
    11490 => 56,
    11491 => 56,
    11492 => 56,
    11493 => 56,
    11494 => 56,
    11495 => 56,
    11496 => 56,
    11497 => 56,
    11498 => 56,
    11499 => 56,
    11500 => 56,
    11501 => 56,
    11502 => 56,
    11503 => 56,
    11504 => 56,
    11505 => 56,
    11506 => 56,
    11507 => 56,
    11508 => 56,
    11509 => 56,
    11510 => 56,
    11511 => 56,
    11512 => 56,
    11513 => 56,
    11514 => 56,
    11515 => 56,
    11516 => 56,
    11517 => 56,
    11518 => 56,
    11519 => 56,
    11520 => 56,
    11521 => 56,
    11522 => 56,
    11523 => 56,
    11524 => 56,
    11525 => 56,
    11526 => 56,
    11527 => 56,
    11528 => 56,
    11529 => 56,
    11530 => 56,
    11531 => 56,
    11532 => 56,
    11533 => 56,
    11534 => 56,
    11535 => 56,
    11536 => 56,
    11537 => 56,
    11538 => 56,
    11539 => 56,
    11540 => 56,
    11541 => 56,
    11542 => 56,
    11543 => 56,
    11544 => 56,
    11545 => 56,
    11546 => 56,
    11547 => 56,
    11548 => 56,
    11549 => 56,
    11550 => 56,
    11551 => 56,
    11552 => 56,
    11553 => 56,
    11554 => 56,
    11555 => 56,
    11556 => 56,
    11557 => 56,
    11558 => 56,
    11559 => 56,
    11560 => 56,
    11561 => 56,
    11562 => 56,
    11563 => 56,
    11564 => 56,
    11565 => 56,
    11566 => 56,
    11567 => 56,
    11568 => 56,
    11569 => 56,
    11570 => 56,
    11571 => 56,
    11572 => 56,
    11573 => 56,
    11574 => 56,
    11575 => 56,
    11576 => 56,
    11577 => 56,
    11578 => 56,
    11579 => 56,
    11580 => 56,
    11581 => 56,
    11582 => 56,
    11583 => 56,
    11584 => 56,
    11585 => 56,
    11586 => 56,
    11587 => 56,
    11588 => 56,
    11589 => 56,
    11590 => 56,
    11591 => 56,
    11592 => 56,
    11593 => 56,
    11594 => 56,
    11595 => 56,
    11596 => 56,
    11597 => 56,
    11598 => 56,
    11599 => 56,
    11600 => 56,
    11601 => 56,
    11602 => 56,
    11603 => 56,
    11604 => 56,
    11605 => 57,
    11606 => 57,
    11607 => 57,
    11608 => 57,
    11609 => 57,
    11610 => 57,
    11611 => 57,
    11612 => 57,
    11613 => 57,
    11614 => 57,
    11615 => 57,
    11616 => 57,
    11617 => 57,
    11618 => 57,
    11619 => 57,
    11620 => 57,
    11621 => 57,
    11622 => 57,
    11623 => 57,
    11624 => 57,
    11625 => 57,
    11626 => 57,
    11627 => 57,
    11628 => 57,
    11629 => 57,
    11630 => 57,
    11631 => 57,
    11632 => 57,
    11633 => 57,
    11634 => 57,
    11635 => 57,
    11636 => 57,
    11637 => 57,
    11638 => 57,
    11639 => 57,
    11640 => 57,
    11641 => 57,
    11642 => 57,
    11643 => 57,
    11644 => 57,
    11645 => 57,
    11646 => 57,
    11647 => 57,
    11648 => 57,
    11649 => 57,
    11650 => 57,
    11651 => 57,
    11652 => 57,
    11653 => 57,
    11654 => 57,
    11655 => 57,
    11656 => 57,
    11657 => 57,
    11658 => 57,
    11659 => 57,
    11660 => 57,
    11661 => 57,
    11662 => 57,
    11663 => 57,
    11664 => 57,
    11665 => 57,
    11666 => 57,
    11667 => 57,
    11668 => 57,
    11669 => 57,
    11670 => 57,
    11671 => 57,
    11672 => 57,
    11673 => 57,
    11674 => 57,
    11675 => 57,
    11676 => 57,
    11677 => 57,
    11678 => 57,
    11679 => 57,
    11680 => 57,
    11681 => 57,
    11682 => 57,
    11683 => 57,
    11684 => 57,
    11685 => 57,
    11686 => 57,
    11687 => 57,
    11688 => 57,
    11689 => 57,
    11690 => 57,
    11691 => 57,
    11692 => 57,
    11693 => 57,
    11694 => 57,
    11695 => 57,
    11696 => 57,
    11697 => 57,
    11698 => 57,
    11699 => 57,
    11700 => 57,
    11701 => 57,
    11702 => 57,
    11703 => 57,
    11704 => 57,
    11705 => 57,
    11706 => 57,
    11707 => 57,
    11708 => 57,
    11709 => 57,
    11710 => 57,
    11711 => 57,
    11712 => 57,
    11713 => 57,
    11714 => 57,
    11715 => 57,
    11716 => 57,
    11717 => 57,
    11718 => 57,
    11719 => 57,
    11720 => 57,
    11721 => 57,
    11722 => 57,
    11723 => 57,
    11724 => 57,
    11725 => 57,
    11726 => 57,
    11727 => 57,
    11728 => 57,
    11729 => 57,
    11730 => 57,
    11731 => 57,
    11732 => 57,
    11733 => 57,
    11734 => 57,
    11735 => 57,
    11736 => 57,
    11737 => 57,
    11738 => 57,
    11739 => 57,
    11740 => 57,
    11741 => 57,
    11742 => 57,
    11743 => 57,
    11744 => 57,
    11745 => 57,
    11746 => 57,
    11747 => 57,
    11748 => 57,
    11749 => 57,
    11750 => 57,
    11751 => 57,
    11752 => 57,
    11753 => 57,
    11754 => 57,
    11755 => 57,
    11756 => 57,
    11757 => 57,
    11758 => 57,
    11759 => 57,
    11760 => 57,
    11761 => 57,
    11762 => 57,
    11763 => 57,
    11764 => 57,
    11765 => 57,
    11766 => 57,
    11767 => 57,
    11768 => 57,
    11769 => 57,
    11770 => 57,
    11771 => 57,
    11772 => 57,
    11773 => 57,
    11774 => 57,
    11775 => 57,
    11776 => 57,
    11777 => 57,
    11778 => 57,
    11779 => 57,
    11780 => 57,
    11781 => 57,
    11782 => 57,
    11783 => 57,
    11784 => 57,
    11785 => 57,
    11786 => 57,
    11787 => 57,
    11788 => 57,
    11789 => 57,
    11790 => 57,
    11791 => 57,
    11792 => 57,
    11793 => 57,
    11794 => 57,
    11795 => 57,
    11796 => 57,
    11797 => 57,
    11798 => 57,
    11799 => 57,
    11800 => 57,
    11801 => 57,
    11802 => 57,
    11803 => 57,
    11804 => 57,
    11805 => 57,
    11806 => 57,
    11807 => 57,
    11808 => 57,
    11809 => 57,
    11810 => 57,
    11811 => 57,
    11812 => 57,
    11813 => 57,
    11814 => 57,
    11815 => 57,
    11816 => 57,
    11817 => 57,
    11818 => 57,
    11819 => 57,
    11820 => 57,
    11821 => 57,
    11822 => 57,
    11823 => 57,
    11824 => 57,
    11825 => 57,
    11826 => 57,
    11827 => 57,
    11828 => 57,
    11829 => 57,
    11830 => 57,
    11831 => 57,
    11832 => 57,
    11833 => 57,
    11834 => 57,
    11835 => 57,
    11836 => 57,
    11837 => 57,
    11838 => 57,
    11839 => 57,
    11840 => 57,
    11841 => 57,
    11842 => 57,
    11843 => 57,
    11844 => 57,
    11845 => 57,
    11846 => 57,
    11847 => 57,
    11848 => 57,
    11849 => 57,
    11850 => 57,
    11851 => 57,
    11852 => 57,
    11853 => 57,
    11854 => 57,
    11855 => 57,
    11856 => 57,
    11857 => 57,
    11858 => 57,
    11859 => 57,
    11860 => 57,
    11861 => 57,
    11862 => 57,
    11863 => 57,
    11864 => 57,
    11865 => 57,
    11866 => 57,
    11867 => 57,
    11868 => 57,
    11869 => 57,
    11870 => 57,
    11871 => 57,
    11872 => 57,
    11873 => 57,
    11874 => 57,
    11875 => 57,
    11876 => 57,
    11877 => 57,
    11878 => 57,
    11879 => 57,
    11880 => 57,
    11881 => 57,
    11882 => 57,
    11883 => 57,
    11884 => 57,
    11885 => 57,
    11886 => 57,
    11887 => 57,
    11888 => 57,
    11889 => 57,
    11890 => 57,
    11891 => 57,
    11892 => 57,
    11893 => 57,
    11894 => 57,
    11895 => 57,
    11896 => 57,
    11897 => 57,
    11898 => 57,
    11899 => 57,
    11900 => 57,
    11901 => 57,
    11902 => 57,
    11903 => 57,
    11904 => 57,
    11905 => 57,
    11906 => 57,
    11907 => 57,
    11908 => 57,
    11909 => 57,
    11910 => 57,
    11911 => 57,
    11912 => 57,
    11913 => 57,
    11914 => 57,
    11915 => 57,
    11916 => 57,
    11917 => 57,
    11918 => 57,
    11919 => 57,
    11920 => 57,
    11921 => 57,
    11922 => 57,
    11923 => 57,
    11924 => 57,
    11925 => 57,
    11926 => 57,
    11927 => 57,
    11928 => 57,
    11929 => 57,
    11930 => 57,
    11931 => 57,
    11932 => 57,
    11933 => 57,
    11934 => 57,
    11935 => 57,
    11936 => 57,
    11937 => 57,
    11938 => 57,
    11939 => 57,
    11940 => 57,
    11941 => 57,
    11942 => 57,
    11943 => 57,
    11944 => 57,
    11945 => 57,
    11946 => 57,
    11947 => 57,
    11948 => 57,
    11949 => 57,
    11950 => 57,
    11951 => 57,
    11952 => 57,
    11953 => 57,
    11954 => 57,
    11955 => 57,
    11956 => 57,
    11957 => 57,
    11958 => 57,
    11959 => 57,
    11960 => 57,
    11961 => 57,
    11962 => 57,
    11963 => 57,
    11964 => 57,
    11965 => 57,
    11966 => 57,
    11967 => 57,
    11968 => 57,
    11969 => 57,
    11970 => 57,
    11971 => 57,
    11972 => 57,
    11973 => 57,
    11974 => 57,
    11975 => 57,
    11976 => 57,
    11977 => 57,
    11978 => 57,
    11979 => 57,
    11980 => 57,
    11981 => 57,
    11982 => 57,
    11983 => 57,
    11984 => 57,
    11985 => 57,
    11986 => 57,
    11987 => 57,
    11988 => 57,
    11989 => 57,
    11990 => 57,
    11991 => 57,
    11992 => 57,
    11993 => 57,
    11994 => 58,
    11995 => 58,
    11996 => 58,
    11997 => 58,
    11998 => 58,
    11999 => 58,
    12000 => 58,
    12001 => 58,
    12002 => 58,
    12003 => 58,
    12004 => 58,
    12005 => 58,
    12006 => 58,
    12007 => 58,
    12008 => 58,
    12009 => 58,
    12010 => 58,
    12011 => 58,
    12012 => 58,
    12013 => 58,
    12014 => 58,
    12015 => 58,
    12016 => 58,
    12017 => 58,
    12018 => 58,
    12019 => 58,
    12020 => 58,
    12021 => 58,
    12022 => 58,
    12023 => 58,
    12024 => 58,
    12025 => 58,
    12026 => 58,
    12027 => 58,
    12028 => 58,
    12029 => 58,
    12030 => 58,
    12031 => 58,
    12032 => 58,
    12033 => 58,
    12034 => 58,
    12035 => 58,
    12036 => 58,
    12037 => 58,
    12038 => 58,
    12039 => 58,
    12040 => 58,
    12041 => 58,
    12042 => 58,
    12043 => 58,
    12044 => 58,
    12045 => 58,
    12046 => 58,
    12047 => 58,
    12048 => 58,
    12049 => 58,
    12050 => 58,
    12051 => 58,
    12052 => 58,
    12053 => 58,
    12054 => 58,
    12055 => 58,
    12056 => 58,
    12057 => 58,
    12058 => 58,
    12059 => 58,
    12060 => 58,
    12061 => 58,
    12062 => 58,
    12063 => 58,
    12064 => 58,
    12065 => 58,
    12066 => 58,
    12067 => 58,
    12068 => 58,
    12069 => 58,
    12070 => 58,
    12071 => 58,
    12072 => 58,
    12073 => 58,
    12074 => 58,
    12075 => 58,
    12076 => 58,
    12077 => 58,
    12078 => 58,
    12079 => 58,
    12080 => 58,
    12081 => 58,
    12082 => 58,
    12083 => 58,
    12084 => 58,
    12085 => 58,
    12086 => 58,
    12087 => 58,
    12088 => 58,
    12089 => 58,
    12090 => 58,
    12091 => 58,
    12092 => 58,
    12093 => 58,
    12094 => 58,
    12095 => 58,
    12096 => 58,
    12097 => 58,
    12098 => 58,
    12099 => 58,
    12100 => 58,
    12101 => 58,
    12102 => 58,
    12103 => 58,
    12104 => 58,
    12105 => 58,
    12106 => 58,
    12107 => 58,
    12108 => 58,
    12109 => 58,
    12110 => 58,
    12111 => 58,
    12112 => 58,
    12113 => 58,
    12114 => 58,
    12115 => 58,
    12116 => 58,
    12117 => 58,
    12118 => 58,
    12119 => 58,
    12120 => 58,
    12121 => 58,
    12122 => 58,
    12123 => 58,
    12124 => 58,
    12125 => 58,
    12126 => 58,
    12127 => 58,
    12128 => 58,
    12129 => 58,
    12130 => 58,
    12131 => 58,
    12132 => 58,
    12133 => 58,
    12134 => 58,
    12135 => 58,
    12136 => 58,
    12137 => 58,
    12138 => 58,
    12139 => 58,
    12140 => 58,
    12141 => 58,
    12142 => 58,
    12143 => 58,
    12144 => 58,
    12145 => 58,
    12146 => 58,
    12147 => 58,
    12148 => 58,
    12149 => 58,
    12150 => 58,
    12151 => 58,
    12152 => 58,
    12153 => 58,
    12154 => 58,
    12155 => 58,
    12156 => 58,
    12157 => 58,
    12158 => 58,
    12159 => 58,
    12160 => 58,
    12161 => 58,
    12162 => 58,
    12163 => 58,
    12164 => 58,
    12165 => 58,
    12166 => 58,
    12167 => 58,
    12168 => 58,
    12169 => 58,
    12170 => 58,
    12171 => 58,
    12172 => 58,
    12173 => 58,
    12174 => 58,
    12175 => 58,
    12176 => 58,
    12177 => 58,
    12178 => 58,
    12179 => 58,
    12180 => 58,
    12181 => 58,
    12182 => 58,
    12183 => 58,
    12184 => 58,
    12185 => 58,
    12186 => 58,
    12187 => 58,
    12188 => 58,
    12189 => 58,
    12190 => 58,
    12191 => 58,
    12192 => 58,
    12193 => 58,
    12194 => 58,
    12195 => 58,
    12196 => 58,
    12197 => 58,
    12198 => 58,
    12199 => 58,
    12200 => 58,
    12201 => 58,
    12202 => 58,
    12203 => 58,
    12204 => 58,
    12205 => 58,
    12206 => 58,
    12207 => 58,
    12208 => 58,
    12209 => 58,
    12210 => 58,
    12211 => 58,
    12212 => 58,
    12213 => 58,
    12214 => 58,
    12215 => 58,
    12216 => 58,
    12217 => 58,
    12218 => 58,
    12219 => 58,
    12220 => 58,
    12221 => 58,
    12222 => 58,
    12223 => 58,
    12224 => 58,
    12225 => 58,
    12226 => 58,
    12227 => 58,
    12228 => 58,
    12229 => 58,
    12230 => 58,
    12231 => 58,
    12232 => 58,
    12233 => 58,
    12234 => 58,
    12235 => 58,
    12236 => 58,
    12237 => 58,
    12238 => 58,
    12239 => 58,
    12240 => 58,
    12241 => 58,
    12242 => 58,
    12243 => 58,
    12244 => 58,
    12245 => 58,
    12246 => 58,
    12247 => 58,
    12248 => 58,
    12249 => 58,
    12250 => 58,
    12251 => 58,
    12252 => 58,
    12253 => 58,
    12254 => 58,
    12255 => 58,
    12256 => 58,
    12257 => 58,
    12258 => 58,
    12259 => 58,
    12260 => 58,
    12261 => 58,
    12262 => 58,
    12263 => 58,
    12264 => 58,
    12265 => 58,
    12266 => 58,
    12267 => 58,
    12268 => 58,
    12269 => 58,
    12270 => 58,
    12271 => 58,
    12272 => 58,
    12273 => 58,
    12274 => 58,
    12275 => 58,
    12276 => 58,
    12277 => 58,
    12278 => 58,
    12279 => 58,
    12280 => 58,
    12281 => 58,
    12282 => 58,
    12283 => 58,
    12284 => 58,
    12285 => 58,
    12286 => 58,
    12287 => 58,
    12288 => 58,
    12289 => 58,
    12290 => 58,
    12291 => 58,
    12292 => 58,
    12293 => 58,
    12294 => 58,
    12295 => 58,
    12296 => 58,
    12297 => 58,
    12298 => 58,
    12299 => 58,
    12300 => 58,
    12301 => 58,
    12302 => 58,
    12303 => 58,
    12304 => 58,
    12305 => 58,
    12306 => 58,
    12307 => 58,
    12308 => 58,
    12309 => 58,
    12310 => 58,
    12311 => 58,
    12312 => 58,
    12313 => 58,
    12314 => 58,
    12315 => 58,
    12316 => 58,
    12317 => 58,
    12318 => 58,
    12319 => 58,
    12320 => 58,
    12321 => 58,
    12322 => 58,
    12323 => 58,
    12324 => 58,
    12325 => 58,
    12326 => 58,
    12327 => 58,
    12328 => 58,
    12329 => 58,
    12330 => 58,
    12331 => 58,
    12332 => 58,
    12333 => 58,
    12334 => 58,
    12335 => 58,
    12336 => 58,
    12337 => 58,
    12338 => 58,
    12339 => 58,
    12340 => 58,
    12341 => 58,
    12342 => 58,
    12343 => 58,
    12344 => 58,
    12345 => 58,
    12346 => 58,
    12347 => 58,
    12348 => 58,
    12349 => 58,
    12350 => 58,
    12351 => 58,
    12352 => 58,
    12353 => 58,
    12354 => 58,
    12355 => 58,
    12356 => 58,
    12357 => 58,
    12358 => 58,
    12359 => 58,
    12360 => 58,
    12361 => 58,
    12362 => 58,
    12363 => 58,
    12364 => 58,
    12365 => 58,
    12366 => 58,
    12367 => 58,
    12368 => 58,
    12369 => 58,
    12370 => 58,
    12371 => 58,
    12372 => 58,
    12373 => 58,
    12374 => 58,
    12375 => 58,
    12376 => 58,
    12377 => 58,
    12378 => 58,
    12379 => 58,
    12380 => 58,
    12381 => 58,
    12382 => 58,
    12383 => 58,
    12384 => 58,
    12385 => 58,
    12386 => 58,
    12387 => 58,
    12388 => 58,
    12389 => 58,
    12390 => 58,
    12391 => 58,
    12392 => 58,
    12393 => 58,
    12394 => 58,
    12395 => 58,
    12396 => 58,
    12397 => 58,
    12398 => 58,
    12399 => 58,
    12400 => 58,
    12401 => 58,
    12402 => 58,
    12403 => 58,
    12404 => 58,
    12405 => 58,
    12406 => 58,
    12407 => 58,
    12408 => 58,
    12409 => 58,
    12410 => 58,
    12411 => 58,
    12412 => 58,
    12413 => 58,
    12414 => 58,
    12415 => 58,
    12416 => 58,
    12417 => 58,
    12418 => 59,
    12419 => 59,
    12420 => 59,
    12421 => 59,
    12422 => 59,
    12423 => 59,
    12424 => 59,
    12425 => 59,
    12426 => 59,
    12427 => 59,
    12428 => 59,
    12429 => 59,
    12430 => 59,
    12431 => 59,
    12432 => 59,
    12433 => 59,
    12434 => 59,
    12435 => 59,
    12436 => 59,
    12437 => 59,
    12438 => 59,
    12439 => 59,
    12440 => 59,
    12441 => 59,
    12442 => 59,
    12443 => 59,
    12444 => 59,
    12445 => 59,
    12446 => 59,
    12447 => 59,
    12448 => 59,
    12449 => 59,
    12450 => 59,
    12451 => 59,
    12452 => 59,
    12453 => 59,
    12454 => 59,
    12455 => 59,
    12456 => 59,
    12457 => 59,
    12458 => 59,
    12459 => 59,
    12460 => 59,
    12461 => 59,
    12462 => 59,
    12463 => 59,
    12464 => 59,
    12465 => 59,
    12466 => 59,
    12467 => 59,
    12468 => 59,
    12469 => 59,
    12470 => 59,
    12471 => 59,
    12472 => 59,
    12473 => 59,
    12474 => 59,
    12475 => 59,
    12476 => 59,
    12477 => 59,
    12478 => 59,
    12479 => 59,
    12480 => 59,
    12481 => 59,
    12482 => 59,
    12483 => 59,
    12484 => 59,
    12485 => 59,
    12486 => 59,
    12487 => 59,
    12488 => 59,
    12489 => 59,
    12490 => 59,
    12491 => 59,
    12492 => 59,
    12493 => 59,
    12494 => 59,
    12495 => 59,
    12496 => 59,
    12497 => 59,
    12498 => 59,
    12499 => 59,
    12500 => 59,
    12501 => 59,
    12502 => 59,
    12503 => 59,
    12504 => 59,
    12505 => 59,
    12506 => 59,
    12507 => 59,
    12508 => 59,
    12509 => 59,
    12510 => 59,
    12511 => 59,
    12512 => 59,
    12513 => 59,
    12514 => 59,
    12515 => 59,
    12516 => 59,
    12517 => 59,
    12518 => 59,
    12519 => 59,
    12520 => 59,
    12521 => 59,
    12522 => 59,
    12523 => 59,
    12524 => 59,
    12525 => 59,
    12526 => 59,
    12527 => 59,
    12528 => 59,
    12529 => 59,
    12530 => 59,
    12531 => 59,
    12532 => 59,
    12533 => 59,
    12534 => 59,
    12535 => 59,
    12536 => 59,
    12537 => 59,
    12538 => 59,
    12539 => 59,
    12540 => 59,
    12541 => 59,
    12542 => 59,
    12543 => 59,
    12544 => 59,
    12545 => 59,
    12546 => 59,
    12547 => 59,
    12548 => 59,
    12549 => 59,
    12550 => 59,
    12551 => 59,
    12552 => 59,
    12553 => 59,
    12554 => 59,
    12555 => 59,
    12556 => 59,
    12557 => 59,
    12558 => 59,
    12559 => 59,
    12560 => 59,
    12561 => 59,
    12562 => 59,
    12563 => 59,
    12564 => 59,
    12565 => 59,
    12566 => 59,
    12567 => 59,
    12568 => 59,
    12569 => 59,
    12570 => 59,
    12571 => 59,
    12572 => 59,
    12573 => 59,
    12574 => 59,
    12575 => 59,
    12576 => 59,
    12577 => 59,
    12578 => 59,
    12579 => 59,
    12580 => 59,
    12581 => 59,
    12582 => 59,
    12583 => 59,
    12584 => 59,
    12585 => 59,
    12586 => 59,
    12587 => 59,
    12588 => 59,
    12589 => 59,
    12590 => 59,
    12591 => 59,
    12592 => 59,
    12593 => 59,
    12594 => 59,
    12595 => 59,
    12596 => 59,
    12597 => 59,
    12598 => 59,
    12599 => 59,
    12600 => 59,
    12601 => 59,
    12602 => 59,
    12603 => 59,
    12604 => 59,
    12605 => 59,
    12606 => 59,
    12607 => 59,
    12608 => 59,
    12609 => 59,
    12610 => 59,
    12611 => 59,
    12612 => 59,
    12613 => 59,
    12614 => 59,
    12615 => 59,
    12616 => 59,
    12617 => 59,
    12618 => 59,
    12619 => 59,
    12620 => 59,
    12621 => 59,
    12622 => 59,
    12623 => 59,
    12624 => 59,
    12625 => 59,
    12626 => 59,
    12627 => 59,
    12628 => 59,
    12629 => 59,
    12630 => 59,
    12631 => 59,
    12632 => 59,
    12633 => 59,
    12634 => 59,
    12635 => 59,
    12636 => 59,
    12637 => 59,
    12638 => 59,
    12639 => 59,
    12640 => 59,
    12641 => 59,
    12642 => 59,
    12643 => 59,
    12644 => 59,
    12645 => 59,
    12646 => 59,
    12647 => 59,
    12648 => 59,
    12649 => 59,
    12650 => 59,
    12651 => 59,
    12652 => 59,
    12653 => 59,
    12654 => 59,
    12655 => 59,
    12656 => 59,
    12657 => 59,
    12658 => 59,
    12659 => 59,
    12660 => 59,
    12661 => 59,
    12662 => 59,
    12663 => 59,
    12664 => 59,
    12665 => 59,
    12666 => 59,
    12667 => 59,
    12668 => 59,
    12669 => 59,
    12670 => 59,
    12671 => 59,
    12672 => 59,
    12673 => 59,
    12674 => 59,
    12675 => 59,
    12676 => 59,
    12677 => 59,
    12678 => 59,
    12679 => 59,
    12680 => 59,
    12681 => 59,
    12682 => 59,
    12683 => 59,
    12684 => 59,
    12685 => 59,
    12686 => 59,
    12687 => 59,
    12688 => 59,
    12689 => 59,
    12690 => 59,
    12691 => 59,
    12692 => 59,
    12693 => 59,
    12694 => 59,
    12695 => 59,
    12696 => 59,
    12697 => 59,
    12698 => 59,
    12699 => 59,
    12700 => 59,
    12701 => 59,
    12702 => 59,
    12703 => 59,
    12704 => 59,
    12705 => 59,
    12706 => 59,
    12707 => 59,
    12708 => 59,
    12709 => 59,
    12710 => 59,
    12711 => 59,
    12712 => 59,
    12713 => 59,
    12714 => 59,
    12715 => 59,
    12716 => 59,
    12717 => 59,
    12718 => 59,
    12719 => 59,
    12720 => 59,
    12721 => 59,
    12722 => 59,
    12723 => 59,
    12724 => 59,
    12725 => 59,
    12726 => 59,
    12727 => 59,
    12728 => 59,
    12729 => 59,
    12730 => 59,
    12731 => 59,
    12732 => 59,
    12733 => 59,
    12734 => 59,
    12735 => 59,
    12736 => 59,
    12737 => 59,
    12738 => 59,
    12739 => 59,
    12740 => 59,
    12741 => 59,
    12742 => 59,
    12743 => 59,
    12744 => 59,
    12745 => 59,
    12746 => 59,
    12747 => 59,
    12748 => 59,
    12749 => 59,
    12750 => 59,
    12751 => 59,
    12752 => 59,
    12753 => 59,
    12754 => 59,
    12755 => 59,
    12756 => 59,
    12757 => 59,
    12758 => 59,
    12759 => 59,
    12760 => 59,
    12761 => 59,
    12762 => 59,
    12763 => 59,
    12764 => 59,
    12765 => 59,
    12766 => 59,
    12767 => 59,
    12768 => 59,
    12769 => 59,
    12770 => 59,
    12771 => 59,
    12772 => 59,
    12773 => 59,
    12774 => 59,
    12775 => 59,
    12776 => 59,
    12777 => 59,
    12778 => 59,
    12779 => 59,
    12780 => 59,
    12781 => 59,
    12782 => 59,
    12783 => 59,
    12784 => 59,
    12785 => 59,
    12786 => 59,
    12787 => 59,
    12788 => 59,
    12789 => 59,
    12790 => 59,
    12791 => 59,
    12792 => 59,
    12793 => 59,
    12794 => 59,
    12795 => 59,
    12796 => 59,
    12797 => 59,
    12798 => 59,
    12799 => 59,
    12800 => 59,
    12801 => 59,
    12802 => 59,
    12803 => 59,
    12804 => 59,
    12805 => 59,
    12806 => 59,
    12807 => 59,
    12808 => 59,
    12809 => 59,
    12810 => 59,
    12811 => 59,
    12812 => 59,
    12813 => 59,
    12814 => 59,
    12815 => 59,
    12816 => 59,
    12817 => 59,
    12818 => 59,
    12819 => 59,
    12820 => 59,
    12821 => 59,
    12822 => 59,
    12823 => 59,
    12824 => 59,
    12825 => 59,
    12826 => 59,
    12827 => 59,
    12828 => 59,
    12829 => 59,
    12830 => 59,
    12831 => 59,
    12832 => 59,
    12833 => 59,
    12834 => 59,
    12835 => 59,
    12836 => 59,
    12837 => 59,
    12838 => 59,
    12839 => 59,
    12840 => 59,
    12841 => 59,
    12842 => 59,
    12843 => 59,
    12844 => 59,
    12845 => 59,
    12846 => 59,
    12847 => 59,
    12848 => 59,
    12849 => 59,
    12850 => 59,
    12851 => 59,
    12852 => 59,
    12853 => 59,
    12854 => 59,
    12855 => 59,
    12856 => 59,
    12857 => 59,
    12858 => 59,
    12859 => 59,
    12860 => 59,
    12861 => 59,
    12862 => 59,
    12863 => 59,
    12864 => 59,
    12865 => 59,
    12866 => 59,
    12867 => 59,
    12868 => 59,
    12869 => 59,
    12870 => 59,
    12871 => 59,
    12872 => 59,
    12873 => 59,
    12874 => 59,
    12875 => 59,
    12876 => 59,
    12877 => 59,
    12878 => 59,
    12879 => 59,
    12880 => 59,
    12881 => 59,
    12882 => 59,
    12883 => 59,
    12884 => 59,
    12885 => 59,
    12886 => 59,
    12887 => 59,
    12888 => 59,
    12889 => 59,
    12890 => 59,
    12891 => 60,
    12892 => 60,
    12893 => 60,
    12894 => 60,
    12895 => 60,
    12896 => 60,
    12897 => 60,
    12898 => 60,
    12899 => 60,
    12900 => 60,
    12901 => 60,
    12902 => 60,
    12903 => 60,
    12904 => 60,
    12905 => 60,
    12906 => 60,
    12907 => 60,
    12908 => 60,
    12909 => 60,
    12910 => 60,
    12911 => 60,
    12912 => 60,
    12913 => 60,
    12914 => 60,
    12915 => 60,
    12916 => 60,
    12917 => 60,
    12918 => 60,
    12919 => 60,
    12920 => 60,
    12921 => 60,
    12922 => 60,
    12923 => 60,
    12924 => 60,
    12925 => 60,
    12926 => 60,
    12927 => 60,
    12928 => 60,
    12929 => 60,
    12930 => 60,
    12931 => 60,
    12932 => 60,
    12933 => 60,
    12934 => 60,
    12935 => 60,
    12936 => 60,
    12937 => 60,
    12938 => 60,
    12939 => 60,
    12940 => 60,
    12941 => 60,
    12942 => 60,
    12943 => 60,
    12944 => 60,
    12945 => 60,
    12946 => 60,
    12947 => 60,
    12948 => 60,
    12949 => 60,
    12950 => 60,
    12951 => 60,
    12952 => 60,
    12953 => 60,
    12954 => 60,
    12955 => 60,
    12956 => 60,
    12957 => 60,
    12958 => 60,
    12959 => 60,
    12960 => 60,
    12961 => 60,
    12962 => 60,
    12963 => 60,
    12964 => 60,
    12965 => 60,
    12966 => 60,
    12967 => 60,
    12968 => 60,
    12969 => 60,
    12970 => 60,
    12971 => 60,
    12972 => 60,
    12973 => 60,
    12974 => 60,
    12975 => 60,
    12976 => 60,
    12977 => 60,
    12978 => 60,
    12979 => 60,
    12980 => 60,
    12981 => 60,
    12982 => 60,
    12983 => 60,
    12984 => 60,
    12985 => 60,
    12986 => 60,
    12987 => 60,
    12988 => 60,
    12989 => 60,
    12990 => 60,
    12991 => 60,
    12992 => 60,
    12993 => 60,
    12994 => 60,
    12995 => 60,
    12996 => 60,
    12997 => 60,
    12998 => 60,
    12999 => 60,
    13000 => 60,
    13001 => 60,
    13002 => 60,
    13003 => 60,
    13004 => 60,
    13005 => 60,
    13006 => 60,
    13007 => 60,
    13008 => 60,
    13009 => 60,
    13010 => 60,
    13011 => 60,
    13012 => 60,
    13013 => 60,
    13014 => 60,
    13015 => 60,
    13016 => 60,
    13017 => 60,
    13018 => 60,
    13019 => 60,
    13020 => 60,
    13021 => 60,
    13022 => 60,
    13023 => 60,
    13024 => 60,
    13025 => 60,
    13026 => 60,
    13027 => 60,
    13028 => 60,
    13029 => 60,
    13030 => 60,
    13031 => 60,
    13032 => 60,
    13033 => 60,
    13034 => 60,
    13035 => 60,
    13036 => 60,
    13037 => 60,
    13038 => 60,
    13039 => 60,
    13040 => 60,
    13041 => 60,
    13042 => 60,
    13043 => 60,
    13044 => 60,
    13045 => 60,
    13046 => 60,
    13047 => 60,
    13048 => 60,
    13049 => 60,
    13050 => 60,
    13051 => 60,
    13052 => 60,
    13053 => 60,
    13054 => 60,
    13055 => 60,
    13056 => 60,
    13057 => 60,
    13058 => 60,
    13059 => 60,
    13060 => 60,
    13061 => 60,
    13062 => 60,
    13063 => 60,
    13064 => 60,
    13065 => 60,
    13066 => 60,
    13067 => 60,
    13068 => 60,
    13069 => 60,
    13070 => 60,
    13071 => 60,
    13072 => 60,
    13073 => 60,
    13074 => 60,
    13075 => 60,
    13076 => 60,
    13077 => 60,
    13078 => 60,
    13079 => 60,
    13080 => 60,
    13081 => 60,
    13082 => 60,
    13083 => 60,
    13084 => 60,
    13085 => 60,
    13086 => 60,
    13087 => 60,
    13088 => 60,
    13089 => 60,
    13090 => 60,
    13091 => 60,
    13092 => 60,
    13093 => 60,
    13094 => 60,
    13095 => 60,
    13096 => 60,
    13097 => 60,
    13098 => 60,
    13099 => 60,
    13100 => 60,
    13101 => 60,
    13102 => 60,
    13103 => 60,
    13104 => 60,
    13105 => 60,
    13106 => 60,
    13107 => 60,
    13108 => 60,
    13109 => 60,
    13110 => 60,
    13111 => 60,
    13112 => 60,
    13113 => 60,
    13114 => 60,
    13115 => 60,
    13116 => 60,
    13117 => 60,
    13118 => 60,
    13119 => 60,
    13120 => 60,
    13121 => 60,
    13122 => 60,
    13123 => 60,
    13124 => 60,
    13125 => 60,
    13126 => 60,
    13127 => 60,
    13128 => 60,
    13129 => 60,
    13130 => 60,
    13131 => 60,
    13132 => 60,
    13133 => 60,
    13134 => 60,
    13135 => 60,
    13136 => 60,
    13137 => 60,
    13138 => 60,
    13139 => 60,
    13140 => 60,
    13141 => 60,
    13142 => 60,
    13143 => 60,
    13144 => 60,
    13145 => 60,
    13146 => 60,
    13147 => 60,
    13148 => 60,
    13149 => 60,
    13150 => 60,
    13151 => 60,
    13152 => 60,
    13153 => 60,
    13154 => 60,
    13155 => 60,
    13156 => 60,
    13157 => 60,
    13158 => 60,
    13159 => 60,
    13160 => 60,
    13161 => 60,
    13162 => 60,
    13163 => 60,
    13164 => 60,
    13165 => 60,
    13166 => 60,
    13167 => 60,
    13168 => 60,
    13169 => 60,
    13170 => 60,
    13171 => 60,
    13172 => 60,
    13173 => 60,
    13174 => 60,
    13175 => 60,
    13176 => 60,
    13177 => 60,
    13178 => 60,
    13179 => 60,
    13180 => 60,
    13181 => 60,
    13182 => 60,
    13183 => 60,
    13184 => 60,
    13185 => 60,
    13186 => 60,
    13187 => 60,
    13188 => 60,
    13189 => 60,
    13190 => 60,
    13191 => 60,
    13192 => 60,
    13193 => 60,
    13194 => 60,
    13195 => 60,
    13196 => 60,
    13197 => 60,
    13198 => 60,
    13199 => 60,
    13200 => 60,
    13201 => 60,
    13202 => 60,
    13203 => 60,
    13204 => 60,
    13205 => 60,
    13206 => 60,
    13207 => 60,
    13208 => 60,
    13209 => 60,
    13210 => 60,
    13211 => 60,
    13212 => 60,
    13213 => 60,
    13214 => 60,
    13215 => 60,
    13216 => 60,
    13217 => 60,
    13218 => 60,
    13219 => 60,
    13220 => 60,
    13221 => 60,
    13222 => 60,
    13223 => 60,
    13224 => 60,
    13225 => 60,
    13226 => 60,
    13227 => 60,
    13228 => 60,
    13229 => 60,
    13230 => 60,
    13231 => 60,
    13232 => 60,
    13233 => 60,
    13234 => 60,
    13235 => 60,
    13236 => 60,
    13237 => 60,
    13238 => 60,
    13239 => 60,
    13240 => 60,
    13241 => 60,
    13242 => 60,
    13243 => 60,
    13244 => 60,
    13245 => 60,
    13246 => 60,
    13247 => 60,
    13248 => 60,
    13249 => 60,
    13250 => 60,
    13251 => 60,
    13252 => 60,
    13253 => 60,
    13254 => 60,
    13255 => 60,
    13256 => 60,
    13257 => 60,
    13258 => 60,
    13259 => 60,
    13260 => 60,
    13261 => 60,
    13262 => 60,
    13263 => 60,
    13264 => 60,
    13265 => 60,
    13266 => 60,
    13267 => 60,
    13268 => 60,
    13269 => 60,
    13270 => 60,
    13271 => 60,
    13272 => 60,
    13273 => 60,
    13274 => 60,
    13275 => 60,
    13276 => 60,
    13277 => 60,
    13278 => 60,
    13279 => 60,
    13280 => 60,
    13281 => 60,
    13282 => 60,
    13283 => 60,
    13284 => 60,
    13285 => 60,
    13286 => 60,
    13287 => 60,
    13288 => 60,
    13289 => 60,
    13290 => 60,
    13291 => 60,
    13292 => 60,
    13293 => 60,
    13294 => 60,
    13295 => 60,
    13296 => 60,
    13297 => 60,
    13298 => 60,
    13299 => 60,
    13300 => 60,
    13301 => 60,
    13302 => 60,
    13303 => 60,
    13304 => 60,
    13305 => 60,
    13306 => 60,
    13307 => 60,
    13308 => 60,
    13309 => 60,
    13310 => 60,
    13311 => 60,
    13312 => 60,
    13313 => 60,
    13314 => 60,
    13315 => 60,
    13316 => 60,
    13317 => 60,
    13318 => 60,
    13319 => 60,
    13320 => 60,
    13321 => 60,
    13322 => 60,
    13323 => 60,
    13324 => 60,
    13325 => 60,
    13326 => 60,
    13327 => 60,
    13328 => 60,
    13329 => 60,
    13330 => 60,
    13331 => 60,
    13332 => 60,
    13333 => 60,
    13334 => 60,
    13335 => 60,
    13336 => 60,
    13337 => 60,
    13338 => 60,
    13339 => 60,
    13340 => 60,
    13341 => 60,
    13342 => 60,
    13343 => 60,
    13344 => 60,
    13345 => 60,
    13346 => 60,
    13347 => 60,
    13348 => 60,
    13349 => 60,
    13350 => 60,
    13351 => 60,
    13352 => 60,
    13353 => 60,
    13354 => 60,
    13355 => 60,
    13356 => 60,
    13357 => 60,
    13358 => 60,
    13359 => 60,
    13360 => 60,
    13361 => 60,
    13362 => 60,
    13363 => 60,
    13364 => 60,
    13365 => 60,
    13366 => 60,
    13367 => 60,
    13368 => 60,
    13369 => 60,
    13370 => 60,
    13371 => 60,
    13372 => 60,
    13373 => 60,
    13374 => 60,
    13375 => 60,
    13376 => 60,
    13377 => 60,
    13378 => 60,
    13379 => 60,
    13380 => 60,
    13381 => 60,
    13382 => 60,
    13383 => 60,
    13384 => 60,
    13385 => 60,
    13386 => 60,
    13387 => 60,
    13388 => 60,
    13389 => 60,
    13390 => 60,
    13391 => 60,
    13392 => 60,
    13393 => 60,
    13394 => 60,
    13395 => 60,
    13396 => 60,
    13397 => 60,
    13398 => 60,
    13399 => 60,
    13400 => 60,
    13401 => 60,
    13402 => 60,
    13403 => 60,
    13404 => 60,
    13405 => 60,
    13406 => 60,
    13407 => 60,
    13408 => 60,
    13409 => 60,
    13410 => 60,
    13411 => 60,
    13412 => 60,
    13413 => 60,
    13414 => 60,
    13415 => 60,
    13416 => 60,
    13417 => 60,
    13418 => 60,
    13419 => 60,
    13420 => 60,
    13421 => 60,
    13422 => 60,
    13423 => 60,
    13424 => 60,
    13425 => 60,
    13426 => 60,
    13427 => 60,
    13428 => 60,
    13429 => 60,
    13430 => 60,
    13431 => 60,
    13432 => 60,
    13433 => 60,
    13434 => 60,
    13435 => 60,
    13436 => 61,
    13437 => 61,
    13438 => 61,
    13439 => 61,
    13440 => 61,
    13441 => 61,
    13442 => 61,
    13443 => 61,
    13444 => 61,
    13445 => 61,
    13446 => 61,
    13447 => 61,
    13448 => 61,
    13449 => 61,
    13450 => 61,
    13451 => 61,
    13452 => 61,
    13453 => 61,
    13454 => 61,
    13455 => 61,
    13456 => 61,
    13457 => 61,
    13458 => 61,
    13459 => 61,
    13460 => 61,
    13461 => 61,
    13462 => 61,
    13463 => 61,
    13464 => 61,
    13465 => 61,
    13466 => 61,
    13467 => 61,
    13468 => 61,
    13469 => 61,
    13470 => 61,
    13471 => 61,
    13472 => 61,
    13473 => 61,
    13474 => 61,
    13475 => 61,
    13476 => 61,
    13477 => 61,
    13478 => 61,
    13479 => 61,
    13480 => 61,
    13481 => 61,
    13482 => 61,
    13483 => 61,
    13484 => 61,
    13485 => 61,
    13486 => 61,
    13487 => 61,
    13488 => 61,
    13489 => 61,
    13490 => 61,
    13491 => 61,
    13492 => 61,
    13493 => 61,
    13494 => 61,
    13495 => 61,
    13496 => 61,
    13497 => 61,
    13498 => 61,
    13499 => 61,
    13500 => 61,
    13501 => 61,
    13502 => 61,
    13503 => 61,
    13504 => 61,
    13505 => 61,
    13506 => 61,
    13507 => 61,
    13508 => 61,
    13509 => 61,
    13510 => 61,
    13511 => 61,
    13512 => 61,
    13513 => 61,
    13514 => 61,
    13515 => 61,
    13516 => 61,
    13517 => 61,
    13518 => 61,
    13519 => 61,
    13520 => 61,
    13521 => 61,
    13522 => 61,
    13523 => 61,
    13524 => 61,
    13525 => 61,
    13526 => 61,
    13527 => 61,
    13528 => 61,
    13529 => 61,
    13530 => 61,
    13531 => 61,
    13532 => 61,
    13533 => 61,
    13534 => 61,
    13535 => 61,
    13536 => 61,
    13537 => 61,
    13538 => 61,
    13539 => 61,
    13540 => 61,
    13541 => 61,
    13542 => 61,
    13543 => 61,
    13544 => 61,
    13545 => 61,
    13546 => 61,
    13547 => 61,
    13548 => 61,
    13549 => 61,
    13550 => 61,
    13551 => 61,
    13552 => 61,
    13553 => 61,
    13554 => 61,
    13555 => 61,
    13556 => 61,
    13557 => 61,
    13558 => 61,
    13559 => 61,
    13560 => 61,
    13561 => 61,
    13562 => 61,
    13563 => 61,
    13564 => 61,
    13565 => 61,
    13566 => 61,
    13567 => 61,
    13568 => 61,
    13569 => 61,
    13570 => 61,
    13571 => 61,
    13572 => 61,
    13573 => 61,
    13574 => 61,
    13575 => 61,
    13576 => 61,
    13577 => 61,
    13578 => 61,
    13579 => 61,
    13580 => 61,
    13581 => 61,
    13582 => 61,
    13583 => 61,
    13584 => 61,
    13585 => 61,
    13586 => 61,
    13587 => 61,
    13588 => 61,
    13589 => 61,
    13590 => 61,
    13591 => 61,
    13592 => 61,
    13593 => 61,
    13594 => 61,
    13595 => 61,
    13596 => 61,
    13597 => 61,
    13598 => 61,
    13599 => 61,
    13600 => 61,
    13601 => 61,
    13602 => 61,
    13603 => 61,
    13604 => 61,
    13605 => 61,
    13606 => 61,
    13607 => 61,
    13608 => 61,
    13609 => 61,
    13610 => 61,
    13611 => 61,
    13612 => 61,
    13613 => 61,
    13614 => 61,
    13615 => 61,
    13616 => 61,
    13617 => 61,
    13618 => 61,
    13619 => 61,
    13620 => 61,
    13621 => 61,
    13622 => 61,
    13623 => 61,
    13624 => 61,
    13625 => 61,
    13626 => 61,
    13627 => 61,
    13628 => 61,
    13629 => 61,
    13630 => 61,
    13631 => 61,
    13632 => 61,
    13633 => 61,
    13634 => 61,
    13635 => 61,
    13636 => 61,
    13637 => 61,
    13638 => 61,
    13639 => 61,
    13640 => 61,
    13641 => 61,
    13642 => 61,
    13643 => 61,
    13644 => 61,
    13645 => 61,
    13646 => 61,
    13647 => 61,
    13648 => 61,
    13649 => 61,
    13650 => 61,
    13651 => 61,
    13652 => 61,
    13653 => 61,
    13654 => 61,
    13655 => 61,
    13656 => 61,
    13657 => 61,
    13658 => 61,
    13659 => 61,
    13660 => 61,
    13661 => 61,
    13662 => 61,
    13663 => 61,
    13664 => 61,
    13665 => 61,
    13666 => 61,
    13667 => 61,
    13668 => 61,
    13669 => 61,
    13670 => 61,
    13671 => 61,
    13672 => 61,
    13673 => 61,
    13674 => 61,
    13675 => 61,
    13676 => 61,
    13677 => 61,
    13678 => 61,
    13679 => 61,
    13680 => 61,
    13681 => 61,
    13682 => 61,
    13683 => 61,
    13684 => 61,
    13685 => 61,
    13686 => 61,
    13687 => 61,
    13688 => 61,
    13689 => 61,
    13690 => 61,
    13691 => 61,
    13692 => 61,
    13693 => 61,
    13694 => 61,
    13695 => 61,
    13696 => 61,
    13697 => 61,
    13698 => 61,
    13699 => 61,
    13700 => 61,
    13701 => 61,
    13702 => 61,
    13703 => 61,
    13704 => 61,
    13705 => 61,
    13706 => 61,
    13707 => 61,
    13708 => 61,
    13709 => 61,
    13710 => 61,
    13711 => 61,
    13712 => 61,
    13713 => 61,
    13714 => 61,
    13715 => 61,
    13716 => 61,
    13717 => 61,
    13718 => 61,
    13719 => 61,
    13720 => 61,
    13721 => 61,
    13722 => 61,
    13723 => 61,
    13724 => 61,
    13725 => 61,
    13726 => 61,
    13727 => 61,
    13728 => 61,
    13729 => 61,
    13730 => 61,
    13731 => 61,
    13732 => 61,
    13733 => 61,
    13734 => 61,
    13735 => 61,
    13736 => 61,
    13737 => 61,
    13738 => 61,
    13739 => 61,
    13740 => 61,
    13741 => 61,
    13742 => 61,
    13743 => 61,
    13744 => 61,
    13745 => 61,
    13746 => 61,
    13747 => 61,
    13748 => 61,
    13749 => 61,
    13750 => 61,
    13751 => 61,
    13752 => 61,
    13753 => 61,
    13754 => 61,
    13755 => 61,
    13756 => 61,
    13757 => 61,
    13758 => 61,
    13759 => 61,
    13760 => 61,
    13761 => 61,
    13762 => 61,
    13763 => 61,
    13764 => 61,
    13765 => 61,
    13766 => 61,
    13767 => 61,
    13768 => 61,
    13769 => 61,
    13770 => 61,
    13771 => 61,
    13772 => 61,
    13773 => 61,
    13774 => 61,
    13775 => 61,
    13776 => 61,
    13777 => 61,
    13778 => 61,
    13779 => 61,
    13780 => 61,
    13781 => 61,
    13782 => 61,
    13783 => 61,
    13784 => 61,
    13785 => 61,
    13786 => 61,
    13787 => 61,
    13788 => 61,
    13789 => 61,
    13790 => 61,
    13791 => 61,
    13792 => 61,
    13793 => 61,
    13794 => 61,
    13795 => 61,
    13796 => 61,
    13797 => 61,
    13798 => 61,
    13799 => 61,
    13800 => 61,
    13801 => 61,
    13802 => 61,
    13803 => 61,
    13804 => 61,
    13805 => 61,
    13806 => 61,
    13807 => 61,
    13808 => 61,
    13809 => 61,
    13810 => 61,
    13811 => 61,
    13812 => 61,
    13813 => 61,
    13814 => 61,
    13815 => 61,
    13816 => 61,
    13817 => 61,
    13818 => 61,
    13819 => 61,
    13820 => 61,
    13821 => 61,
    13822 => 61,
    13823 => 61,
    13824 => 61,
    13825 => 61,
    13826 => 61,
    13827 => 61,
    13828 => 61,
    13829 => 61,
    13830 => 61,
    13831 => 61,
    13832 => 61,
    13833 => 61,
    13834 => 61,
    13835 => 61,
    13836 => 61,
    13837 => 61,
    13838 => 61,
    13839 => 61,
    13840 => 61,
    13841 => 61,
    13842 => 61,
    13843 => 61,
    13844 => 61,
    13845 => 61,
    13846 => 61,
    13847 => 61,
    13848 => 61,
    13849 => 61,
    13850 => 61,
    13851 => 61,
    13852 => 61,
    13853 => 61,
    13854 => 61,
    13855 => 61,
    13856 => 61,
    13857 => 61,
    13858 => 61,
    13859 => 61,
    13860 => 61,
    13861 => 61,
    13862 => 61,
    13863 => 61,
    13864 => 61,
    13865 => 61,
    13866 => 61,
    13867 => 61,
    13868 => 61,
    13869 => 61,
    13870 => 61,
    13871 => 61,
    13872 => 61,
    13873 => 61,
    13874 => 61,
    13875 => 61,
    13876 => 61,
    13877 => 61,
    13878 => 61,
    13879 => 61,
    13880 => 61,
    13881 => 61,
    13882 => 61,
    13883 => 61,
    13884 => 61,
    13885 => 61,
    13886 => 61,
    13887 => 61,
    13888 => 61,
    13889 => 61,
    13890 => 61,
    13891 => 61,
    13892 => 61,
    13893 => 61,
    13894 => 61,
    13895 => 61,
    13896 => 61,
    13897 => 61,
    13898 => 61,
    13899 => 61,
    13900 => 61,
    13901 => 61,
    13902 => 61,
    13903 => 61,
    13904 => 61,
    13905 => 61,
    13906 => 61,
    13907 => 61,
    13908 => 61,
    13909 => 61,
    13910 => 61,
    13911 => 61,
    13912 => 61,
    13913 => 61,
    13914 => 61,
    13915 => 61,
    13916 => 61,
    13917 => 61,
    13918 => 61,
    13919 => 61,
    13920 => 61,
    13921 => 61,
    13922 => 61,
    13923 => 61,
    13924 => 61,
    13925 => 61,
    13926 => 61,
    13927 => 61,
    13928 => 61,
    13929 => 61,
    13930 => 61,
    13931 => 61,
    13932 => 61,
    13933 => 61,
    13934 => 61,
    13935 => 61,
    13936 => 61,
    13937 => 61,
    13938 => 61,
    13939 => 61,
    13940 => 61,
    13941 => 61,
    13942 => 61,
    13943 => 61,
    13944 => 61,
    13945 => 61,
    13946 => 61,
    13947 => 61,
    13948 => 61,
    13949 => 61,
    13950 => 61,
    13951 => 61,
    13952 => 61,
    13953 => 61,
    13954 => 61,
    13955 => 61,
    13956 => 61,
    13957 => 61,
    13958 => 61,
    13959 => 61,
    13960 => 61,
    13961 => 61,
    13962 => 61,
    13963 => 61,
    13964 => 61,
    13965 => 61,
    13966 => 61,
    13967 => 61,
    13968 => 61,
    13969 => 61,
    13970 => 61,
    13971 => 61,
    13972 => 61,
    13973 => 61,
    13974 => 61,
    13975 => 61,
    13976 => 61,
    13977 => 61,
    13978 => 61,
    13979 => 61,
    13980 => 61,
    13981 => 61,
    13982 => 61,
    13983 => 61,
    13984 => 61,
    13985 => 61,
    13986 => 61,
    13987 => 61,
    13988 => 61,
    13989 => 61,
    13990 => 61,
    13991 => 61,
    13992 => 61,
    13993 => 61,
    13994 => 61,
    13995 => 61,
    13996 => 61,
    13997 => 61,
    13998 => 61,
    13999 => 61,
    14000 => 61,
    14001 => 61,
    14002 => 61,
    14003 => 61,
    14004 => 61,
    14005 => 61,
    14006 => 61,
    14007 => 61,
    14008 => 61,
    14009 => 61,
    14010 => 61,
    14011 => 61,
    14012 => 61,
    14013 => 61,
    14014 => 61,
    14015 => 61,
    14016 => 61,
    14017 => 61,
    14018 => 61,
    14019 => 61,
    14020 => 61,
    14021 => 61,
    14022 => 61,
    14023 => 61,
    14024 => 61,
    14025 => 61,
    14026 => 61,
    14027 => 61,
    14028 => 61,
    14029 => 61,
    14030 => 61,
    14031 => 61,
    14032 => 61,
    14033 => 61,
    14034 => 61,
    14035 => 61,
    14036 => 61,
    14037 => 61,
    14038 => 61,
    14039 => 61,
    14040 => 61,
    14041 => 61,
    14042 => 61,
    14043 => 61,
    14044 => 61,
    14045 => 61,
    14046 => 61,
    14047 => 61,
    14048 => 61,
    14049 => 61,
    14050 => 61,
    14051 => 61,
    14052 => 61,
    14053 => 61,
    14054 => 61,
    14055 => 61,
    14056 => 61,
    14057 => 61,
    14058 => 61,
    14059 => 61,
    14060 => 61,
    14061 => 61,
    14062 => 61,
    14063 => 61,
    14064 => 61,
    14065 => 61,
    14066 => 61,
    14067 => 61,
    14068 => 61,
    14069 => 61,
    14070 => 61,
    14071 => 61,
    14072 => 61,
    14073 => 61,
    14074 => 61,
    14075 => 61,
    14076 => 61,
    14077 => 61,
    14078 => 61,
    14079 => 61,
    14080 => 61,
    14081 => 61,
    14082 => 61,
    14083 => 61,
    14084 => 61,
    14085 => 61,
    14086 => 61,
    14087 => 61,
    14088 => 61,
    14089 => 61,
    14090 => 61,
    14091 => 61,
    14092 => 61,
    14093 => 61,
    14094 => 61,
    14095 => 61,
    14096 => 61,
    14097 => 61,
    14098 => 61,
    14099 => 61,
    14100 => 61,
    14101 => 61,
    14102 => 61,
    14103 => 61,
    14104 => 62,
    14105 => 62,
    14106 => 62,
    14107 => 62,
    14108 => 62,
    14109 => 62,
    14110 => 62,
    14111 => 62,
    14112 => 62,
    14113 => 62,
    14114 => 62,
    14115 => 62,
    14116 => 62,
    14117 => 62,
    14118 => 62,
    14119 => 62,
    14120 => 62,
    14121 => 62,
    14122 => 62,
    14123 => 62,
    14124 => 62,
    14125 => 62,
    14126 => 62,
    14127 => 62,
    14128 => 62,
    14129 => 62,
    14130 => 62,
    14131 => 62,
    14132 => 62,
    14133 => 62,
    14134 => 62,
    14135 => 62,
    14136 => 62,
    14137 => 62,
    14138 => 62,
    14139 => 62,
    14140 => 62,
    14141 => 62,
    14142 => 62,
    14143 => 62,
    14144 => 62,
    14145 => 62,
    14146 => 62,
    14147 => 62,
    14148 => 62,
    14149 => 62,
    14150 => 62,
    14151 => 62,
    14152 => 62,
    14153 => 62,
    14154 => 62,
    14155 => 62,
    14156 => 62,
    14157 => 62,
    14158 => 62,
    14159 => 62,
    14160 => 62,
    14161 => 62,
    14162 => 62,
    14163 => 62,
    14164 => 62,
    14165 => 62,
    14166 => 62,
    14167 => 62,
    14168 => 62,
    14169 => 62,
    14170 => 62,
    14171 => 62,
    14172 => 62,
    14173 => 62,
    14174 => 62,
    14175 => 62,
    14176 => 62,
    14177 => 62,
    14178 => 62,
    14179 => 62,
    14180 => 62,
    14181 => 62,
    14182 => 62,
    14183 => 62,
    14184 => 62,
    14185 => 62,
    14186 => 62,
    14187 => 62,
    14188 => 62,
    14189 => 62,
    14190 => 62,
    14191 => 62,
    14192 => 62,
    14193 => 62,
    14194 => 62,
    14195 => 62,
    14196 => 62,
    14197 => 62,
    14198 => 62,
    14199 => 62,
    14200 => 62,
    14201 => 62,
    14202 => 62,
    14203 => 62,
    14204 => 62,
    14205 => 62,
    14206 => 62,
    14207 => 62,
    14208 => 62,
    14209 => 62,
    14210 => 62,
    14211 => 62,
    14212 => 62,
    14213 => 62,
    14214 => 62,
    14215 => 62,
    14216 => 62,
    14217 => 62,
    14218 => 62,
    14219 => 62,
    14220 => 62,
    14221 => 62,
    14222 => 62,
    14223 => 62,
    14224 => 62,
    14225 => 62,
    14226 => 62,
    14227 => 62,
    14228 => 62,
    14229 => 62,
    14230 => 62,
    14231 => 62,
    14232 => 62,
    14233 => 62,
    14234 => 62,
    14235 => 62,
    14236 => 62,
    14237 => 62,
    14238 => 62,
    14239 => 62,
    14240 => 62,
    14241 => 62,
    14242 => 62,
    14243 => 62,
    14244 => 62,
    14245 => 62,
    14246 => 62,
    14247 => 62,
    14248 => 62,
    14249 => 62,
    14250 => 62,
    14251 => 62,
    14252 => 62,
    14253 => 62,
    14254 => 62,
    14255 => 62,
    14256 => 62,
    14257 => 62,
    14258 => 62,
    14259 => 62,
    14260 => 62,
    14261 => 62,
    14262 => 62,
    14263 => 62,
    14264 => 62,
    14265 => 62,
    14266 => 62,
    14267 => 62,
    14268 => 62,
    14269 => 62,
    14270 => 62,
    14271 => 62,
    14272 => 62,
    14273 => 62,
    14274 => 62,
    14275 => 62,
    14276 => 62,
    14277 => 62,
    14278 => 62,
    14279 => 62,
    14280 => 62,
    14281 => 62,
    14282 => 62,
    14283 => 62,
    14284 => 62,
    14285 => 62,
    14286 => 62,
    14287 => 62,
    14288 => 62,
    14289 => 62,
    14290 => 62,
    14291 => 62,
    14292 => 62,
    14293 => 62,
    14294 => 62,
    14295 => 62,
    14296 => 62,
    14297 => 62,
    14298 => 62,
    14299 => 62,
    14300 => 62,
    14301 => 62,
    14302 => 62,
    14303 => 62,
    14304 => 62,
    14305 => 62,
    14306 => 62,
    14307 => 62,
    14308 => 62,
    14309 => 62,
    14310 => 62,
    14311 => 62,
    14312 => 62,
    14313 => 62,
    14314 => 62,
    14315 => 62,
    14316 => 62,
    14317 => 62,
    14318 => 62,
    14319 => 62,
    14320 => 62,
    14321 => 62,
    14322 => 62,
    14323 => 62,
    14324 => 62,
    14325 => 62,
    14326 => 62,
    14327 => 62,
    14328 => 62,
    14329 => 62,
    14330 => 62,
    14331 => 62,
    14332 => 62,
    14333 => 62,
    14334 => 62,
    14335 => 62,
    14336 => 62,
    14337 => 62,
    14338 => 62,
    14339 => 62,
    14340 => 62,
    14341 => 62,
    14342 => 62,
    14343 => 62,
    14344 => 62,
    14345 => 62,
    14346 => 62,
    14347 => 62,
    14348 => 62,
    14349 => 62,
    14350 => 62,
    14351 => 62,
    14352 => 62,
    14353 => 62,
    14354 => 62,
    14355 => 62,
    14356 => 62,
    14357 => 62,
    14358 => 62,
    14359 => 62,
    14360 => 62,
    14361 => 62,
    14362 => 62,
    14363 => 62,
    14364 => 62,
    14365 => 62,
    14366 => 62,
    14367 => 62,
    14368 => 62,
    14369 => 62,
    14370 => 62,
    14371 => 62,
    14372 => 62,
    14373 => 62,
    14374 => 62,
    14375 => 62,
    14376 => 62,
    14377 => 62,
    14378 => 62,
    14379 => 62,
    14380 => 62,
    14381 => 62,
    14382 => 62,
    14383 => 62,
    14384 => 62,
    14385 => 62,
    14386 => 62,
    14387 => 62,
    14388 => 62,
    14389 => 62,
    14390 => 62,
    14391 => 62,
    14392 => 62,
    14393 => 62,
    14394 => 62,
    14395 => 62,
    14396 => 62,
    14397 => 62,
    14398 => 62,
    14399 => 62,
    14400 => 62,
    14401 => 62,
    14402 => 62,
    14403 => 62,
    14404 => 62,
    14405 => 62,
    14406 => 62,
    14407 => 62,
    14408 => 62,
    14409 => 62,
    14410 => 62,
    14411 => 62,
    14412 => 62,
    14413 => 62,
    14414 => 62,
    14415 => 62,
    14416 => 62,
    14417 => 62,
    14418 => 62,
    14419 => 62,
    14420 => 62,
    14421 => 62,
    14422 => 62,
    14423 => 62,
    14424 => 62,
    14425 => 62,
    14426 => 62,
    14427 => 62,
    14428 => 62,
    14429 => 62,
    14430 => 62,
    14431 => 62,
    14432 => 62,
    14433 => 62,
    14434 => 62,
    14435 => 62,
    14436 => 62,
    14437 => 62,
    14438 => 62,
    14439 => 62,
    14440 => 62,
    14441 => 62,
    14442 => 62,
    14443 => 62,
    14444 => 62,
    14445 => 62,
    14446 => 62,
    14447 => 62,
    14448 => 62,
    14449 => 62,
    14450 => 62,
    14451 => 62,
    14452 => 62,
    14453 => 62,
    14454 => 62,
    14455 => 62,
    14456 => 62,
    14457 => 62,
    14458 => 62,
    14459 => 62,
    14460 => 62,
    14461 => 62,
    14462 => 62,
    14463 => 62,
    14464 => 62,
    14465 => 62,
    14466 => 62,
    14467 => 62,
    14468 => 62,
    14469 => 62,
    14470 => 62,
    14471 => 62,
    14472 => 62,
    14473 => 62,
    14474 => 62,
    14475 => 62,
    14476 => 62,
    14477 => 62,
    14478 => 62,
    14479 => 62,
    14480 => 62,
    14481 => 62,
    14482 => 62,
    14483 => 62,
    14484 => 62,
    14485 => 62,
    14486 => 62,
    14487 => 62,
    14488 => 62,
    14489 => 62,
    14490 => 62,
    14491 => 62,
    14492 => 62,
    14493 => 62,
    14494 => 62,
    14495 => 62,
    14496 => 62,
    14497 => 62,
    14498 => 62,
    14499 => 62,
    14500 => 62,
    14501 => 62,
    14502 => 62,
    14503 => 62,
    14504 => 62,
    14505 => 62,
    14506 => 62,
    14507 => 62,
    14508 => 62,
    14509 => 62,
    14510 => 62,
    14511 => 62,
    14512 => 62,
    14513 => 62,
    14514 => 62,
    14515 => 62,
    14516 => 62,
    14517 => 62,
    14518 => 62,
    14519 => 62,
    14520 => 62,
    14521 => 62,
    14522 => 62,
    14523 => 62,
    14524 => 62,
    14525 => 62,
    14526 => 62,
    14527 => 62,
    14528 => 62,
    14529 => 62,
    14530 => 62,
    14531 => 62,
    14532 => 62,
    14533 => 62,
    14534 => 62,
    14535 => 62,
    14536 => 62,
    14537 => 62,
    14538 => 62,
    14539 => 62,
    14540 => 62,
    14541 => 62,
    14542 => 62,
    14543 => 62,
    14544 => 62,
    14545 => 62,
    14546 => 62,
    14547 => 62,
    14548 => 62,
    14549 => 62,
    14550 => 62,
    14551 => 62,
    14552 => 62,
    14553 => 62,
    14554 => 62,
    14555 => 62,
    14556 => 62,
    14557 => 62,
    14558 => 62,
    14559 => 62,
    14560 => 62,
    14561 => 62,
    14562 => 62,
    14563 => 62,
    14564 => 62,
    14565 => 62,
    14566 => 62,
    14567 => 62,
    14568 => 62,
    14569 => 62,
    14570 => 62,
    14571 => 62,
    14572 => 62,
    14573 => 62,
    14574 => 62,
    14575 => 62,
    14576 => 62,
    14577 => 62,
    14578 => 62,
    14579 => 62,
    14580 => 62,
    14581 => 62,
    14582 => 62,
    14583 => 62,
    14584 => 62,
    14585 => 62,
    14586 => 62,
    14587 => 62,
    14588 => 62,
    14589 => 62,
    14590 => 62,
    14591 => 62,
    14592 => 62,
    14593 => 62,
    14594 => 62,
    14595 => 62,
    14596 => 62,
    14597 => 62,
    14598 => 62,
    14599 => 62,
    14600 => 62,
    14601 => 62,
    14602 => 62,
    14603 => 62,
    14604 => 62,
    14605 => 62,
    14606 => 62,
    14607 => 62,
    14608 => 62,
    14609 => 62,
    14610 => 62,
    14611 => 62,
    14612 => 62,
    14613 => 62,
    14614 => 62,
    14615 => 62,
    14616 => 62,
    14617 => 62,
    14618 => 62,
    14619 => 62,
    14620 => 62,
    14621 => 62,
    14622 => 62,
    14623 => 62,
    14624 => 62,
    14625 => 62,
    14626 => 62,
    14627 => 62,
    14628 => 62,
    14629 => 62,
    14630 => 62,
    14631 => 62,
    14632 => 62,
    14633 => 62,
    14634 => 62,
    14635 => 62,
    14636 => 62,
    14637 => 62,
    14638 => 62,
    14639 => 62,
    14640 => 62,
    14641 => 62,
    14642 => 62,
    14643 => 62,
    14644 => 62,
    14645 => 62,
    14646 => 62,
    14647 => 62,
    14648 => 62,
    14649 => 62,
    14650 => 62,
    14651 => 62,
    14652 => 62,
    14653 => 62,
    14654 => 62,
    14655 => 62,
    14656 => 62,
    14657 => 62,
    14658 => 62,
    14659 => 62,
    14660 => 62,
    14661 => 62,
    14662 => 62,
    14663 => 62,
    14664 => 62,
    14665 => 62,
    14666 => 62,
    14667 => 62,
    14668 => 62,
    14669 => 62,
    14670 => 62,
    14671 => 62,
    14672 => 62,
    14673 => 62,
    14674 => 62,
    14675 => 62,
    14676 => 62,
    14677 => 62,
    14678 => 62,
    14679 => 62,
    14680 => 62,
    14681 => 62,
    14682 => 62,
    14683 => 62,
    14684 => 62,
    14685 => 62,
    14686 => 62,
    14687 => 62,
    14688 => 62,
    14689 => 62,
    14690 => 62,
    14691 => 62,
    14692 => 62,
    14693 => 62,
    14694 => 62,
    14695 => 62,
    14696 => 62,
    14697 => 62,
    14698 => 62,
    14699 => 62,
    14700 => 62,
    14701 => 62,
    14702 => 62,
    14703 => 62,
    14704 => 62,
    14705 => 62,
    14706 => 62,
    14707 => 62,
    14708 => 62,
    14709 => 62,
    14710 => 62,
    14711 => 62,
    14712 => 62,
    14713 => 62,
    14714 => 62,
    14715 => 62,
    14716 => 62,
    14717 => 62,
    14718 => 62,
    14719 => 62,
    14720 => 62,
    14721 => 62,
    14722 => 62,
    14723 => 62,
    14724 => 62,
    14725 => 62,
    14726 => 62,
    14727 => 62,
    14728 => 62,
    14729 => 62,
    14730 => 62,
    14731 => 62,
    14732 => 62,
    14733 => 62,
    14734 => 62,
    14735 => 62,
    14736 => 62,
    14737 => 62,
    14738 => 62,
    14739 => 62,
    14740 => 62,
    14741 => 62,
    14742 => 62,
    14743 => 62,
    14744 => 62,
    14745 => 62,
    14746 => 62,
    14747 => 62,
    14748 => 62,
    14749 => 62,
    14750 => 62,
    14751 => 62,
    14752 => 62,
    14753 => 62,
    14754 => 62,
    14755 => 62,
    14756 => 62,
    14757 => 62,
    14758 => 62,
    14759 => 62,
    14760 => 62,
    14761 => 62,
    14762 => 62,
    14763 => 62,
    14764 => 62,
    14765 => 62,
    14766 => 62,
    14767 => 62,
    14768 => 62,
    14769 => 62,
    14770 => 62,
    14771 => 62,
    14772 => 62,
    14773 => 62,
    14774 => 62,
    14775 => 62,
    14776 => 62,
    14777 => 62,
    14778 => 62,
    14779 => 62,
    14780 => 62,
    14781 => 62,
    14782 => 62,
    14783 => 62,
    14784 => 62,
    14785 => 62,
    14786 => 62,
    14787 => 62,
    14788 => 62,
    14789 => 62,
    14790 => 62,
    14791 => 62,
    14792 => 62,
    14793 => 62,
    14794 => 62,
    14795 => 62,
    14796 => 62,
    14797 => 62,
    14798 => 62,
    14799 => 62,
    14800 => 62,
    14801 => 62,
    14802 => 62,
    14803 => 62,
    14804 => 62,
    14805 => 62,
    14806 => 62,
    14807 => 62,
    14808 => 62,
    14809 => 62,
    14810 => 62,
    14811 => 62,
    14812 => 62,
    14813 => 62,
    14814 => 62,
    14815 => 62,
    14816 => 62,
    14817 => 62,
    14818 => 62,
    14819 => 62,
    14820 => 62,
    14821 => 62,
    14822 => 62,
    14823 => 62,
    14824 => 62,
    14825 => 62,
    14826 => 62,
    14827 => 62,
    14828 => 62,
    14829 => 62,
    14830 => 62,
    14831 => 62,
    14832 => 62,
    14833 => 62,
    14834 => 62,
    14835 => 62,
    14836 => 62,
    14837 => 62,
    14838 => 62,
    14839 => 62,
    14840 => 62,
    14841 => 62,
    14842 => 62,
    14843 => 62,
    14844 => 62,
    14845 => 62,
    14846 => 62,
    14847 => 62,
    14848 => 62,
    14849 => 62,
    14850 => 62,
    14851 => 62,
    14852 => 62,
    14853 => 62,
    14854 => 62,
    14855 => 62,
    14856 => 62,
    14857 => 62,
    14858 => 62,
    14859 => 62,
    14860 => 62,
    14861 => 62,
    14862 => 62,
    14863 => 62,
    14864 => 62,
    14865 => 62,
    14866 => 62,
    14867 => 62,
    14868 => 62,
    14869 => 62,
    14870 => 62,
    14871 => 62,
    14872 => 62,
    14873 => 62,
    14874 => 62,
    14875 => 62,
    14876 => 62,
    14877 => 62,
    14878 => 62,
    14879 => 62,
    14880 => 62,
    14881 => 62,
    14882 => 62,
    14883 => 62,
    14884 => 62,
    14885 => 62,
    14886 => 62,
    14887 => 62,
    14888 => 62,
    14889 => 62,
    14890 => 62,
    14891 => 62,
    14892 => 62,
    14893 => 62,
    14894 => 62,
    14895 => 62,
    14896 => 62,
    14897 => 62,
    14898 => 62,
    14899 => 62,
    14900 => 62,
    14901 => 62,
    14902 => 62,
    14903 => 62,
    14904 => 62,
    14905 => 62,
    14906 => 62,
    14907 => 62,
    14908 => 62,
    14909 => 62,
    14910 => 62,
    14911 => 62,
    14912 => 62,
    14913 => 62,
    14914 => 62,
    14915 => 62,
    14916 => 62,
    14917 => 62,
    14918 => 62,
    14919 => 62,
    14920 => 62,
    14921 => 62,
    14922 => 62,
    14923 => 62,
    14924 => 62,
    14925 => 62,
    14926 => 62,
    14927 => 62,
    14928 => 62,
    14929 => 62,
    14930 => 62,
    14931 => 62,
    14932 => 62,
    14933 => 62,
    14934 => 62,
    14935 => 62,
    14936 => 62,
    14937 => 62,
    14938 => 62,
    14939 => 62,
    14940 => 62,
    14941 => 62,
    14942 => 62,
    14943 => 62,
    14944 => 62,
    14945 => 62,
    14946 => 62,
    14947 => 62,
    14948 => 62,
    14949 => 62,
    14950 => 62,
    14951 => 62,
    14952 => 62,
    14953 => 62,
    14954 => 62,
    14955 => 62,
    14956 => 62,
    14957 => 62,
    14958 => 62,
    14959 => 62,
    14960 => 62,
    14961 => 62,
    14962 => 62,
    14963 => 62,
    14964 => 62,
    14965 => 62,
    14966 => 62,
    14967 => 62,
    14968 => 62,
    14969 => 62,
    14970 => 62,
    14971 => 62,
    14972 => 62,
    14973 => 62,
    14974 => 62,
    14975 => 62,
    14976 => 62,
    14977 => 62,
    14978 => 62,
    14979 => 62,
    14980 => 62,
    14981 => 62,
    14982 => 62,
    14983 => 62,
    14984 => 62,
    14985 => 62,
    14986 => 62,
    14987 => 62,
    14988 => 62,
    14989 => 62,
    14990 => 62,
    14991 => 62,
    14992 => 62,
    14993 => 62,
    14994 => 62,
    14995 => 62,
    14996 => 62,
    14997 => 62,
    14998 => 62,
    14999 => 62,
    15000 => 62,
    15001 => 62,
    15002 => 62,
    15003 => 62,
    15004 => 62,
    15005 => 62,
    15006 => 62,
    15007 => 62,
    15008 => 62,
    15009 => 62,
    15010 => 62,
    15011 => 62,
    15012 => 62,
    15013 => 62,
    15014 => 62,
    15015 => 62,
    15016 => 62,
    15017 => 62,
    15018 => 62,
    15019 => 62,
    15020 => 62,
    15021 => 62,
    15022 => 62,
    15023 => 62,
    15024 => 62,
    15025 => 62,
    15026 => 62,
    15027 => 62,
    15028 => 62,
    15029 => 62,
    15030 => 62,
    15031 => 62,
    15032 => 62,
    15033 => 62,
    15034 => 62,
    15035 => 62,
    15036 => 62,
    15037 => 62,
    15038 => 62,
    15039 => 62,
    15040 => 62,
    15041 => 62,
    15042 => 62,
    15043 => 62,
    15044 => 62,
    15045 => 62,
    15046 => 62,
    15047 => 62,
    15048 => 62,
    15049 => 62,
    15050 => 62,
    15051 => 62,
    15052 => 62,
    15053 => 62,
    15054 => 62,
    15055 => 62,
    15056 => 62,
    15057 => 62,
    15058 => 62,
    15059 => 62,
    15060 => 62,
    15061 => 62,
    15062 => 62,
    15063 => 62,
    15064 => 62,
    15065 => 62,
    15066 => 62,
    15067 => 62,
    15068 => 62,
    15069 => 62,
    15070 => 63,
    15071 => 63,
    15072 => 63,
    15073 => 63,
    15074 => 63,
    15075 => 63,
    15076 => 63,
    15077 => 63,
    15078 => 63,
    15079 => 63,
    15080 => 63,
    15081 => 63,
    15082 => 63,
    15083 => 63,
    15084 => 63,
    15085 => 63,
    15086 => 63,
    15087 => 63,
    15088 => 63,
    15089 => 63,
    15090 => 63,
    15091 => 63,
    15092 => 63,
    15093 => 63,
    15094 => 63,
    15095 => 63,
    15096 => 63,
    15097 => 63,
    15098 => 63,
    15099 => 63,
    15100 => 63,
    15101 => 63,
    15102 => 63,
    15103 => 63,
    15104 => 63,
    15105 => 63,
    15106 => 63,
    15107 => 63,
    15108 => 63,
    15109 => 63,
    15110 => 63,
    15111 => 63,
    15112 => 63,
    15113 => 63,
    15114 => 63,
    15115 => 63,
    15116 => 63,
    15117 => 63,
    15118 => 63,
    15119 => 63,
    15120 => 63,
    15121 => 63,
    15122 => 63,
    15123 => 63,
    15124 => 63,
    15125 => 63,
    15126 => 63,
    15127 => 63,
    15128 => 63,
    15129 => 63,
    15130 => 63,
    15131 => 63,
    15132 => 63,
    15133 => 63,
    15134 => 63,
    15135 => 63,
    15136 => 63,
    15137 => 63,
    15138 => 63,
    15139 => 63,
    15140 => 63,
    15141 => 63,
    15142 => 63,
    15143 => 63,
    15144 => 63,
    15145 => 63,
    15146 => 63,
    15147 => 63,
    15148 => 63,
    15149 => 63,
    15150 => 63,
    15151 => 63,
    15152 => 63,
    15153 => 63,
    15154 => 63,
    15155 => 63,
    15156 => 63,
    15157 => 63,
    15158 => 63,
    15159 => 63,
    15160 => 63,
    15161 => 63,
    15162 => 63,
    15163 => 63,
    15164 => 63,
    15165 => 63,
    15166 => 63,
    15167 => 63,
    15168 => 63,
    15169 => 63,
    15170 => 63,
    15171 => 63,
    15172 => 63,
    15173 => 63,
    15174 => 63,
    15175 => 63,
    15176 => 63,
    15177 => 63,
    15178 => 63,
    15179 => 63,
    15180 => 63,
    15181 => 63,
    15182 => 63,
    15183 => 63,
    15184 => 63,
    15185 => 63,
    15186 => 63,
    15187 => 63,
    15188 => 63,
    15189 => 63,
    15190 => 63,
    15191 => 63,
    15192 => 63,
    15193 => 63,
    15194 => 63,
    15195 => 63,
    15196 => 63,
    15197 => 63,
    15198 => 63,
    15199 => 63,
    15200 => 63,
    15201 => 63,
    15202 => 63,
    15203 => 63,
    15204 => 63,
    15205 => 63,
    15206 => 63,
    15207 => 63,
    15208 => 63,
    15209 => 63,
    15210 => 63,
    15211 => 63,
    15212 => 63,
    15213 => 63,
    15214 => 63,
    15215 => 63,
    15216 => 63,
    15217 => 63,
    15218 => 63,
    15219 => 63,
    15220 => 63,
    15221 => 63,
    15222 => 63,
    15223 => 63,
    15224 => 63,
    15225 => 63,
    15226 => 63,
    15227 => 63,
    15228 => 63,
    15229 => 63,
    15230 => 63,
    15231 => 63,
    15232 => 63,
    15233 => 63,
    15234 => 63,
    15235 => 63,
    15236 => 63,
    15237 => 63,
    15238 => 63,
    15239 => 63,
    15240 => 63,
    15241 => 63,
    15242 => 63,
    15243 => 63,
    15244 => 63,
    15245 => 63,
    15246 => 63,
    15247 => 63,
    15248 => 63,
    15249 => 63,
    15250 => 63,
    15251 => 63,
    15252 => 63,
    15253 => 63,
    15254 => 63,
    15255 => 63,
    15256 => 63,
    15257 => 63,
    15258 => 63,
    15259 => 63,
    15260 => 63,
    15261 => 63,
    15262 => 63,
    15263 => 63,
    15264 => 63,
    15265 => 63,
    15266 => 63,
    15267 => 63,
    15268 => 63,
    15269 => 63,
    15270 => 63,
    15271 => 63,
    15272 => 63,
    15273 => 63,
    15274 => 63,
    15275 => 63,
    15276 => 63,
    15277 => 63,
    15278 => 63,
    15279 => 63,
    15280 => 63,
    15281 => 63,
    15282 => 63,
    15283 => 63,
    15284 => 63,
    15285 => 63,
    15286 => 63,
    15287 => 63,
    15288 => 63,
    15289 => 63,
    15290 => 63,
    15291 => 63,
    15292 => 63,
    15293 => 63,
    15294 => 63,
    15295 => 63,
    15296 => 63,
    15297 => 63,
    15298 => 63,
    15299 => 63,
    15300 => 63,
    15301 => 63,
    15302 => 63,
    15303 => 63,
    15304 => 63,
    15305 => 63,
    15306 => 63,
    15307 => 63,
    15308 => 63,
    15309 => 63,
    15310 => 63,
    15311 => 63,
    15312 => 63,
    15313 => 63,
    15314 => 63,
    15315 => 63,
    15316 => 63,
    15317 => 63,
    15318 => 63,
    15319 => 63,
    15320 => 63,
    15321 => 63,
    15322 => 63,
    15323 => 63,
    15324 => 63,
    15325 => 63,
    15326 => 63,
    15327 => 63,
    15328 => 63,
    15329 => 63,
    15330 => 63,
    15331 => 63,
    15332 => 63,
    15333 => 63,
    15334 => 63,
    15335 => 63,
    15336 => 63,
    15337 => 63,
    15338 => 63,
    15339 => 63,
    15340 => 63,
    15341 => 63,
    15342 => 63,
    15343 => 63,
    15344 => 63,
    15345 => 63,
    15346 => 63,
    15347 => 63,
    15348 => 63,
    15349 => 63,
    15350 => 63,
    15351 => 63,
    15352 => 63,
    15353 => 63,
    15354 => 63,
    15355 => 63,
    15356 => 63,
    15357 => 63,
    15358 => 63,
    15359 => 63,
    15360 => 63,
    15361 => 63,
    15362 => 63,
    15363 => 63,
    15364 => 63,
    15365 => 63,
    15366 => 63,
    15367 => 63,
    15368 => 63,
    15369 => 63,
    15370 => 63,
    15371 => 63,
    15372 => 63,
    15373 => 63,
    15374 => 63,
    15375 => 63,
    15376 => 63,
    15377 => 63,
    15378 => 63,
    15379 => 63,
    15380 => 63,
    15381 => 63,
    15382 => 63,
    15383 => 63,
    15384 => 63,
    15385 => 63,
    15386 => 63,
    15387 => 63,
    15388 => 63,
    15389 => 63,
    15390 => 63,
    15391 => 63,
    15392 => 63,
    15393 => 63,
    15394 => 63,
    15395 => 63,
    15396 => 63,
    15397 => 63,
    15398 => 63,
    15399 => 63,
    15400 => 63,
    15401 => 63,
    15402 => 63,
    15403 => 63,
    15404 => 63,
    15405 => 63,
    15406 => 63,
    15407 => 63,
    15408 => 63,
    15409 => 63,
    15410 => 63,
    15411 => 63,
    15412 => 63,
    15413 => 63,
    15414 => 63,
    15415 => 63,
    15416 => 63,
    15417 => 63,
    15418 => 63,
    15419 => 63,
    15420 => 63,
    15421 => 63,
    15422 => 63,
    15423 => 63,
    15424 => 63,
    15425 => 63,
    15426 => 63,
    15427 => 63,
    15428 => 63,
    15429 => 63,
    15430 => 63,
    15431 => 63,
    15432 => 63,
    15433 => 63,
    15434 => 63,
    15435 => 63,
    15436 => 63,
    15437 => 63,
    15438 => 63,
    15439 => 63,
    15440 => 63,
    15441 => 63,
    15442 => 63,
    15443 => 63,
    15444 => 63,
    15445 => 63,
    15446 => 63,
    15447 => 63,
    15448 => 63,
    15449 => 63,
    15450 => 63,
    15451 => 63,
    15452 => 63,
    15453 => 63,
    15454 => 63,
    15455 => 63,
    15456 => 63,
    15457 => 63,
    15458 => 63,
    15459 => 63,
    15460 => 63,
    15461 => 63,
    15462 => 63,
    15463 => 63,
    15464 => 63,
    15465 => 63,
    15466 => 63,
    15467 => 63,
    15468 => 63,
    15469 => 63,
    15470 => 63,
    15471 => 63,
    15472 => 63,
    15473 => 63,
    15474 => 63,
    15475 => 63,
    15476 => 63,
    15477 => 63,
    15478 => 63,
    15479 => 63,
    15480 => 63,
    15481 => 63,
    15482 => 63,
    15483 => 63,
    15484 => 63,
    15485 => 63,
    15486 => 63,
    15487 => 63,
    15488 => 63,
    15489 => 63,
    15490 => 63,
    15491 => 63,
    15492 => 63,
    15493 => 63,
    15494 => 63,
    15495 => 63,
    15496 => 63,
    15497 => 63,
    15498 => 63,
    15499 => 63,
    15500 => 63,
    15501 => 63,
    15502 => 63,
    15503 => 63,
    15504 => 63,
    15505 => 63,
    15506 => 63,
    15507 => 63,
    15508 => 63,
    15509 => 63,
    15510 => 63,
    15511 => 63,
    15512 => 63,
    15513 => 63,
    15514 => 63,
    15515 => 63,
    15516 => 63,
    15517 => 63,
    15518 => 63,
    15519 => 63,
    15520 => 63,
    15521 => 63,
    15522 => 63,
    15523 => 63,
    15524 => 63,
    15525 => 63,
    15526 => 63,
    15527 => 63,
    15528 => 63,
    15529 => 63,
    15530 => 63,
    15531 => 63,
    15532 => 63,
    15533 => 63,
    15534 => 63,
    15535 => 63,
    15536 => 63,
    15537 => 63,
    15538 => 63,
    15539 => 63,
    15540 => 63,
    15541 => 63,
    15542 => 63,
    15543 => 63,
    15544 => 63,
    15545 => 63,
    15546 => 63,
    15547 => 63,
    15548 => 63,
    15549 => 63,
    15550 => 63,
    15551 => 63,
    15552 => 63,
    15553 => 63,
    15554 => 63,
    15555 => 63,
    15556 => 63,
    15557 => 63,
    15558 => 63,
    15559 => 63,
    15560 => 63,
    15561 => 63,
    15562 => 63,
    15563 => 63,
    15564 => 63,
    15565 => 63,
    15566 => 63,
    15567 => 63,
    15568 => 63,
    15569 => 63,
    15570 => 63,
    15571 => 63,
    15572 => 63,
    15573 => 63,
    15574 => 63,
    15575 => 63,
    15576 => 63,
    15577 => 63,
    15578 => 63,
    15579 => 63,
    15580 => 63,
    15581 => 63,
    15582 => 63,
    15583 => 63,
    15584 => 63,
    15585 => 63,
    15586 => 63,
    15587 => 63,
    15588 => 63,
    15589 => 63,
    15590 => 63,
    15591 => 63,
    15592 => 63,
    15593 => 63,
    15594 => 63,
    15595 => 63,
    15596 => 63,
    15597 => 63,
    15598 => 63,
    15599 => 63,
    15600 => 63,
    15601 => 63,
    15602 => 63,
    15603 => 63,
    15604 => 63,
    15605 => 63,
    15606 => 63,
    15607 => 63,
    15608 => 63,
    15609 => 63,
    15610 => 63,
    15611 => 63,
    15612 => 63,
    15613 => 63,
    15614 => 63,
    15615 => 63,
    15616 => 63,
    15617 => 63,
    15618 => 63,
    15619 => 63,
    15620 => 63,
    15621 => 63,
    15622 => 63,
    15623 => 63,
    15624 => 63,
    15625 => 63,
    15626 => 63,
    15627 => 63,
    15628 => 63,
    15629 => 63,
    15630 => 63,
    15631 => 63,
    15632 => 63,
    15633 => 63,
    15634 => 63,
    15635 => 63,
    15636 => 63,
    15637 => 63,
    15638 => 63,
    15639 => 63,
    15640 => 63,
    15641 => 63,
    15642 => 63,
    15643 => 63,
    15644 => 63,
    15645 => 63,
    15646 => 63,
    15647 => 63,
    15648 => 63,
    15649 => 63,
    15650 => 63,
    15651 => 63,
    15652 => 63,
    15653 => 63,
    15654 => 63,
    15655 => 63,
    15656 => 63,
    15657 => 63,
    15658 => 63,
    15659 => 63,
    15660 => 63,
    15661 => 63,
    15662 => 63,
    15663 => 63,
    15664 => 63,
    15665 => 63,
    15666 => 63,
    15667 => 63,
    15668 => 63,
    15669 => 63,
    15670 => 63,
    15671 => 63,
    15672 => 63,
    15673 => 63,
    15674 => 63,
    15675 => 63,
    15676 => 63,
    15677 => 63,
    15678 => 63,
    15679 => 63,
    15680 => 63,
    15681 => 63,
    15682 => 63,
    15683 => 63,
    15684 => 63,
    15685 => 63,
    15686 => 63,
    15687 => 63,
    15688 => 63,
    15689 => 63,
    15690 => 63,
    15691 => 63,
    15692 => 63,
    15693 => 63,
    15694 => 63,
    15695 => 63,
    15696 => 63,
    15697 => 63,
    15698 => 63,
    15699 => 63,
    15700 => 63,
    15701 => 63,
    15702 => 63,
    15703 => 63,
    15704 => 63,
    15705 => 63,
    15706 => 63,
    15707 => 63,
    15708 => 63,
    15709 => 63,
    15710 => 63,
    15711 => 63,
    15712 => 63,
    15713 => 63,
    15714 => 63,
    15715 => 63,
    15716 => 63,
    15717 => 63,
    15718 => 63,
    15719 => 63,
    15720 => 63,
    15721 => 63,
    15722 => 63,
    15723 => 63,
    15724 => 63,
    15725 => 63,
    15726 => 63,
    15727 => 63,
    15728 => 63,
    15729 => 63,
    15730 => 63,
    15731 => 63,
    15732 => 63,
    15733 => 63,
    15734 => 63,
    15735 => 63,
    15736 => 63,
    15737 => 63,
    15738 => 63,
    15739 => 63,
    15740 => 63,
    15741 => 63,
    15742 => 63,
    15743 => 63,
    15744 => 63,
    15745 => 63,
    15746 => 63,
    15747 => 63,
    15748 => 63,
    15749 => 63,
    15750 => 63,
    15751 => 63,
    15752 => 63,
    15753 => 63,
    15754 => 63,
    15755 => 63,
    15756 => 63,
    15757 => 63,
    15758 => 63,
    15759 => 63,
    15760 => 63,
    15761 => 63,
    15762 => 63,
    15763 => 63,
    15764 => 63,
    15765 => 63,
    15766 => 63,
    15767 => 63,
    15768 => 63,
    15769 => 63,
    15770 => 63,
    15771 => 63,
    15772 => 63,
    15773 => 63,
    15774 => 63,
    15775 => 63,
    15776 => 63,
    15777 => 63,
    15778 => 63,
    15779 => 63,
    15780 => 63,
    15781 => 63,
    15782 => 63,
    15783 => 63,
    15784 => 63,
    15785 => 63,
    15786 => 63,
    15787 => 63,
    15788 => 63,
    15789 => 63,
    15790 => 63,
    15791 => 63,
    15792 => 63,
    15793 => 63,
    15794 => 63,
    15795 => 63,
    15796 => 63,
    15797 => 63,
    15798 => 63,
    15799 => 63,
    15800 => 63,
    15801 => 63,
    15802 => 63,
    15803 => 63,
    15804 => 63,
    15805 => 63,
    15806 => 63,
    15807 => 63,
    15808 => 63,
    15809 => 63,
    15810 => 63,
    15811 => 63,
    15812 => 63,
    15813 => 63,
    15814 => 63,
    15815 => 63,
    15816 => 63,
    15817 => 63,
    15818 => 63,
    15819 => 63,
    15820 => 63,
    15821 => 63,
    15822 => 63,
    15823 => 63,
    15824 => 63,
    15825 => 63,
    15826 => 63,
    15827 => 63,
    15828 => 63,
    15829 => 63,
    15830 => 63,
    15831 => 63,
    15832 => 63,
    15833 => 63,
    15834 => 63,
    15835 => 63,
    15836 => 63,
    15837 => 63,
    15838 => 63,
    15839 => 63,
    15840 => 63,
    15841 => 63,
    15842 => 63,
    15843 => 63,
    15844 => 63,
    15845 => 63,
    15846 => 63,
    15847 => 63,
    15848 => 63,
    15849 => 63,
    15850 => 63,
    15851 => 63,
    15852 => 63,
    15853 => 63,
    15854 => 63,
    15855 => 63,
    15856 => 63,
    15857 => 63,
    15858 => 63,
    15859 => 63,
    15860 => 63,
    15861 => 63,
    15862 => 63,
    15863 => 63,
    15864 => 63,
    15865 => 63,
    15866 => 63,
    15867 => 63,
    15868 => 63,
    15869 => 63,
    15870 => 63,
    15871 => 63,
    15872 => 63,
    15873 => 63,
    15874 => 63,
    15875 => 63,
    15876 => 63,
    15877 => 63,
    15878 => 63,
    15879 => 63,
    15880 => 63,
    15881 => 63,
    15882 => 63,
    15883 => 63,
    15884 => 63,
    15885 => 63,
    15886 => 63,
    15887 => 63,
    15888 => 63,
    15889 => 63,
    15890 => 63,
    15891 => 63,
    15892 => 63,
    15893 => 63,
    15894 => 63,
    15895 => 63,
    15896 => 63,
    15897 => 63,
    15898 => 63,
    15899 => 63,
    15900 => 63,
    15901 => 63,
    15902 => 63,
    15903 => 63,
    15904 => 63,
    15905 => 63,
    15906 => 63,
    15907 => 63,
    15908 => 63,
    15909 => 63,
    15910 => 63,
    15911 => 63,
    15912 => 63,
    15913 => 63,
    15914 => 63,
    15915 => 63,
    15916 => 63,
    15917 => 63,
    15918 => 63,
    15919 => 63,
    15920 => 63,
    15921 => 63,
    15922 => 63,
    15923 => 63,
    15924 => 63,
    15925 => 63,
    15926 => 63,
    15927 => 63,
    15928 => 63,
    15929 => 63,
    15930 => 63,
    15931 => 63,
    15932 => 63,
    15933 => 63,
    15934 => 63,
    15935 => 63,
    15936 => 63,
    15937 => 63,
    15938 => 63,
    15939 => 63,
    15940 => 63,
    15941 => 63,
    15942 => 63,
    15943 => 63,
    15944 => 63,
    15945 => 63,
    15946 => 63,
    15947 => 63,
    15948 => 63,
    15949 => 63,
    15950 => 63,
    15951 => 63,
    15952 => 63,
    15953 => 63,
    15954 => 63,
    15955 => 63,
    15956 => 63,
    15957 => 63,
    15958 => 63,
    15959 => 63,
    15960 => 63,
    15961 => 63,
    15962 => 63,
    15963 => 63,
    15964 => 63,
    15965 => 63,
    15966 => 63,
    15967 => 63,
    15968 => 63,
    15969 => 63,
    15970 => 63,
    15971 => 63,
    15972 => 63,
    15973 => 63,
    15974 => 63,
    15975 => 63,
    15976 => 63,
    15977 => 63,
    15978 => 63,
    15979 => 63,
    15980 => 63,
    15981 => 63,
    15982 => 63,
    15983 => 63,
    15984 => 63,
    15985 => 63,
    15986 => 63,
    15987 => 63,
    15988 => 63,
    15989 => 63,
    15990 => 63,
    15991 => 63,
    15992 => 63,
    15993 => 63,
    15994 => 63,
    15995 => 63,
    15996 => 63,
    15997 => 63,
    15998 => 63,
    15999 => 63,
    16000 => 63,
    16001 => 63,
    16002 => 63,
    16003 => 63,
    16004 => 63,
    16005 => 63,
    16006 => 63,
    16007 => 63,
    16008 => 63,
    16009 => 63,
    16010 => 63,
    16011 => 63,
    16012 => 63,
    16013 => 63,
    16014 => 63,
    16015 => 63,
    16016 => 63,
    16017 => 63,
    16018 => 63,
    16019 => 63,
    16020 => 63,
    16021 => 63,
    16022 => 63,
    16023 => 63,
    16024 => 63,
    16025 => 63,
    16026 => 63,
    16027 => 63,
    16028 => 63,
    16029 => 63,
    16030 => 63,
    16031 => 63,
    16032 => 63,
    16033 => 63,
    16034 => 63,
    16035 => 63,
    16036 => 63,
    16037 => 63,
    16038 => 63,
    16039 => 63,
    16040 => 63,
    16041 => 63,
    16042 => 63,
    16043 => 63,
    16044 => 63,
    16045 => 63,
    16046 => 63,
    16047 => 63,
    16048 => 63,
    16049 => 63,
    16050 => 63,
    16051 => 63,
    16052 => 63,
    16053 => 63,
    16054 => 63,
    16055 => 63,
    16056 => 63,
    16057 => 63,
    16058 => 63,
    16059 => 63,
    16060 => 63,
    16061 => 63,
    16062 => 63,
    16063 => 63,
    16064 => 63,
    16065 => 63,
    16066 => 63,
    16067 => 63,
    16068 => 63,
    16069 => 63,
    16070 => 63,
    16071 => 63,
    16072 => 63,
    16073 => 63,
    16074 => 63,
    16075 => 63,
    16076 => 63,
    16077 => 63,
    16078 => 63,
    16079 => 63,
    16080 => 63,
    16081 => 63,
    16082 => 63,
    16083 => 63,
    16084 => 63,
    16085 => 63,
    16086 => 63,
    16087 => 63,
    16088 => 63,
    16089 => 63,
    16090 => 63,
    16091 => 63,
    16092 => 63,
    16093 => 63,
    16094 => 63,
    16095 => 63,
    16096 => 63,
    16097 => 63,
    16098 => 63,
    16099 => 63,
    16100 => 63,
    16101 => 63,
    16102 => 63,
    16103 => 63,
    16104 => 63,
    16105 => 63,
    16106 => 63,
    16107 => 63,
    16108 => 63,
    16109 => 63,
    16110 => 63,
    16111 => 63,
    16112 => 63,
    16113 => 63,
    16114 => 63,
    16115 => 63,
    16116 => 63,
    16117 => 63,
    16118 => 63,
    16119 => 63,
    16120 => 63,
    16121 => 63,
    16122 => 63,
    16123 => 63,
    16124 => 63,
    16125 => 63,
    16126 => 63,
    16127 => 63,
    16128 => 63,
    16129 => 63,
    16130 => 63,
    16131 => 63,
    16132 => 63,
    16133 => 63,
    16134 => 63,
    16135 => 63,
    16136 => 63,
    16137 => 63,
    16138 => 63,
    16139 => 63,
    16140 => 63,
    16141 => 63,
    16142 => 63,
    16143 => 63,
    16144 => 63,
    16145 => 63,
    16146 => 63,
    16147 => 63,
    16148 => 63,
    16149 => 63,
    16150 => 63,
    16151 => 63,
    16152 => 63,
    16153 => 63,
    16154 => 63,
    16155 => 63,
    16156 => 63,
    16157 => 63,
    16158 => 63,
    16159 => 63,
    16160 => 63,
    16161 => 63,
    16162 => 63,
    16163 => 63,
    16164 => 63,
    16165 => 63,
    16166 => 63,
    16167 => 63,
    16168 => 63,
    16169 => 63,
    16170 => 63,
    16171 => 63,
    16172 => 63,
    16173 => 63,
    16174 => 63,
    16175 => 63,
    16176 => 63,
    16177 => 63,
    16178 => 63,
    16179 => 63,
    16180 => 63,
    16181 => 63,
    16182 => 63,
    16183 => 63,
    16184 => 63,
    16185 => 63,
    16186 => 63,
    16187 => 63,
    16188 => 63,
    16189 => 63,
    16190 => 63,
    16191 => 63,
    16192 => 63,
    16193 => 63,
    16194 => 63,
    16195 => 63,
    16196 => 63,
    16197 => 63,
    16198 => 63,
    16199 => 63,
    16200 => 63,
    16201 => 63,
    16202 => 63,
    16203 => 63,
    16204 => 63,
    16205 => 63,
    16206 => 63,
    16207 => 63,
    16208 => 63,
    16209 => 63,
    16210 => 63,
    16211 => 63,
    16212 => 63,
    16213 => 63,
    16214 => 63,
    16215 => 63,
    16216 => 63,
    16217 => 63,
    16218 => 63,
    16219 => 63,
    16220 => 63,
    16221 => 63,
    16222 => 63,
    16223 => 63,
    16224 => 63,
    16225 => 63,
    16226 => 63,
    16227 => 63,
    16228 => 63,
    16229 => 63,
    16230 => 63,
    16231 => 63,
    16232 => 63,
    16233 => 63,
    16234 => 63,
    16235 => 63,
    16236 => 63,
    16237 => 63,
    16238 => 63,
    16239 => 63,
    16240 => 63,
    16241 => 63,
    16242 => 63,
    16243 => 63,
    16244 => 63,
    16245 => 63,
    16246 => 63,
    16247 => 63,
    16248 => 63,
    16249 => 63,
    16250 => 63,
    16251 => 63,
    16252 => 63,
    16253 => 63,
    16254 => 63,
    16255 => 63,
    16256 => 63,
    16257 => 63,
    16258 => 63,
    16259 => 63,
    16260 => 63,
    16261 => 63,
    16262 => 63,
    16263 => 63,
    16264 => 63,
    16265 => 63,
    16266 => 63,
    16267 => 63,
    16268 => 63,
    16269 => 63,
    16270 => 63,
    16271 => 63,
    16272 => 63,
    16273 => 63,
    16274 => 63,
    16275 => 63,
    16276 => 63,
    16277 => 63,
    16278 => 63,
    16279 => 63,
    16280 => 63,
    16281 => 63,
    16282 => 63,
    16283 => 63,
    16284 => 63,
    16285 => 63,
    16286 => 63,
    16287 => 63,
    16288 => 63,
    16289 => 63,
    16290 => 63,
    16291 => 63,
    16292 => 63,
    16293 => 63,
    16294 => 63,
    16295 => 63,
    16296 => 63,
    16297 => 63,
    16298 => 63,
    16299 => 63,
    16300 => 63,
    16301 => 63,
    16302 => 63,
    16303 => 63,
    16304 => 63,
    16305 => 63,
    16306 => 63,
    16307 => 63,
    16308 => 63,
    16309 => 63,
    16310 => 63,
    16311 => 63,
    16312 => 63,
    16313 => 63,
    16314 => 63,
    16315 => 63,
    16316 => 63,
    16317 => 63,
    16318 => 63,
    16319 => 63,
    16320 => 63,
    16321 => 63,
    16322 => 63,
    16323 => 63,
    16324 => 63,
    16325 => 63,
    16326 => 63,
    16327 => 63,
    16328 => 63,
    16329 => 63,
    16330 => 63,
    16331 => 63,
    16332 => 63,
    16333 => 63,
    16334 => 63,
    16335 => 63,
    16336 => 63,
    16337 => 63,
    16338 => 63,
    16339 => 63,
    16340 => 63,
    16341 => 63,
    16342 => 63,
    16343 => 63,
    16344 => 63,
    16345 => 63,
    16346 => 63,
    16347 => 63,
    16348 => 63,
    16349 => 63,
    16350 => 63,
    16351 => 63,
    16352 => 63,
    16353 => 63,
    16354 => 63,
    16355 => 63,
    16356 => 63,
    16357 => 63,
    16358 => 63,
    16359 => 63,
    16360 => 63,
    16361 => 63,
    16362 => 63,
    16363 => 63,
    16364 => 63,
    16365 => 63,
    16366 => 63,
    16367 => 63,
    16368 => 63,
    16369 => 63,
    16370 => 63,
    16371 => 63,
    16372 => 63,
    16373 => 63,
    16374 => 63,
    16375 => 63,
    16376 => 63,
    16377 => 63,
    16378 => 63,
    16379 => 63,
    16380 => 63,
    16381 => 63,
    16382 => 63,
    16383 => 63,
    16384 => 63,
    16385 => 63,
    16386 => 63,
    16387 => 63,
    16388 => 63,
    16389 => 63,
    16390 => 63,
    16391 => 63,
    16392 => 63,
    16393 => 63,
    16394 => 63,
    16395 => 63,
    16396 => 63,
    16397 => 63,
    16398 => 63,
    16399 => 63,
    16400 => 63,
    16401 => 63,
    16402 => 63,
    16403 => 63,
    16404 => 63,
    16405 => 63,
    16406 => 63,
    16407 => 63,
    16408 => 63,
    16409 => 63,
    16410 => 63,
    16411 => 63,
    16412 => 63,
    16413 => 63,
    16414 => 63,
    16415 => 63,
    16416 => 63,
    16417 => 63,
    16418 => 63,
    16419 => 63,
    16420 => 63,
    16421 => 63,
    16422 => 63,
    16423 => 63,
    16424 => 63,
    16425 => 63,
    16426 => 63,
    16427 => 63,
    16428 => 63,
    16429 => 63,
    16430 => 63,
    16431 => 63,
    16432 => 63,
    16433 => 63,
    16434 => 63,
    16435 => 63,
    16436 => 63,
    16437 => 63,
    16438 => 63,
    16439 => 63,
    16440 => 63,
    16441 => 63,
    16442 => 63,
    16443 => 63,
    16444 => 63,
    16445 => 63,
    16446 => 63,
    16447 => 63,
    16448 => 63,
    16449 => 63,
    16450 => 63,
    16451 => 63,
    16452 => 63,
    16453 => 63,
    16454 => 63,
    16455 => 63,
    16456 => 63,
    16457 => 63,
    16458 => 63,
    16459 => 63,
    16460 => 63,
    16461 => 63,
    16462 => 63,
    16463 => 63,
    16464 => 63,
    16465 => 63,
    16466 => 63,
    16467 => 63,
    16468 => 63,
    16469 => 63,
    16470 => 63,
    16471 => 63,
    16472 => 63,
    16473 => 63,
    16474 => 63,
    16475 => 63,
    16476 => 63,
    16477 => 63,
    16478 => 63,
    16479 => 63,
    16480 => 63,
    16481 => 63,
    16482 => 63,
    16483 => 63,
    16484 => 63,
    16485 => 63,
    16486 => 63,
    16487 => 63,
    16488 => 63,
    16489 => 63,
    16490 => 63,
    16491 => 63,
    16492 => 63,
    16493 => 63,
    16494 => 63,
    16495 => 63,
    16496 => 63,
    16497 => 63,
    16498 => 63,
    16499 => 63,
    16500 => 63,
    16501 => 63,
    16502 => 63,
    16503 => 63,
    16504 => 63,
    16505 => 63,
    16506 => 63,
    16507 => 63,
    16508 => 63,
    16509 => 63,
    16510 => 63,
    16511 => 63,
    16512 => 63,
    16513 => 63,
    16514 => 63,
    16515 => 63,
    16516 => 63,
    16517 => 63,
    16518 => 63,
    16519 => 63,
    16520 => 63,
    16521 => 63,
    16522 => 63,
    16523 => 63,
    16524 => 63,
    16525 => 63,
    16526 => 63,
    16527 => 63,
    16528 => 63,
    16529 => 63,
    16530 => 63,
    16531 => 63,
    16532 => 63,
    16533 => 63,
    16534 => 63,
    16535 => 63,
    16536 => 63,
    16537 => 63,
    16538 => 63,
    16539 => 63,
    16540 => 63,
    16541 => 63,
    16542 => 63,
    16543 => 63,
    16544 => 63,
    16545 => 63,
    16546 => 63,
    16547 => 63,
    16548 => 63,
    16549 => 63,
    16550 => 63,
    16551 => 63,
    16552 => 63,
    16553 => 63,
    16554 => 63,
    16555 => 63,
    16556 => 63,
    16557 => 63,
    16558 => 63,
    16559 => 63,
    16560 => 63,
    16561 => 63,
    16562 => 63,
    16563 => 63,
    16564 => 63,
    16565 => 63,
    16566 => 63,
    16567 => 63,
    16568 => 63,
    16569 => 63,
    16570 => 63,
    16571 => 63,
    16572 => 63,
    16573 => 63,
    16574 => 63,
    16575 => 63,
    16576 => 63,
    16577 => 63,
    16578 => 63,
    16579 => 63,
    16580 => 63,
    16581 => 63,
    16582 => 63,
    16583 => 63,
    16584 => 63,
    16585 => 63,
    16586 => 63,
    16587 => 63,
    16588 => 63,
    16589 => 63,
    16590 => 63,
    16591 => 63,
    16592 => 63,
    16593 => 63,
    16594 => 63,
    16595 => 63,
    16596 => 63,
    16597 => 63,
    16598 => 63,
    16599 => 63,
    16600 => 63,
    16601 => 63,
    16602 => 63,
    16603 => 63,
    16604 => 63,
    16605 => 63,
    16606 => 63,
    16607 => 63,
    16608 => 63,
    16609 => 63,
    16610 => 63,
    16611 => 63,
    16612 => 63,
    16613 => 63,
    16614 => 63,
    16615 => 63,
    16616 => 63,
    16617 => 63,
    16618 => 63,
    16619 => 63,
    16620 => 63,
    16621 => 63,
    16622 => 63,
    16623 => 63,
    16624 => 63,
    16625 => 63,
    16626 => 63,
    16627 => 63,
    16628 => 63,
    16629 => 63,
    16630 => 63,
    16631 => 63,
    16632 => 63,
    16633 => 63,
    16634 => 63,
    16635 => 63,
    16636 => 63,
    16637 => 63,
    16638 => 63,
    16639 => 63,
    16640 => 63,
    16641 => 63,
    16642 => 63,
    16643 => 63,
    16644 => 63,
    16645 => 63,
    16646 => 63,
    16647 => 63,
    16648 => 63,
    16649 => 63,
    16650 => 63,
    16651 => 63,
    16652 => 63,
    16653 => 63,
    16654 => 63,
    16655 => 63,
    16656 => 63,
    16657 => 63,
    16658 => 63,
    16659 => 63,
    16660 => 63,
    16661 => 63,
    16662 => 63,
    16663 => 63,
    16664 => 63,
    16665 => 63,
    16666 => 63,
    16667 => 63,
    16668 => 63,
    16669 => 63,
    16670 => 63,
    16671 => 63,
    16672 => 63,
    16673 => 63,
    16674 => 63,
    16675 => 63,
    16676 => 63,
    16677 => 63,
    16678 => 63,
    16679 => 63,
    16680 => 63,
    16681 => 63,
    16682 => 63,
    16683 => 63,
    16684 => 63,
    16685 => 63,
    16686 => 63,
    16687 => 63,
    16688 => 63,
    16689 => 63,
    16690 => 63,
    16691 => 63,
    16692 => 63,
    16693 => 63,
    16694 => 63,
    16695 => 63,
    16696 => 63,
    16697 => 63,
    16698 => 63,
    16699 => 63,
    16700 => 63,
    16701 => 63,
    16702 => 63,
    16703 => 63,
    16704 => 63,
    16705 => 63,
    16706 => 63,
    16707 => 63,
    16708 => 63,
    16709 => 63,
    16710 => 63,
    16711 => 63,
    16712 => 63,
    16713 => 63,
    16714 => 63,
    16715 => 63,
    16716 => 63,
    16717 => 63,
    16718 => 63,
    16719 => 63,
    16720 => 63,
    16721 => 63,
    16722 => 63,
    16723 => 63,
    16724 => 63,
    16725 => 63,
    16726 => 63,
    16727 => 63,
    16728 => 63,
    16729 => 63,
    16730 => 63,
    16731 => 63,
    16732 => 63,
    16733 => 63,
    16734 => 63,
    16735 => 63,
    16736 => 63,
    16737 => 63,
    16738 => 63,
    16739 => 63,
    16740 => 63,
    16741 => 63,
    16742 => 63,
    16743 => 63,
    16744 => 63,
    16745 => 63,
    16746 => 63,
    16747 => 63,
    16748 => 63,
    16749 => 63,
    16750 => 63,
    16751 => 63,
    16752 => 63,
    16753 => 63,
    16754 => 63,
    16755 => 63,
    16756 => 63,
    16757 => 63,
    16758 => 63,
    16759 => 63,
    16760 => 63,
    16761 => 63,
    16762 => 63,
    16763 => 63,
    16764 => 63,
    16765 => 63,
    16766 => 63,
    16767 => 63,
    16768 => 63,
    16769 => 63,
    16770 => 63,
    16771 => 63,
    16772 => 63,
    16773 => 63,
    16774 => 63,
    16775 => 63,
    16776 => 63,
    16777 => 63,
    16778 => 63,
    16779 => 63,
    16780 => 63,
    16781 => 63,
    16782 => 63,
    16783 => 63,
    16784 => 63,
    16785 => 63,
    16786 => 63,
    16787 => 63,
    16788 => 63,
    16789 => 63,
    16790 => 63,
    16791 => 63,
    16792 => 63,
    16793 => 63,
    16794 => 63,
    16795 => 63,
    16796 => 63,
    16797 => 63,
    16798 => 63,
    16799 => 63,
    16800 => 63,
    16801 => 63,
    16802 => 63,
    16803 => 63,
    16804 => 63,
    16805 => 63,
    16806 => 63,
    16807 => 63,
    16808 => 63,
    16809 => 63,
    16810 => 63,
    16811 => 63,
    16812 => 63,
    16813 => 63,
    16814 => 63,
    16815 => 63,
    16816 => 63,
    16817 => 63,
    16818 => 63,
    16819 => 63,
    16820 => 63,
    16821 => 63,
    16822 => 63,
    16823 => 63,
    16824 => 63,
    16825 => 63,
    16826 => 63,
    16827 => 63,
    16828 => 63,
    16829 => 63,
    16830 => 63,
    16831 => 63,
    16832 => 63,
    16833 => 63,
    16834 => 63,
    16835 => 63,
    16836 => 63,
    16837 => 63,
    16838 => 63,
    16839 => 63,
    16840 => 63,
    16841 => 63,
    16842 => 63,
    16843 => 63,
    16844 => 63,
    16845 => 63,
    16846 => 63,
    16847 => 63,
    16848 => 63,
    16849 => 63,
    16850 => 63,
    16851 => 63,
    16852 => 63,
    16853 => 63,
    16854 => 63,
    16855 => 63,
    16856 => 63,
    16857 => 63,
    16858 => 63,
    16859 => 63,
    16860 => 63,
    16861 => 63,
    16862 => 63,
    16863 => 63,
    16864 => 63,
    16865 => 63,
    16866 => 63,
    16867 => 63,
    16868 => 63,
    16869 => 63,
    16870 => 63,
    16871 => 63,
    16872 => 63,
    16873 => 63,
    16874 => 63,
    16875 => 63,
    16876 => 63,
    16877 => 63,
    16878 => 63,
    16879 => 63,
    16880 => 63,
    16881 => 63,
    16882 => 63,
    16883 => 63,
    16884 => 63,
    16885 => 63,
    16886 => 63,
    16887 => 63,
    16888 => 63,
    16889 => 63,
    16890 => 63,
    16891 => 63,
    16892 => 63,
    16893 => 63,
    16894 => 63,
    16895 => 63,
    16896 => 63,
    16897 => 63,
    16898 => 63,
    16899 => 63,
    16900 => 63,
    16901 => 63,
    16902 => 63,
    16903 => 63,
    16904 => 63,
    16905 => 63,
    16906 => 63,
    16907 => 63,
    16908 => 63,
    16909 => 63,
    16910 => 63,
    16911 => 63,
    16912 => 63,
    16913 => 63,
    16914 => 63,
    16915 => 63,
    16916 => 63,
    16917 => 63,
    16918 => 63,
    16919 => 63,
    16920 => 63,
    16921 => 63,
    16922 => 63,
    16923 => 63,
    16924 => 63,
    16925 => 63,
    16926 => 63,
    16927 => 63,
    16928 => 63,
    16929 => 63,
    16930 => 63,
    16931 => 63,
    16932 => 63,
    16933 => 63,
    16934 => 63,
    16935 => 63,
    16936 => 63,
    16937 => 63,
    16938 => 63,
    16939 => 63,
    16940 => 63,
    16941 => 63,
    16942 => 63,
    16943 => 63,
    16944 => 63,
    16945 => 63,
    16946 => 63,
    16947 => 63,
    16948 => 63,
    16949 => 63,
    16950 => 63,
    16951 => 63,
    16952 => 63,
    16953 => 63,
    16954 => 63,
    16955 => 63,
    16956 => 63,
    16957 => 63,
    16958 => 63,
    16959 => 63,
    16960 => 63,
    16961 => 63,
    16962 => 63,
    16963 => 63,
    16964 => 63,
    16965 => 63,
    16966 => 63,
    16967 => 63,
    16968 => 63,
    16969 => 63,
    16970 => 63,
    16971 => 63,
    16972 => 63,
    16973 => 63,
    16974 => 63,
    16975 => 63,
    16976 => 63,
    16977 => 63,
    16978 => 63,
    16979 => 63,
    16980 => 63,
    16981 => 63,
    16982 => 63,
    16983 => 63,
    16984 => 63,
    16985 => 63,
    16986 => 63,
    16987 => 63,
    16988 => 63,
    16989 => 63,
    16990 => 63,
    16991 => 63,
    16992 => 63,
    16993 => 63,
    16994 => 63,
    16995 => 63,
    16996 => 63,
    16997 => 63,
    16998 => 63,
    16999 => 63,
    17000 => 63,
    17001 => 63,
    17002 => 63,
    17003 => 63,
    17004 => 63,
    17005 => 63,
    17006 => 63,
    17007 => 63,
    17008 => 63,
    17009 => 63,
    17010 => 63,
    17011 => 63,
    17012 => 63,
    17013 => 63,
    17014 => 63,
    17015 => 63,
    17016 => 63,
    17017 => 63,
    17018 => 63,
    17019 => 63,
    17020 => 63,
    17021 => 63,
    17022 => 63,
    17023 => 63,
    17024 => 63,
    17025 => 63,
    17026 => 63,
    17027 => 63,
    17028 => 63,
    17029 => 63,
    17030 => 63,
    17031 => 63,
    17032 => 63,
    17033 => 63,
    17034 => 63,
    17035 => 63,
    17036 => 63,
    17037 => 63,
    17038 => 63,
    17039 => 63,
    17040 => 63,
    17041 => 63,
    17042 => 63,
    17043 => 63,
    17044 => 63,
    17045 => 63,
    17046 => 63,
    17047 => 63,
    17048 => 63,
    17049 => 63,
    17050 => 63,
    17051 => 63,
    17052 => 63,
    17053 => 63,
    17054 => 63,
    17055 => 63,
    17056 => 63,
    17057 => 63,
    17058 => 63,
    17059 => 63,
    17060 => 63,
    17061 => 63,
    17062 => 63,
    17063 => 63,
    17064 => 63,
    17065 => 63,
    17066 => 63,
    17067 => 63,
    17068 => 63,
    17069 => 63,
    17070 => 63,
    17071 => 63,
    17072 => 63,
    17073 => 63,
    17074 => 63,
    17075 => 63,
    17076 => 63,
    17077 => 63,
    17078 => 63,
    17079 => 63,
    17080 => 63,
    17081 => 63,
    17082 => 63,
    17083 => 63,
    17084 => 63,
    17085 => 63,
    17086 => 63,
    17087 => 63,
    17088 => 63,
    17089 => 63,
    17090 => 63,
    17091 => 63,
    17092 => 63,
    17093 => 63,
    17094 => 63,
    17095 => 63,
    17096 => 63,
    17097 => 63,
    17098 => 63,
    17099 => 63,
    17100 => 63,
    17101 => 63,
    17102 => 63,
    17103 => 63,
    17104 => 63,
    17105 => 63,
    17106 => 63,
    17107 => 63,
    17108 => 63,
    17109 => 63,
    17110 => 63,
    17111 => 63,
    17112 => 63,
    17113 => 63,
    17114 => 63,
    17115 => 63,
    17116 => 63,
    17117 => 63,
    17118 => 63,
    17119 => 63,
    17120 => 63,
    17121 => 63,
    17122 => 63,
    17123 => 63,
    17124 => 63,
    17125 => 63,
    17126 => 63,
    17127 => 63,
    17128 => 63,
    17129 => 63,
    17130 => 63,
    17131 => 63,
    17132 => 63,
    17133 => 63,
    17134 => 63,
    17135 => 63,
    17136 => 63,
    17137 => 63,
    17138 => 63,
    17139 => 63,
    17140 => 63,
    17141 => 63,
    17142 => 63,
    17143 => 63,
    17144 => 63,
    17145 => 63,
    17146 => 63,
    17147 => 63,
    17148 => 63,
    17149 => 63,
    17150 => 63,
    17151 => 63,
    17152 => 63,
    17153 => 63,
    17154 => 63,
    17155 => 63,
    17156 => 63,
    17157 => 63,
    17158 => 63,
    17159 => 63,
    17160 => 63,
    17161 => 63,
    17162 => 63,
    17163 => 63,
    17164 => 63,
    17165 => 63,
    17166 => 63,
    17167 => 63,
    17168 => 63,
    17169 => 63,
    17170 => 63,
    17171 => 63,
    17172 => 63,
    17173 => 63,
    17174 => 63,
    17175 => 63,
    17176 => 63,
    17177 => 63,
    17178 => 63,
    17179 => 63,
    17180 => 63,
    17181 => 63,
    17182 => 63,
    17183 => 63,
    17184 => 63,
    17185 => 63,
    17186 => 63,
    17187 => 63,
    17188 => 63,
    17189 => 63,
    17190 => 63,
    17191 => 63,
    17192 => 63,
    17193 => 63,
    17194 => 63,
    17195 => 63,
    17196 => 63,
    17197 => 63,
    17198 => 63,
    17199 => 63,
    17200 => 63,
    17201 => 63,
    17202 => 63,
    17203 => 63,
    17204 => 63,
    17205 => 63,
    17206 => 63,
    17207 => 63,
    17208 => 63,
    17209 => 63,
    17210 => 63,
    17211 => 63,
    17212 => 63,
    17213 => 63,
    17214 => 63,
    17215 => 63,
    17216 => 63,
    17217 => 63,
    17218 => 63,
    17219 => 63,
    17220 => 63,
    17221 => 63,
    17222 => 63,
    17223 => 63,
    17224 => 63,
    17225 => 63,
    17226 => 63,
    17227 => 63,
    17228 => 63,
    17229 => 63,
    17230 => 63,
    17231 => 63,
    17232 => 63,
    17233 => 63,
    17234 => 63,
    17235 => 63,
    17236 => 63,
    17237 => 63,
    17238 => 63,
    17239 => 63,
    17240 => 63,
    17241 => 63,
    17242 => 63,
    17243 => 63,
    17244 => 63,
    17245 => 63,
    17246 => 63,
    17247 => 63,
    17248 => 63,
    17249 => 63,
    17250 => 63,
    17251 => 63,
    17252 => 63,
    17253 => 63,
    17254 => 63,
    17255 => 63,
    17256 => 63,
    17257 => 63,
    17258 => 63,
    17259 => 63,
    17260 => 63,
    17261 => 63,
    17262 => 63,
    17263 => 63,
    17264 => 63,
    17265 => 63,
    17266 => 63,
    17267 => 63,
    17268 => 63,
    17269 => 63,
    17270 => 63,
    17271 => 63,
    17272 => 63,
    17273 => 63,
    17274 => 63,
    17275 => 63,
    17276 => 63,
    17277 => 63,
    17278 => 63,
    17279 => 63,
    17280 => 63,
    17281 => 63,
    17282 => 63,
    17283 => 63,
    17284 => 63,
    17285 => 63,
    17286 => 63,
    17287 => 63,
    17288 => 63,
    17289 => 63,
    17290 => 63,
    17291 => 63,
    17292 => 63,
    17293 => 63,
    17294 => 63,
    17295 => 63,
    17296 => 63,
    17297 => 63,
    17298 => 63,
    17299 => 63,
    17300 => 63,
    17301 => 63,
    17302 => 63,
    17303 => 63,
    17304 => 63,
    17305 => 63,
    17306 => 63,
    17307 => 63,
    17308 => 63,
    17309 => 63,
    17310 => 63,
    17311 => 63,
    17312 => 63,
    17313 => 63,
    17314 => 63,
    17315 => 63,
    17316 => 63,
    17317 => 63,
    17318 => 63,
    17319 => 63,
    17320 => 63,
    17321 => 63,
    17322 => 63,
    17323 => 63,
    17324 => 63,
    17325 => 63,
    17326 => 63,
    17327 => 63,
    17328 => 63,
    17329 => 63,
    17330 => 63,
    17331 => 63,
    17332 => 63,
    17333 => 63,
    17334 => 63,
    17335 => 63,
    17336 => 63,
    17337 => 63,
    17338 => 63,
    17339 => 63,
    17340 => 63,
    17341 => 63,
    17342 => 63,
    17343 => 63,
    17344 => 63,
    17345 => 63,
    17346 => 63,
    17347 => 63,
    17348 => 63,
    17349 => 63,
    17350 => 63,
    17351 => 63,
    17352 => 63,
    17353 => 63,
    17354 => 63,
    17355 => 63,
    17356 => 63,
    17357 => 63,
    17358 => 63,
    17359 => 63,
    17360 => 63,
    17361 => 63,
    17362 => 63,
    17363 => 63,
    17364 => 63,
    17365 => 63,
    17366 => 63,
    17367 => 63,
    17368 => 63,
    17369 => 63,
    17370 => 63,
    17371 => 63,
    17372 => 63,
    17373 => 63,
    17374 => 63,
    17375 => 63,
    17376 => 63,
    17377 => 63,
    17378 => 63,
    17379 => 63,
    17380 => 63,
    17381 => 63,
    17382 => 63,
    17383 => 63,
    17384 => 63,
    17385 => 63,
    17386 => 63,
    17387 => 63,
    17388 => 63,
    17389 => 63,
    17390 => 63,
    17391 => 63,
    17392 => 63,
    17393 => 63,
    17394 => 63,
    17395 => 63,
    17396 => 63,
    17397 => 63,
    17398 => 63,
    17399 => 63,
    17400 => 63,
    17401 => 63,
    17402 => 63,
    17403 => 63,
    17404 => 63,
    17405 => 63,
    17406 => 63,
    17407 => 63,
    17408 => 63,
    17409 => 63,
    17410 => 63,
    17411 => 63,
    17412 => 63,
    17413 => 63,
    17414 => 63,
    17415 => 63,
    17416 => 63,
    17417 => 63,
    17418 => 63,
    17419 => 63,
    17420 => 63,
    17421 => 63,
    17422 => 63,
    17423 => 63,
    17424 => 63,
    17425 => 63,
    17426 => 63,
    17427 => 63,
    17428 => 63,
    17429 => 63,
    17430 => 63,
    17431 => 63,
    17432 => 63,
    17433 => 63,
    17434 => 63,
    17435 => 63,
    17436 => 63,
    17437 => 63,
    17438 => 63,
    17439 => 63,
    17440 => 63,
    17441 => 63,
    17442 => 63,
    17443 => 63,
    17444 => 63,
    17445 => 63,
    17446 => 63,
    17447 => 63,
    17448 => 63,
    17449 => 63,
    17450 => 63,
    17451 => 63,
    17452 => 63,
    17453 => 63,
    17454 => 63,
    17455 => 63,
    17456 => 63,
    17457 => 63,
    17458 => 63,
    17459 => 63,
    17460 => 63,
    17461 => 63,
    17462 => 63,
    17463 => 63,
    17464 => 63,
    17465 => 63,
    17466 => 63,
    17467 => 63,
    17468 => 63,
    17469 => 63,
    17470 => 63,
    17471 => 63,
    17472 => 63,
    17473 => 63,
    17474 => 63,
    17475 => 63,
    17476 => 63,
    17477 => 63,
    17478 => 63,
    17479 => 63,
    17480 => 63,
    17481 => 63,
    17482 => 63,
    17483 => 63,
    17484 => 63,
    17485 => 63,
    17486 => 63,
    17487 => 63,
    17488 => 63,
    17489 => 63,
    17490 => 63,
    17491 => 63,
    17492 => 63,
    17493 => 63,
    17494 => 63,
    17495 => 63,
    17496 => 63,
    17497 => 63,
    17498 => 63,
    17499 => 63,
    17500 => 63,
    17501 => 63,
    17502 => 63,
    17503 => 63,
    17504 => 63,
    17505 => 63,
    17506 => 63,
    17507 => 63,
    17508 => 63,
    17509 => 63,
    17510 => 63,
    17511 => 63,
    17512 => 63,
    17513 => 63,
    17514 => 63,
    17515 => 63,
    17516 => 63,
    17517 => 63,
    17518 => 63,
    17519 => 63,
    17520 => 63,
    17521 => 63,
    17522 => 63,
    17523 => 63,
    17524 => 63,
    17525 => 63,
    17526 => 63,
    17527 => 63,
    17528 => 63,
    17529 => 63,
    17530 => 63,
    17531 => 63,
    17532 => 63,
    17533 => 63,
    17534 => 63,
    17535 => 63,
    17536 => 63,
    17537 => 63,
    17538 => 63,
    17539 => 63,
    17540 => 63,
    17541 => 63,
    17542 => 63,
    17543 => 63,
    17544 => 63,
    17545 => 63,
    17546 => 63,
    17547 => 63,
    17548 => 63,
    17549 => 63,
    17550 => 63,
    17551 => 63,
    17552 => 63,
    17553 => 63,
    17554 => 63,
    17555 => 63,
    17556 => 63,
    17557 => 63,
    17558 => 63,
    17559 => 63,
    17560 => 63,
    17561 => 63,
    17562 => 63,
    17563 => 63,
    17564 => 63,
    17565 => 63,
    17566 => 63,
    17567 => 63,
    17568 => 63,
    17569 => 63,
    17570 => 63,
    17571 => 63,
    17572 => 63,
    17573 => 63,
    17574 => 63,
    17575 => 63,
    17576 => 63,
    17577 => 63,
    17578 => 63,
    17579 => 63,
    17580 => 63,
    17581 => 63,
    17582 => 63,
    17583 => 63,
    17584 => 63,
    17585 => 63,
    17586 => 63,
    17587 => 63,
    17588 => 63,
    17589 => 63,
    17590 => 63,
    17591 => 63,
    17592 => 63,
    17593 => 63,
    17594 => 63,
    17595 => 63,
    17596 => 63,
    17597 => 63,
    17598 => 63,
    17599 => 63,
    17600 => 63,
    17601 => 63,
    17602 => 63,
    17603 => 63,
    17604 => 63,
    17605 => 63,
    17606 => 63,
    17607 => 63,
    17608 => 63,
    17609 => 63,
    17610 => 63,
    17611 => 63,
    17612 => 63,
    17613 => 63,
    17614 => 63,
    17615 => 63,
    17616 => 63,
    17617 => 63,
    17618 => 63,
    17619 => 63,
    17620 => 63,
    17621 => 63,
    17622 => 63,
    17623 => 63,
    17624 => 63,
    17625 => 63,
    17626 => 63,
    17627 => 63,
    17628 => 63,
    17629 => 63,
    17630 => 63,
    17631 => 63,
    17632 => 63,
    17633 => 63,
    17634 => 63,
    17635 => 63,
    17636 => 63,
    17637 => 63,
    17638 => 63,
    17639 => 63,
    17640 => 63,
    17641 => 63,
    17642 => 63,
    17643 => 63,
    17644 => 63,
    17645 => 63,
    17646 => 63,
    17647 => 63,
    17648 => 63,
    17649 => 63,
    17650 => 63,
    17651 => 63,
    17652 => 63,
    17653 => 63,
    17654 => 63,
    17655 => 63,
    17656 => 63,
    17657 => 63,
    17658 => 63,
    17659 => 63,
    17660 => 63,
    17661 => 63,
    17662 => 63,
    17663 => 63,
    17664 => 63,
    17665 => 63,
    17666 => 63,
    17667 => 63,
    17668 => 63,
    17669 => 63,
    17670 => 63,
    17671 => 63,
    17672 => 63,
    17673 => 63,
    17674 => 63,
    17675 => 63,
    17676 => 63,
    17677 => 63,
    17678 => 63,
    17679 => 63,
    17680 => 63,
    17681 => 63,
    17682 => 63,
    17683 => 63,
    17684 => 63,
    17685 => 63,
    17686 => 63,
    17687 => 63,
    17688 => 63,
    17689 => 63,
    17690 => 63,
    17691 => 63,
    17692 => 63,
    17693 => 63,
    17694 => 63,
    17695 => 63,
    17696 => 63,
    17697 => 63,
    17698 => 63,
    17699 => 62,
    17700 => 62,
    17701 => 62,
    17702 => 62,
    17703 => 62,
    17704 => 62,
    17705 => 62,
    17706 => 62,
    17707 => 62,
    17708 => 62,
    17709 => 62,
    17710 => 62,
    17711 => 62,
    17712 => 62,
    17713 => 62,
    17714 => 62,
    17715 => 62,
    17716 => 62,
    17717 => 62,
    17718 => 62,
    17719 => 62,
    17720 => 62,
    17721 => 62,
    17722 => 62,
    17723 => 62,
    17724 => 62,
    17725 => 62,
    17726 => 62,
    17727 => 62,
    17728 => 62,
    17729 => 62,
    17730 => 62,
    17731 => 62,
    17732 => 62,
    17733 => 62,
    17734 => 62,
    17735 => 62,
    17736 => 62,
    17737 => 62,
    17738 => 62,
    17739 => 62,
    17740 => 62,
    17741 => 62,
    17742 => 62,
    17743 => 62,
    17744 => 62,
    17745 => 62,
    17746 => 62,
    17747 => 62,
    17748 => 62,
    17749 => 62,
    17750 => 62,
    17751 => 62,
    17752 => 62,
    17753 => 62,
    17754 => 62,
    17755 => 62,
    17756 => 62,
    17757 => 62,
    17758 => 62,
    17759 => 62,
    17760 => 62,
    17761 => 62,
    17762 => 62,
    17763 => 62,
    17764 => 62,
    17765 => 62,
    17766 => 62,
    17767 => 62,
    17768 => 62,
    17769 => 62,
    17770 => 62,
    17771 => 62,
    17772 => 62,
    17773 => 62,
    17774 => 62,
    17775 => 62,
    17776 => 62,
    17777 => 62,
    17778 => 62,
    17779 => 62,
    17780 => 62,
    17781 => 62,
    17782 => 62,
    17783 => 62,
    17784 => 62,
    17785 => 62,
    17786 => 62,
    17787 => 62,
    17788 => 62,
    17789 => 62,
    17790 => 62,
    17791 => 62,
    17792 => 62,
    17793 => 62,
    17794 => 62,
    17795 => 62,
    17796 => 62,
    17797 => 62,
    17798 => 62,
    17799 => 62,
    17800 => 62,
    17801 => 62,
    17802 => 62,
    17803 => 62,
    17804 => 62,
    17805 => 62,
    17806 => 62,
    17807 => 62,
    17808 => 62,
    17809 => 62,
    17810 => 62,
    17811 => 62,
    17812 => 62,
    17813 => 62,
    17814 => 62,
    17815 => 62,
    17816 => 62,
    17817 => 62,
    17818 => 62,
    17819 => 62,
    17820 => 62,
    17821 => 62,
    17822 => 62,
    17823 => 62,
    17824 => 62,
    17825 => 62,
    17826 => 62,
    17827 => 62,
    17828 => 62,
    17829 => 62,
    17830 => 62,
    17831 => 62,
    17832 => 62,
    17833 => 62,
    17834 => 62,
    17835 => 62,
    17836 => 62,
    17837 => 62,
    17838 => 62,
    17839 => 62,
    17840 => 62,
    17841 => 62,
    17842 => 62,
    17843 => 62,
    17844 => 62,
    17845 => 62,
    17846 => 62,
    17847 => 62,
    17848 => 62,
    17849 => 62,
    17850 => 62,
    17851 => 62,
    17852 => 62,
    17853 => 62,
    17854 => 62,
    17855 => 62,
    17856 => 62,
    17857 => 62,
    17858 => 62,
    17859 => 62,
    17860 => 62,
    17861 => 62,
    17862 => 62,
    17863 => 62,
    17864 => 62,
    17865 => 62,
    17866 => 62,
    17867 => 62,
    17868 => 62,
    17869 => 62,
    17870 => 62,
    17871 => 62,
    17872 => 62,
    17873 => 62,
    17874 => 62,
    17875 => 62,
    17876 => 62,
    17877 => 62,
    17878 => 62,
    17879 => 62,
    17880 => 62,
    17881 => 62,
    17882 => 62,
    17883 => 62,
    17884 => 62,
    17885 => 62,
    17886 => 62,
    17887 => 62,
    17888 => 62,
    17889 => 62,
    17890 => 62,
    17891 => 62,
    17892 => 62,
    17893 => 62,
    17894 => 62,
    17895 => 62,
    17896 => 62,
    17897 => 62,
    17898 => 62,
    17899 => 62,
    17900 => 62,
    17901 => 62,
    17902 => 62,
    17903 => 62,
    17904 => 62,
    17905 => 62,
    17906 => 62,
    17907 => 62,
    17908 => 62,
    17909 => 62,
    17910 => 62,
    17911 => 62,
    17912 => 62,
    17913 => 62,
    17914 => 62,
    17915 => 62,
    17916 => 62,
    17917 => 62,
    17918 => 62,
    17919 => 62,
    17920 => 62,
    17921 => 62,
    17922 => 62,
    17923 => 62,
    17924 => 62,
    17925 => 62,
    17926 => 62,
    17927 => 62,
    17928 => 62,
    17929 => 62,
    17930 => 62,
    17931 => 62,
    17932 => 62,
    17933 => 62,
    17934 => 62,
    17935 => 62,
    17936 => 62,
    17937 => 62,
    17938 => 62,
    17939 => 62,
    17940 => 62,
    17941 => 62,
    17942 => 62,
    17943 => 62,
    17944 => 62,
    17945 => 62,
    17946 => 62,
    17947 => 62,
    17948 => 62,
    17949 => 62,
    17950 => 62,
    17951 => 62,
    17952 => 62,
    17953 => 62,
    17954 => 62,
    17955 => 62,
    17956 => 62,
    17957 => 62,
    17958 => 62,
    17959 => 62,
    17960 => 62,
    17961 => 62,
    17962 => 62,
    17963 => 62,
    17964 => 62,
    17965 => 62,
    17966 => 62,
    17967 => 62,
    17968 => 62,
    17969 => 62,
    17970 => 62,
    17971 => 62,
    17972 => 62,
    17973 => 62,
    17974 => 62,
    17975 => 62,
    17976 => 62,
    17977 => 62,
    17978 => 62,
    17979 => 62,
    17980 => 62,
    17981 => 62,
    17982 => 62,
    17983 => 62,
    17984 => 62,
    17985 => 62,
    17986 => 62,
    17987 => 62,
    17988 => 62,
    17989 => 62,
    17990 => 62,
    17991 => 62,
    17992 => 62,
    17993 => 62,
    17994 => 62,
    17995 => 62,
    17996 => 62,
    17997 => 62,
    17998 => 62,
    17999 => 62,
    18000 => 62,
    18001 => 62,
    18002 => 62,
    18003 => 62,
    18004 => 62,
    18005 => 62,
    18006 => 62,
    18007 => 62,
    18008 => 62,
    18009 => 62,
    18010 => 62,
    18011 => 62,
    18012 => 62,
    18013 => 62,
    18014 => 62,
    18015 => 62,
    18016 => 62,
    18017 => 62,
    18018 => 62,
    18019 => 62,
    18020 => 62,
    18021 => 62,
    18022 => 62,
    18023 => 62,
    18024 => 62,
    18025 => 62,
    18026 => 62,
    18027 => 62,
    18028 => 62,
    18029 => 62,
    18030 => 62,
    18031 => 62,
    18032 => 62,
    18033 => 62,
    18034 => 62,
    18035 => 62,
    18036 => 62,
    18037 => 62,
    18038 => 62,
    18039 => 62,
    18040 => 62,
    18041 => 62,
    18042 => 62,
    18043 => 62,
    18044 => 62,
    18045 => 62,
    18046 => 62,
    18047 => 62,
    18048 => 62,
    18049 => 62,
    18050 => 62,
    18051 => 62,
    18052 => 62,
    18053 => 62,
    18054 => 62,
    18055 => 62,
    18056 => 62,
    18057 => 62,
    18058 => 62,
    18059 => 62,
    18060 => 62,
    18061 => 62,
    18062 => 62,
    18063 => 62,
    18064 => 62,
    18065 => 62,
    18066 => 62,
    18067 => 62,
    18068 => 62,
    18069 => 62,
    18070 => 62,
    18071 => 62,
    18072 => 62,
    18073 => 62,
    18074 => 62,
    18075 => 62,
    18076 => 62,
    18077 => 62,
    18078 => 62,
    18079 => 62,
    18080 => 62,
    18081 => 62,
    18082 => 62,
    18083 => 62,
    18084 => 62,
    18085 => 62,
    18086 => 62,
    18087 => 62,
    18088 => 62,
    18089 => 62,
    18090 => 62,
    18091 => 62,
    18092 => 62,
    18093 => 62,
    18094 => 62,
    18095 => 62,
    18096 => 62,
    18097 => 62,
    18098 => 62,
    18099 => 62,
    18100 => 62,
    18101 => 62,
    18102 => 62,
    18103 => 62,
    18104 => 62,
    18105 => 62,
    18106 => 62,
    18107 => 62,
    18108 => 62,
    18109 => 62,
    18110 => 62,
    18111 => 62,
    18112 => 62,
    18113 => 62,
    18114 => 62,
    18115 => 62,
    18116 => 62,
    18117 => 62,
    18118 => 62,
    18119 => 62,
    18120 => 62,
    18121 => 62,
    18122 => 62,
    18123 => 62,
    18124 => 62,
    18125 => 62,
    18126 => 62,
    18127 => 62,
    18128 => 62,
    18129 => 62,
    18130 => 62,
    18131 => 62,
    18132 => 62,
    18133 => 62,
    18134 => 62,
    18135 => 62,
    18136 => 62,
    18137 => 62,
    18138 => 62,
    18139 => 62,
    18140 => 62,
    18141 => 62,
    18142 => 62,
    18143 => 62,
    18144 => 62,
    18145 => 62,
    18146 => 62,
    18147 => 62,
    18148 => 62,
    18149 => 62,
    18150 => 62,
    18151 => 62,
    18152 => 62,
    18153 => 62,
    18154 => 62,
    18155 => 62,
    18156 => 62,
    18157 => 62,
    18158 => 62,
    18159 => 62,
    18160 => 62,
    18161 => 62,
    18162 => 62,
    18163 => 62,
    18164 => 62,
    18165 => 62,
    18166 => 62,
    18167 => 62,
    18168 => 62,
    18169 => 62,
    18170 => 62,
    18171 => 62,
    18172 => 62,
    18173 => 62,
    18174 => 62,
    18175 => 62,
    18176 => 62,
    18177 => 62,
    18178 => 62,
    18179 => 62,
    18180 => 62,
    18181 => 62,
    18182 => 62,
    18183 => 62,
    18184 => 62,
    18185 => 62,
    18186 => 62,
    18187 => 62,
    18188 => 62,
    18189 => 62,
    18190 => 62,
    18191 => 62,
    18192 => 62,
    18193 => 62,
    18194 => 62,
    18195 => 62,
    18196 => 62,
    18197 => 62,
    18198 => 62,
    18199 => 62,
    18200 => 62,
    18201 => 62,
    18202 => 62,
    18203 => 62,
    18204 => 62,
    18205 => 62,
    18206 => 62,
    18207 => 62,
    18208 => 62,
    18209 => 62,
    18210 => 62,
    18211 => 62,
    18212 => 62,
    18213 => 62,
    18214 => 62,
    18215 => 62,
    18216 => 62,
    18217 => 62,
    18218 => 62,
    18219 => 62,
    18220 => 62,
    18221 => 62,
    18222 => 62,
    18223 => 62,
    18224 => 62,
    18225 => 62,
    18226 => 62,
    18227 => 62,
    18228 => 62,
    18229 => 62,
    18230 => 62,
    18231 => 62,
    18232 => 62,
    18233 => 62,
    18234 => 62,
    18235 => 62,
    18236 => 62,
    18237 => 62,
    18238 => 62,
    18239 => 62,
    18240 => 62,
    18241 => 62,
    18242 => 62,
    18243 => 62,
    18244 => 62,
    18245 => 62,
    18246 => 62,
    18247 => 62,
    18248 => 62,
    18249 => 62,
    18250 => 62,
    18251 => 62,
    18252 => 62,
    18253 => 62,
    18254 => 62,
    18255 => 62,
    18256 => 62,
    18257 => 62,
    18258 => 62,
    18259 => 62,
    18260 => 62,
    18261 => 62,
    18262 => 62,
    18263 => 62,
    18264 => 62,
    18265 => 62,
    18266 => 62,
    18267 => 62,
    18268 => 62,
    18269 => 62,
    18270 => 62,
    18271 => 62,
    18272 => 62,
    18273 => 62,
    18274 => 62,
    18275 => 62,
    18276 => 62,
    18277 => 62,
    18278 => 62,
    18279 => 62,
    18280 => 62,
    18281 => 62,
    18282 => 62,
    18283 => 62,
    18284 => 62,
    18285 => 62,
    18286 => 62,
    18287 => 62,
    18288 => 62,
    18289 => 62,
    18290 => 62,
    18291 => 62,
    18292 => 62,
    18293 => 62,
    18294 => 62,
    18295 => 62,
    18296 => 62,
    18297 => 62,
    18298 => 62,
    18299 => 62,
    18300 => 62,
    18301 => 62,
    18302 => 62,
    18303 => 62,
    18304 => 62,
    18305 => 62,
    18306 => 62,
    18307 => 62,
    18308 => 62,
    18309 => 62,
    18310 => 62,
    18311 => 62,
    18312 => 62,
    18313 => 62,
    18314 => 62,
    18315 => 62,
    18316 => 62,
    18317 => 62,
    18318 => 62,
    18319 => 62,
    18320 => 62,
    18321 => 62,
    18322 => 62,
    18323 => 62,
    18324 => 62,
    18325 => 62,
    18326 => 62,
    18327 => 62,
    18328 => 62,
    18329 => 62,
    18330 => 62,
    18331 => 62,
    18332 => 62,
    18333 => 62,
    18334 => 62,
    18335 => 62,
    18336 => 62,
    18337 => 62,
    18338 => 62,
    18339 => 62,
    18340 => 62,
    18341 => 62,
    18342 => 62,
    18343 => 62,
    18344 => 62,
    18345 => 62,
    18346 => 62,
    18347 => 62,
    18348 => 62,
    18349 => 62,
    18350 => 62,
    18351 => 62,
    18352 => 62,
    18353 => 62,
    18354 => 62,
    18355 => 62,
    18356 => 62,
    18357 => 62,
    18358 => 62,
    18359 => 62,
    18360 => 62,
    18361 => 62,
    18362 => 62,
    18363 => 62,
    18364 => 62,
    18365 => 62,
    18366 => 62,
    18367 => 62,
    18368 => 62,
    18369 => 62,
    18370 => 62,
    18371 => 62,
    18372 => 62,
    18373 => 62,
    18374 => 62,
    18375 => 62,
    18376 => 62,
    18377 => 62,
    18378 => 62,
    18379 => 62,
    18380 => 62,
    18381 => 62,
    18382 => 62,
    18383 => 62,
    18384 => 62,
    18385 => 62,
    18386 => 62,
    18387 => 62,
    18388 => 62,
    18389 => 62,
    18390 => 62,
    18391 => 62,
    18392 => 62,
    18393 => 62,
    18394 => 62,
    18395 => 62,
    18396 => 62,
    18397 => 62,
    18398 => 62,
    18399 => 62,
    18400 => 62,
    18401 => 62,
    18402 => 62,
    18403 => 62,
    18404 => 62,
    18405 => 62,
    18406 => 62,
    18407 => 62,
    18408 => 62,
    18409 => 62,
    18410 => 62,
    18411 => 62,
    18412 => 62,
    18413 => 62,
    18414 => 62,
    18415 => 62,
    18416 => 62,
    18417 => 62,
    18418 => 62,
    18419 => 62,
    18420 => 62,
    18421 => 62,
    18422 => 62,
    18423 => 62,
    18424 => 62,
    18425 => 62,
    18426 => 62,
    18427 => 62,
    18428 => 62,
    18429 => 62,
    18430 => 62,
    18431 => 62,
    18432 => 62,
    18433 => 62,
    18434 => 62,
    18435 => 62,
    18436 => 62,
    18437 => 62,
    18438 => 62,
    18439 => 62,
    18440 => 62,
    18441 => 62,
    18442 => 62,
    18443 => 62,
    18444 => 62,
    18445 => 62,
    18446 => 62,
    18447 => 62,
    18448 => 62,
    18449 => 62,
    18450 => 62,
    18451 => 62,
    18452 => 62,
    18453 => 62,
    18454 => 62,
    18455 => 62,
    18456 => 62,
    18457 => 62,
    18458 => 62,
    18459 => 62,
    18460 => 62,
    18461 => 62,
    18462 => 62,
    18463 => 62,
    18464 => 62,
    18465 => 62,
    18466 => 62,
    18467 => 62,
    18468 => 62,
    18469 => 62,
    18470 => 62,
    18471 => 62,
    18472 => 62,
    18473 => 62,
    18474 => 62,
    18475 => 62,
    18476 => 62,
    18477 => 62,
    18478 => 62,
    18479 => 62,
    18480 => 62,
    18481 => 62,
    18482 => 62,
    18483 => 62,
    18484 => 62,
    18485 => 62,
    18486 => 62,
    18487 => 62,
    18488 => 62,
    18489 => 62,
    18490 => 62,
    18491 => 62,
    18492 => 62,
    18493 => 62,
    18494 => 62,
    18495 => 62,
    18496 => 62,
    18497 => 62,
    18498 => 62,
    18499 => 62,
    18500 => 62,
    18501 => 62,
    18502 => 62,
    18503 => 62,
    18504 => 62,
    18505 => 62,
    18506 => 62,
    18507 => 62,
    18508 => 62,
    18509 => 62,
    18510 => 62,
    18511 => 62,
    18512 => 62,
    18513 => 62,
    18514 => 62,
    18515 => 62,
    18516 => 62,
    18517 => 62,
    18518 => 62,
    18519 => 62,
    18520 => 62,
    18521 => 62,
    18522 => 62,
    18523 => 62,
    18524 => 62,
    18525 => 62,
    18526 => 62,
    18527 => 62,
    18528 => 62,
    18529 => 62,
    18530 => 62,
    18531 => 62,
    18532 => 62,
    18533 => 62,
    18534 => 62,
    18535 => 62,
    18536 => 62,
    18537 => 62,
    18538 => 62,
    18539 => 62,
    18540 => 62,
    18541 => 62,
    18542 => 62,
    18543 => 62,
    18544 => 62,
    18545 => 62,
    18546 => 62,
    18547 => 62,
    18548 => 62,
    18549 => 62,
    18550 => 62,
    18551 => 62,
    18552 => 62,
    18553 => 62,
    18554 => 62,
    18555 => 62,
    18556 => 62,
    18557 => 62,
    18558 => 62,
    18559 => 62,
    18560 => 62,
    18561 => 62,
    18562 => 62,
    18563 => 62,
    18564 => 62,
    18565 => 62,
    18566 => 62,
    18567 => 62,
    18568 => 62,
    18569 => 62,
    18570 => 62,
    18571 => 62,
    18572 => 62,
    18573 => 62,
    18574 => 62,
    18575 => 62,
    18576 => 62,
    18577 => 62,
    18578 => 62,
    18579 => 62,
    18580 => 62,
    18581 => 62,
    18582 => 62,
    18583 => 62,
    18584 => 62,
    18585 => 62,
    18586 => 62,
    18587 => 62,
    18588 => 62,
    18589 => 62,
    18590 => 62,
    18591 => 62,
    18592 => 62,
    18593 => 62,
    18594 => 62,
    18595 => 62,
    18596 => 62,
    18597 => 62,
    18598 => 62,
    18599 => 62,
    18600 => 62,
    18601 => 62,
    18602 => 62,
    18603 => 62,
    18604 => 62,
    18605 => 62,
    18606 => 62,
    18607 => 62,
    18608 => 62,
    18609 => 62,
    18610 => 62,
    18611 => 62,
    18612 => 62,
    18613 => 62,
    18614 => 62,
    18615 => 62,
    18616 => 62,
    18617 => 62,
    18618 => 62,
    18619 => 62,
    18620 => 62,
    18621 => 62,
    18622 => 62,
    18623 => 62,
    18624 => 62,
    18625 => 62,
    18626 => 62,
    18627 => 62,
    18628 => 62,
    18629 => 62,
    18630 => 62,
    18631 => 62,
    18632 => 62,
    18633 => 62,
    18634 => 62,
    18635 => 62,
    18636 => 62,
    18637 => 62,
    18638 => 62,
    18639 => 62,
    18640 => 62,
    18641 => 62,
    18642 => 62,
    18643 => 62,
    18644 => 62,
    18645 => 62,
    18646 => 62,
    18647 => 62,
    18648 => 62,
    18649 => 62,
    18650 => 62,
    18651 => 62,
    18652 => 62,
    18653 => 62,
    18654 => 62,
    18655 => 62,
    18656 => 62,
    18657 => 62,
    18658 => 62,
    18659 => 62,
    18660 => 62,
    18661 => 62,
    18662 => 62,
    18663 => 62,
    18664 => 62,
    18665 => 61,
    18666 => 61,
    18667 => 61,
    18668 => 61,
    18669 => 61,
    18670 => 61,
    18671 => 61,
    18672 => 61,
    18673 => 61,
    18674 => 61,
    18675 => 61,
    18676 => 61,
    18677 => 61,
    18678 => 61,
    18679 => 61,
    18680 => 61,
    18681 => 61,
    18682 => 61,
    18683 => 61,
    18684 => 61,
    18685 => 61,
    18686 => 61,
    18687 => 61,
    18688 => 61,
    18689 => 61,
    18690 => 61,
    18691 => 61,
    18692 => 61,
    18693 => 61,
    18694 => 61,
    18695 => 61,
    18696 => 61,
    18697 => 61,
    18698 => 61,
    18699 => 61,
    18700 => 61,
    18701 => 61,
    18702 => 61,
    18703 => 61,
    18704 => 61,
    18705 => 61,
    18706 => 61,
    18707 => 61,
    18708 => 61,
    18709 => 61,
    18710 => 61,
    18711 => 61,
    18712 => 61,
    18713 => 61,
    18714 => 61,
    18715 => 61,
    18716 => 61,
    18717 => 61,
    18718 => 61,
    18719 => 61,
    18720 => 61,
    18721 => 61,
    18722 => 61,
    18723 => 61,
    18724 => 61,
    18725 => 61,
    18726 => 61,
    18727 => 61,
    18728 => 61,
    18729 => 61,
    18730 => 61,
    18731 => 61,
    18732 => 61,
    18733 => 61,
    18734 => 61,
    18735 => 61,
    18736 => 61,
    18737 => 61,
    18738 => 61,
    18739 => 61,
    18740 => 61,
    18741 => 61,
    18742 => 61,
    18743 => 61,
    18744 => 61,
    18745 => 61,
    18746 => 61,
    18747 => 61,
    18748 => 61,
    18749 => 61,
    18750 => 61,
    18751 => 61,
    18752 => 61,
    18753 => 61,
    18754 => 61,
    18755 => 61,
    18756 => 61,
    18757 => 61,
    18758 => 61,
    18759 => 61,
    18760 => 61,
    18761 => 61,
    18762 => 61,
    18763 => 61,
    18764 => 61,
    18765 => 61,
    18766 => 61,
    18767 => 61,
    18768 => 61,
    18769 => 61,
    18770 => 61,
    18771 => 61,
    18772 => 61,
    18773 => 61,
    18774 => 61,
    18775 => 61,
    18776 => 61,
    18777 => 61,
    18778 => 61,
    18779 => 61,
    18780 => 61,
    18781 => 61,
    18782 => 61,
    18783 => 61,
    18784 => 61,
    18785 => 61,
    18786 => 61,
    18787 => 61,
    18788 => 61,
    18789 => 61,
    18790 => 61,
    18791 => 61,
    18792 => 61,
    18793 => 61,
    18794 => 61,
    18795 => 61,
    18796 => 61,
    18797 => 61,
    18798 => 61,
    18799 => 61,
    18800 => 61,
    18801 => 61,
    18802 => 61,
    18803 => 61,
    18804 => 61,
    18805 => 61,
    18806 => 61,
    18807 => 61,
    18808 => 61,
    18809 => 61,
    18810 => 61,
    18811 => 61,
    18812 => 61,
    18813 => 61,
    18814 => 61,
    18815 => 61,
    18816 => 61,
    18817 => 61,
    18818 => 61,
    18819 => 61,
    18820 => 61,
    18821 => 61,
    18822 => 61,
    18823 => 61,
    18824 => 61,
    18825 => 61,
    18826 => 61,
    18827 => 61,
    18828 => 61,
    18829 => 61,
    18830 => 61,
    18831 => 61,
    18832 => 61,
    18833 => 61,
    18834 => 61,
    18835 => 61,
    18836 => 61,
    18837 => 61,
    18838 => 61,
    18839 => 61,
    18840 => 61,
    18841 => 61,
    18842 => 61,
    18843 => 61,
    18844 => 61,
    18845 => 61,
    18846 => 61,
    18847 => 61,
    18848 => 61,
    18849 => 61,
    18850 => 61,
    18851 => 61,
    18852 => 61,
    18853 => 61,
    18854 => 61,
    18855 => 61,
    18856 => 61,
    18857 => 61,
    18858 => 61,
    18859 => 61,
    18860 => 61,
    18861 => 61,
    18862 => 61,
    18863 => 61,
    18864 => 61,
    18865 => 61,
    18866 => 61,
    18867 => 61,
    18868 => 61,
    18869 => 61,
    18870 => 61,
    18871 => 61,
    18872 => 61,
    18873 => 61,
    18874 => 61,
    18875 => 61,
    18876 => 61,
    18877 => 61,
    18878 => 61,
    18879 => 61,
    18880 => 61,
    18881 => 61,
    18882 => 61,
    18883 => 61,
    18884 => 61,
    18885 => 61,
    18886 => 61,
    18887 => 61,
    18888 => 61,
    18889 => 61,
    18890 => 61,
    18891 => 61,
    18892 => 61,
    18893 => 61,
    18894 => 61,
    18895 => 61,
    18896 => 61,
    18897 => 61,
    18898 => 61,
    18899 => 61,
    18900 => 61,
    18901 => 61,
    18902 => 61,
    18903 => 61,
    18904 => 61,
    18905 => 61,
    18906 => 61,
    18907 => 61,
    18908 => 61,
    18909 => 61,
    18910 => 61,
    18911 => 61,
    18912 => 61,
    18913 => 61,
    18914 => 61,
    18915 => 61,
    18916 => 61,
    18917 => 61,
    18918 => 61,
    18919 => 61,
    18920 => 61,
    18921 => 61,
    18922 => 61,
    18923 => 61,
    18924 => 61,
    18925 => 61,
    18926 => 61,
    18927 => 61,
    18928 => 61,
    18929 => 61,
    18930 => 61,
    18931 => 61,
    18932 => 61,
    18933 => 61,
    18934 => 61,
    18935 => 61,
    18936 => 61,
    18937 => 61,
    18938 => 61,
    18939 => 61,
    18940 => 61,
    18941 => 61,
    18942 => 61,
    18943 => 61,
    18944 => 61,
    18945 => 61,
    18946 => 61,
    18947 => 61,
    18948 => 61,
    18949 => 61,
    18950 => 61,
    18951 => 61,
    18952 => 61,
    18953 => 61,
    18954 => 61,
    18955 => 61,
    18956 => 61,
    18957 => 61,
    18958 => 61,
    18959 => 61,
    18960 => 61,
    18961 => 61,
    18962 => 61,
    18963 => 61,
    18964 => 61,
    18965 => 61,
    18966 => 61,
    18967 => 61,
    18968 => 61,
    18969 => 61,
    18970 => 61,
    18971 => 61,
    18972 => 61,
    18973 => 61,
    18974 => 61,
    18975 => 61,
    18976 => 61,
    18977 => 61,
    18978 => 61,
    18979 => 61,
    18980 => 61,
    18981 => 61,
    18982 => 61,
    18983 => 61,
    18984 => 61,
    18985 => 61,
    18986 => 61,
    18987 => 61,
    18988 => 61,
    18989 => 61,
    18990 => 61,
    18991 => 61,
    18992 => 61,
    18993 => 61,
    18994 => 61,
    18995 => 61,
    18996 => 61,
    18997 => 61,
    18998 => 61,
    18999 => 61,
    19000 => 61,
    19001 => 61,
    19002 => 61,
    19003 => 61,
    19004 => 61,
    19005 => 61,
    19006 => 61,
    19007 => 61,
    19008 => 61,
    19009 => 61,
    19010 => 61,
    19011 => 61,
    19012 => 61,
    19013 => 61,
    19014 => 61,
    19015 => 61,
    19016 => 61,
    19017 => 61,
    19018 => 61,
    19019 => 61,
    19020 => 61,
    19021 => 61,
    19022 => 61,
    19023 => 61,
    19024 => 61,
    19025 => 61,
    19026 => 61,
    19027 => 61,
    19028 => 61,
    19029 => 61,
    19030 => 61,
    19031 => 61,
    19032 => 61,
    19033 => 61,
    19034 => 61,
    19035 => 61,
    19036 => 61,
    19037 => 61,
    19038 => 61,
    19039 => 61,
    19040 => 61,
    19041 => 61,
    19042 => 61,
    19043 => 61,
    19044 => 61,
    19045 => 61,
    19046 => 61,
    19047 => 61,
    19048 => 61,
    19049 => 61,
    19050 => 61,
    19051 => 61,
    19052 => 61,
    19053 => 61,
    19054 => 61,
    19055 => 61,
    19056 => 61,
    19057 => 61,
    19058 => 61,
    19059 => 61,
    19060 => 61,
    19061 => 61,
    19062 => 61,
    19063 => 61,
    19064 => 61,
    19065 => 61,
    19066 => 61,
    19067 => 61,
    19068 => 61,
    19069 => 61,
    19070 => 61,
    19071 => 61,
    19072 => 61,
    19073 => 61,
    19074 => 61,
    19075 => 61,
    19076 => 61,
    19077 => 61,
    19078 => 61,
    19079 => 61,
    19080 => 61,
    19081 => 61,
    19082 => 61,
    19083 => 61,
    19084 => 61,
    19085 => 61,
    19086 => 61,
    19087 => 61,
    19088 => 61,
    19089 => 61,
    19090 => 61,
    19091 => 61,
    19092 => 61,
    19093 => 61,
    19094 => 61,
    19095 => 61,
    19096 => 61,
    19097 => 61,
    19098 => 61,
    19099 => 61,
    19100 => 61,
    19101 => 61,
    19102 => 61,
    19103 => 61,
    19104 => 61,
    19105 => 61,
    19106 => 61,
    19107 => 61,
    19108 => 61,
    19109 => 61,
    19110 => 61,
    19111 => 61,
    19112 => 61,
    19113 => 61,
    19114 => 61,
    19115 => 61,
    19116 => 61,
    19117 => 61,
    19118 => 61,
    19119 => 61,
    19120 => 61,
    19121 => 61,
    19122 => 61,
    19123 => 61,
    19124 => 61,
    19125 => 61,
    19126 => 61,
    19127 => 61,
    19128 => 61,
    19129 => 61,
    19130 => 61,
    19131 => 61,
    19132 => 61,
    19133 => 61,
    19134 => 61,
    19135 => 61,
    19136 => 61,
    19137 => 61,
    19138 => 61,
    19139 => 61,
    19140 => 61,
    19141 => 61,
    19142 => 61,
    19143 => 61,
    19144 => 61,
    19145 => 61,
    19146 => 61,
    19147 => 61,
    19148 => 61,
    19149 => 61,
    19150 => 61,
    19151 => 61,
    19152 => 61,
    19153 => 61,
    19154 => 61,
    19155 => 61,
    19156 => 61,
    19157 => 61,
    19158 => 61,
    19159 => 61,
    19160 => 61,
    19161 => 61,
    19162 => 61,
    19163 => 61,
    19164 => 61,
    19165 => 61,
    19166 => 61,
    19167 => 61,
    19168 => 61,
    19169 => 61,
    19170 => 61,
    19171 => 61,
    19172 => 61,
    19173 => 61,
    19174 => 61,
    19175 => 61,
    19176 => 61,
    19177 => 61,
    19178 => 61,
    19179 => 61,
    19180 => 61,
    19181 => 61,
    19182 => 61,
    19183 => 61,
    19184 => 61,
    19185 => 61,
    19186 => 61,
    19187 => 61,
    19188 => 61,
    19189 => 61,
    19190 => 61,
    19191 => 61,
    19192 => 61,
    19193 => 61,
    19194 => 61,
    19195 => 61,
    19196 => 61,
    19197 => 61,
    19198 => 61,
    19199 => 61,
    19200 => 61,
    19201 => 61,
    19202 => 61,
    19203 => 61,
    19204 => 61,
    19205 => 61,
    19206 => 61,
    19207 => 61,
    19208 => 61,
    19209 => 61,
    19210 => 61,
    19211 => 61,
    19212 => 61,
    19213 => 61,
    19214 => 61,
    19215 => 61,
    19216 => 61,
    19217 => 61,
    19218 => 61,
    19219 => 61,
    19220 => 61,
    19221 => 61,
    19222 => 61,
    19223 => 61,
    19224 => 61,
    19225 => 61,
    19226 => 61,
    19227 => 61,
    19228 => 61,
    19229 => 61,
    19230 => 61,
    19231 => 61,
    19232 => 61,
    19233 => 61,
    19234 => 61,
    19235 => 61,
    19236 => 61,
    19237 => 61,
    19238 => 61,
    19239 => 61,
    19240 => 61,
    19241 => 61,
    19242 => 61,
    19243 => 61,
    19244 => 61,
    19245 => 61,
    19246 => 61,
    19247 => 61,
    19248 => 61,
    19249 => 61,
    19250 => 61,
    19251 => 61,
    19252 => 61,
    19253 => 61,
    19254 => 61,
    19255 => 61,
    19256 => 61,
    19257 => 61,
    19258 => 61,
    19259 => 61,
    19260 => 61,
    19261 => 61,
    19262 => 61,
    19263 => 61,
    19264 => 61,
    19265 => 61,
    19266 => 61,
    19267 => 61,
    19268 => 61,
    19269 => 61,
    19270 => 61,
    19271 => 61,
    19272 => 61,
    19273 => 61,
    19274 => 61,
    19275 => 61,
    19276 => 61,
    19277 => 61,
    19278 => 61,
    19279 => 61,
    19280 => 61,
    19281 => 61,
    19282 => 61,
    19283 => 61,
    19284 => 61,
    19285 => 61,
    19286 => 61,
    19287 => 61,
    19288 => 61,
    19289 => 61,
    19290 => 61,
    19291 => 61,
    19292 => 61,
    19293 => 61,
    19294 => 61,
    19295 => 61,
    19296 => 61,
    19297 => 61,
    19298 => 61,
    19299 => 61,
    19300 => 61,
    19301 => 61,
    19302 => 61,
    19303 => 61,
    19304 => 61,
    19305 => 61,
    19306 => 61,
    19307 => 61,
    19308 => 61,
    19309 => 61,
    19310 => 61,
    19311 => 61,
    19312 => 61,
    19313 => 61,
    19314 => 61,
    19315 => 61,
    19316 => 61,
    19317 => 61,
    19318 => 61,
    19319 => 61,
    19320 => 61,
    19321 => 61,
    19322 => 61,
    19323 => 61,
    19324 => 61,
    19325 => 61,
    19326 => 61,
    19327 => 61,
    19328 => 61,
    19329 => 61,
    19330 => 61,
    19331 => 61,
    19332 => 61,
    19333 => 60,
    19334 => 60,
    19335 => 60,
    19336 => 60,
    19337 => 60,
    19338 => 60,
    19339 => 60,
    19340 => 60,
    19341 => 60,
    19342 => 60,
    19343 => 60,
    19344 => 60,
    19345 => 60,
    19346 => 60,
    19347 => 60,
    19348 => 60,
    19349 => 60,
    19350 => 60,
    19351 => 60,
    19352 => 60,
    19353 => 60,
    19354 => 60,
    19355 => 60,
    19356 => 60,
    19357 => 60,
    19358 => 60,
    19359 => 60,
    19360 => 60,
    19361 => 60,
    19362 => 60,
    19363 => 60,
    19364 => 60,
    19365 => 60,
    19366 => 60,
    19367 => 60,
    19368 => 60,
    19369 => 60,
    19370 => 60,
    19371 => 60,
    19372 => 60,
    19373 => 60,
    19374 => 60,
    19375 => 60,
    19376 => 60,
    19377 => 60,
    19378 => 60,
    19379 => 60,
    19380 => 60,
    19381 => 60,
    19382 => 60,
    19383 => 60,
    19384 => 60,
    19385 => 60,
    19386 => 60,
    19387 => 60,
    19388 => 60,
    19389 => 60,
    19390 => 60,
    19391 => 60,
    19392 => 60,
    19393 => 60,
    19394 => 60,
    19395 => 60,
    19396 => 60,
    19397 => 60,
    19398 => 60,
    19399 => 60,
    19400 => 60,
    19401 => 60,
    19402 => 60,
    19403 => 60,
    19404 => 60,
    19405 => 60,
    19406 => 60,
    19407 => 60,
    19408 => 60,
    19409 => 60,
    19410 => 60,
    19411 => 60,
    19412 => 60,
    19413 => 60,
    19414 => 60,
    19415 => 60,
    19416 => 60,
    19417 => 60,
    19418 => 60,
    19419 => 60,
    19420 => 60,
    19421 => 60,
    19422 => 60,
    19423 => 60,
    19424 => 60,
    19425 => 60,
    19426 => 60,
    19427 => 60,
    19428 => 60,
    19429 => 60,
    19430 => 60,
    19431 => 60,
    19432 => 60,
    19433 => 60,
    19434 => 60,
    19435 => 60,
    19436 => 60,
    19437 => 60,
    19438 => 60,
    19439 => 60,
    19440 => 60,
    19441 => 60,
    19442 => 60,
    19443 => 60,
    19444 => 60,
    19445 => 60,
    19446 => 60,
    19447 => 60,
    19448 => 60,
    19449 => 60,
    19450 => 60,
    19451 => 60,
    19452 => 60,
    19453 => 60,
    19454 => 60,
    19455 => 60,
    19456 => 60,
    19457 => 60,
    19458 => 60,
    19459 => 60,
    19460 => 60,
    19461 => 60,
    19462 => 60,
    19463 => 60,
    19464 => 60,
    19465 => 60,
    19466 => 60,
    19467 => 60,
    19468 => 60,
    19469 => 60,
    19470 => 60,
    19471 => 60,
    19472 => 60,
    19473 => 60,
    19474 => 60,
    19475 => 60,
    19476 => 60,
    19477 => 60,
    19478 => 60,
    19479 => 60,
    19480 => 60,
    19481 => 60,
    19482 => 60,
    19483 => 60,
    19484 => 60,
    19485 => 60,
    19486 => 60,
    19487 => 60,
    19488 => 60,
    19489 => 60,
    19490 => 60,
    19491 => 60,
    19492 => 60,
    19493 => 60,
    19494 => 60,
    19495 => 60,
    19496 => 60,
    19497 => 60,
    19498 => 60,
    19499 => 60,
    19500 => 60,
    19501 => 60,
    19502 => 60,
    19503 => 60,
    19504 => 60,
    19505 => 60,
    19506 => 60,
    19507 => 60,
    19508 => 60,
    19509 => 60,
    19510 => 60,
    19511 => 60,
    19512 => 60,
    19513 => 60,
    19514 => 60,
    19515 => 60,
    19516 => 60,
    19517 => 60,
    19518 => 60,
    19519 => 60,
    19520 => 60,
    19521 => 60,
    19522 => 60,
    19523 => 60,
    19524 => 60,
    19525 => 60,
    19526 => 60,
    19527 => 60,
    19528 => 60,
    19529 => 60,
    19530 => 60,
    19531 => 60,
    19532 => 60,
    19533 => 60,
    19534 => 60,
    19535 => 60,
    19536 => 60,
    19537 => 60,
    19538 => 60,
    19539 => 60,
    19540 => 60,
    19541 => 60,
    19542 => 60,
    19543 => 60,
    19544 => 60,
    19545 => 60,
    19546 => 60,
    19547 => 60,
    19548 => 60,
    19549 => 60,
    19550 => 60,
    19551 => 60,
    19552 => 60,
    19553 => 60,
    19554 => 60,
    19555 => 60,
    19556 => 60,
    19557 => 60,
    19558 => 60,
    19559 => 60,
    19560 => 60,
    19561 => 60,
    19562 => 60,
    19563 => 60,
    19564 => 60,
    19565 => 60,
    19566 => 60,
    19567 => 60,
    19568 => 60,
    19569 => 60,
    19570 => 60,
    19571 => 60,
    19572 => 60,
    19573 => 60,
    19574 => 60,
    19575 => 60,
    19576 => 60,
    19577 => 60,
    19578 => 60,
    19579 => 60,
    19580 => 60,
    19581 => 60,
    19582 => 60,
    19583 => 60,
    19584 => 60,
    19585 => 60,
    19586 => 60,
    19587 => 60,
    19588 => 60,
    19589 => 60,
    19590 => 60,
    19591 => 60,
    19592 => 60,
    19593 => 60,
    19594 => 60,
    19595 => 60,
    19596 => 60,
    19597 => 60,
    19598 => 60,
    19599 => 60,
    19600 => 60,
    19601 => 60,
    19602 => 60,
    19603 => 60,
    19604 => 60,
    19605 => 60,
    19606 => 60,
    19607 => 60,
    19608 => 60,
    19609 => 60,
    19610 => 60,
    19611 => 60,
    19612 => 60,
    19613 => 60,
    19614 => 60,
    19615 => 60,
    19616 => 60,
    19617 => 60,
    19618 => 60,
    19619 => 60,
    19620 => 60,
    19621 => 60,
    19622 => 60,
    19623 => 60,
    19624 => 60,
    19625 => 60,
    19626 => 60,
    19627 => 60,
    19628 => 60,
    19629 => 60,
    19630 => 60,
    19631 => 60,
    19632 => 60,
    19633 => 60,
    19634 => 60,
    19635 => 60,
    19636 => 60,
    19637 => 60,
    19638 => 60,
    19639 => 60,
    19640 => 60,
    19641 => 60,
    19642 => 60,
    19643 => 60,
    19644 => 60,
    19645 => 60,
    19646 => 60,
    19647 => 60,
    19648 => 60,
    19649 => 60,
    19650 => 60,
    19651 => 60,
    19652 => 60,
    19653 => 60,
    19654 => 60,
    19655 => 60,
    19656 => 60,
    19657 => 60,
    19658 => 60,
    19659 => 60,
    19660 => 60,
    19661 => 60,
    19662 => 60,
    19663 => 60,
    19664 => 60,
    19665 => 60,
    19666 => 60,
    19667 => 60,
    19668 => 60,
    19669 => 60,
    19670 => 60,
    19671 => 60,
    19672 => 60,
    19673 => 60,
    19674 => 60,
    19675 => 60,
    19676 => 60,
    19677 => 60,
    19678 => 60,
    19679 => 60,
    19680 => 60,
    19681 => 60,
    19682 => 60,
    19683 => 60,
    19684 => 60,
    19685 => 60,
    19686 => 60,
    19687 => 60,
    19688 => 60,
    19689 => 60,
    19690 => 60,
    19691 => 60,
    19692 => 60,
    19693 => 60,
    19694 => 60,
    19695 => 60,
    19696 => 60,
    19697 => 60,
    19698 => 60,
    19699 => 60,
    19700 => 60,
    19701 => 60,
    19702 => 60,
    19703 => 60,
    19704 => 60,
    19705 => 60,
    19706 => 60,
    19707 => 60,
    19708 => 60,
    19709 => 60,
    19710 => 60,
    19711 => 60,
    19712 => 60,
    19713 => 60,
    19714 => 60,
    19715 => 60,
    19716 => 60,
    19717 => 60,
    19718 => 60,
    19719 => 60,
    19720 => 60,
    19721 => 60,
    19722 => 60,
    19723 => 60,
    19724 => 60,
    19725 => 60,
    19726 => 60,
    19727 => 60,
    19728 => 60,
    19729 => 60,
    19730 => 60,
    19731 => 60,
    19732 => 60,
    19733 => 60,
    19734 => 60,
    19735 => 60,
    19736 => 60,
    19737 => 60,
    19738 => 60,
    19739 => 60,
    19740 => 60,
    19741 => 60,
    19742 => 60,
    19743 => 60,
    19744 => 60,
    19745 => 60,
    19746 => 60,
    19747 => 60,
    19748 => 60,
    19749 => 60,
    19750 => 60,
    19751 => 60,
    19752 => 60,
    19753 => 60,
    19754 => 60,
    19755 => 60,
    19756 => 60,
    19757 => 60,
    19758 => 60,
    19759 => 60,
    19760 => 60,
    19761 => 60,
    19762 => 60,
    19763 => 60,
    19764 => 60,
    19765 => 60,
    19766 => 60,
    19767 => 60,
    19768 => 60,
    19769 => 60,
    19770 => 60,
    19771 => 60,
    19772 => 60,
    19773 => 60,
    19774 => 60,
    19775 => 60,
    19776 => 60,
    19777 => 60,
    19778 => 60,
    19779 => 60,
    19780 => 60,
    19781 => 60,
    19782 => 60,
    19783 => 60,
    19784 => 60,
    19785 => 60,
    19786 => 60,
    19787 => 60,
    19788 => 60,
    19789 => 60,
    19790 => 60,
    19791 => 60,
    19792 => 60,
    19793 => 60,
    19794 => 60,
    19795 => 60,
    19796 => 60,
    19797 => 60,
    19798 => 60,
    19799 => 60,
    19800 => 60,
    19801 => 60,
    19802 => 60,
    19803 => 60,
    19804 => 60,
    19805 => 60,
    19806 => 60,
    19807 => 60,
    19808 => 60,
    19809 => 60,
    19810 => 60,
    19811 => 60,
    19812 => 60,
    19813 => 60,
    19814 => 60,
    19815 => 60,
    19816 => 60,
    19817 => 60,
    19818 => 60,
    19819 => 60,
    19820 => 60,
    19821 => 60,
    19822 => 60,
    19823 => 60,
    19824 => 60,
    19825 => 60,
    19826 => 60,
    19827 => 60,
    19828 => 60,
    19829 => 60,
    19830 => 60,
    19831 => 60,
    19832 => 60,
    19833 => 60,
    19834 => 60,
    19835 => 60,
    19836 => 60,
    19837 => 60,
    19838 => 60,
    19839 => 60,
    19840 => 60,
    19841 => 60,
    19842 => 60,
    19843 => 60,
    19844 => 60,
    19845 => 60,
    19846 => 60,
    19847 => 60,
    19848 => 60,
    19849 => 60,
    19850 => 60,
    19851 => 60,
    19852 => 60,
    19853 => 60,
    19854 => 60,
    19855 => 60,
    19856 => 60,
    19857 => 60,
    19858 => 60,
    19859 => 60,
    19860 => 60,
    19861 => 60,
    19862 => 60,
    19863 => 60,
    19864 => 60,
    19865 => 60,
    19866 => 60,
    19867 => 60,
    19868 => 60,
    19869 => 60,
    19870 => 60,
    19871 => 60,
    19872 => 60,
    19873 => 60,
    19874 => 60,
    19875 => 60,
    19876 => 60,
    19877 => 60,
    19878 => 59,
    19879 => 59,
    19880 => 59,
    19881 => 59,
    19882 => 59,
    19883 => 59,
    19884 => 59,
    19885 => 59,
    19886 => 59,
    19887 => 59,
    19888 => 59,
    19889 => 59,
    19890 => 59,
    19891 => 59,
    19892 => 59,
    19893 => 59,
    19894 => 59,
    19895 => 59,
    19896 => 59,
    19897 => 59,
    19898 => 59,
    19899 => 59,
    19900 => 59,
    19901 => 59,
    19902 => 59,
    19903 => 59,
    19904 => 59,
    19905 => 59,
    19906 => 59,
    19907 => 59,
    19908 => 59,
    19909 => 59,
    19910 => 59,
    19911 => 59,
    19912 => 59,
    19913 => 59,
    19914 => 59,
    19915 => 59,
    19916 => 59,
    19917 => 59,
    19918 => 59,
    19919 => 59,
    19920 => 59,
    19921 => 59,
    19922 => 59,
    19923 => 59,
    19924 => 59,
    19925 => 59,
    19926 => 59,
    19927 => 59,
    19928 => 59,
    19929 => 59,
    19930 => 59,
    19931 => 59,
    19932 => 59,
    19933 => 59,
    19934 => 59,
    19935 => 59,
    19936 => 59,
    19937 => 59,
    19938 => 59,
    19939 => 59,
    19940 => 59,
    19941 => 59,
    19942 => 59,
    19943 => 59,
    19944 => 59,
    19945 => 59,
    19946 => 59,
    19947 => 59,
    19948 => 59,
    19949 => 59,
    19950 => 59,
    19951 => 59,
    19952 => 59,
    19953 => 59,
    19954 => 59,
    19955 => 59,
    19956 => 59,
    19957 => 59,
    19958 => 59,
    19959 => 59,
    19960 => 59,
    19961 => 59,
    19962 => 59,
    19963 => 59,
    19964 => 59,
    19965 => 59,
    19966 => 59,
    19967 => 59,
    19968 => 59,
    19969 => 59,
    19970 => 59,
    19971 => 59,
    19972 => 59,
    19973 => 59,
    19974 => 59,
    19975 => 59,
    19976 => 59,
    19977 => 59,
    19978 => 59,
    19979 => 59,
    19980 => 59,
    19981 => 59,
    19982 => 59,
    19983 => 59,
    19984 => 59,
    19985 => 59,
    19986 => 59,
    19987 => 59,
    19988 => 59,
    19989 => 59,
    19990 => 59,
    19991 => 59,
    19992 => 59,
    19993 => 59,
    19994 => 59,
    19995 => 59,
    19996 => 59,
    19997 => 59,
    19998 => 59,
    19999 => 59,
    20000 => 59,
    20001 => 59,
    20002 => 59,
    20003 => 59,
    20004 => 59,
    20005 => 59,
    20006 => 59,
    20007 => 59,
    20008 => 59,
    20009 => 59,
    20010 => 59,
    20011 => 59,
    20012 => 59,
    20013 => 59,
    20014 => 59,
    20015 => 59,
    20016 => 59,
    20017 => 59,
    20018 => 59,
    20019 => 59,
    20020 => 59,
    20021 => 59,
    20022 => 59,
    20023 => 59,
    20024 => 59,
    20025 => 59,
    20026 => 59,
    20027 => 59,
    20028 => 59,
    20029 => 59,
    20030 => 59,
    20031 => 59,
    20032 => 59,
    20033 => 59,
    20034 => 59,
    20035 => 59,
    20036 => 59,
    20037 => 59,
    20038 => 59,
    20039 => 59,
    20040 => 59,
    20041 => 59,
    20042 => 59,
    20043 => 59,
    20044 => 59,
    20045 => 59,
    20046 => 59,
    20047 => 59,
    20048 => 59,
    20049 => 59,
    20050 => 59,
    20051 => 59,
    20052 => 59,
    20053 => 59,
    20054 => 59,
    20055 => 59,
    20056 => 59,
    20057 => 59,
    20058 => 59,
    20059 => 59,
    20060 => 59,
    20061 => 59,
    20062 => 59,
    20063 => 59,
    20064 => 59,
    20065 => 59,
    20066 => 59,
    20067 => 59,
    20068 => 59,
    20069 => 59,
    20070 => 59,
    20071 => 59,
    20072 => 59,
    20073 => 59,
    20074 => 59,
    20075 => 59,
    20076 => 59,
    20077 => 59,
    20078 => 59,
    20079 => 59,
    20080 => 59,
    20081 => 59,
    20082 => 59,
    20083 => 59,
    20084 => 59,
    20085 => 59,
    20086 => 59,
    20087 => 59,
    20088 => 59,
    20089 => 59,
    20090 => 59,
    20091 => 59,
    20092 => 59,
    20093 => 59,
    20094 => 59,
    20095 => 59,
    20096 => 59,
    20097 => 59,
    20098 => 59,
    20099 => 59,
    20100 => 59,
    20101 => 59,
    20102 => 59,
    20103 => 59,
    20104 => 59,
    20105 => 59,
    20106 => 59,
    20107 => 59,
    20108 => 59,
    20109 => 59,
    20110 => 59,
    20111 => 59,
    20112 => 59,
    20113 => 59,
    20114 => 59,
    20115 => 59,
    20116 => 59,
    20117 => 59,
    20118 => 59,
    20119 => 59,
    20120 => 59,
    20121 => 59,
    20122 => 59,
    20123 => 59,
    20124 => 59,
    20125 => 59,
    20126 => 59,
    20127 => 59,
    20128 => 59,
    20129 => 59,
    20130 => 59,
    20131 => 59,
    20132 => 59,
    20133 => 59,
    20134 => 59,
    20135 => 59,
    20136 => 59,
    20137 => 59,
    20138 => 59,
    20139 => 59,
    20140 => 59,
    20141 => 59,
    20142 => 59,
    20143 => 59,
    20144 => 59,
    20145 => 59,
    20146 => 59,
    20147 => 59,
    20148 => 59,
    20149 => 59,
    20150 => 59,
    20151 => 59,
    20152 => 59,
    20153 => 59,
    20154 => 59,
    20155 => 59,
    20156 => 59,
    20157 => 59,
    20158 => 59,
    20159 => 59,
    20160 => 59,
    20161 => 59,
    20162 => 59,
    20163 => 59,
    20164 => 59,
    20165 => 59,
    20166 => 59,
    20167 => 59,
    20168 => 59,
    20169 => 59,
    20170 => 59,
    20171 => 59,
    20172 => 59,
    20173 => 59,
    20174 => 59,
    20175 => 59,
    20176 => 59,
    20177 => 59,
    20178 => 59,
    20179 => 59,
    20180 => 59,
    20181 => 59,
    20182 => 59,
    20183 => 59,
    20184 => 59,
    20185 => 59,
    20186 => 59,
    20187 => 59,
    20188 => 59,
    20189 => 59,
    20190 => 59,
    20191 => 59,
    20192 => 59,
    20193 => 59,
    20194 => 59,
    20195 => 59,
    20196 => 59,
    20197 => 59,
    20198 => 59,
    20199 => 59,
    20200 => 59,
    20201 => 59,
    20202 => 59,
    20203 => 59,
    20204 => 59,
    20205 => 59,
    20206 => 59,
    20207 => 59,
    20208 => 59,
    20209 => 59,
    20210 => 59,
    20211 => 59,
    20212 => 59,
    20213 => 59,
    20214 => 59,
    20215 => 59,
    20216 => 59,
    20217 => 59,
    20218 => 59,
    20219 => 59,
    20220 => 59,
    20221 => 59,
    20222 => 59,
    20223 => 59,
    20224 => 59,
    20225 => 59,
    20226 => 59,
    20227 => 59,
    20228 => 59,
    20229 => 59,
    20230 => 59,
    20231 => 59,
    20232 => 59,
    20233 => 59,
    20234 => 59,
    20235 => 59,
    20236 => 59,
    20237 => 59,
    20238 => 59,
    20239 => 59,
    20240 => 59,
    20241 => 59,
    20242 => 59,
    20243 => 59,
    20244 => 59,
    20245 => 59,
    20246 => 59,
    20247 => 59,
    20248 => 59,
    20249 => 59,
    20250 => 59,
    20251 => 59,
    20252 => 59,
    20253 => 59,
    20254 => 59,
    20255 => 59,
    20256 => 59,
    20257 => 59,
    20258 => 59,
    20259 => 59,
    20260 => 59,
    20261 => 59,
    20262 => 59,
    20263 => 59,
    20264 => 59,
    20265 => 59,
    20266 => 59,
    20267 => 59,
    20268 => 59,
    20269 => 59,
    20270 => 59,
    20271 => 59,
    20272 => 59,
    20273 => 59,
    20274 => 59,
    20275 => 59,
    20276 => 59,
    20277 => 59,
    20278 => 59,
    20279 => 59,
    20280 => 59,
    20281 => 59,
    20282 => 59,
    20283 => 59,
    20284 => 59,
    20285 => 59,
    20286 => 59,
    20287 => 59,
    20288 => 59,
    20289 => 59,
    20290 => 59,
    20291 => 59,
    20292 => 59,
    20293 => 59,
    20294 => 59,
    20295 => 59,
    20296 => 59,
    20297 => 59,
    20298 => 59,
    20299 => 59,
    20300 => 59,
    20301 => 59,
    20302 => 59,
    20303 => 59,
    20304 => 59,
    20305 => 59,
    20306 => 59,
    20307 => 59,
    20308 => 59,
    20309 => 59,
    20310 => 59,
    20311 => 59,
    20312 => 59,
    20313 => 59,
    20314 => 59,
    20315 => 59,
    20316 => 59,
    20317 => 59,
    20318 => 59,
    20319 => 59,
    20320 => 59,
    20321 => 59,
    20322 => 59,
    20323 => 59,
    20324 => 59,
    20325 => 59,
    20326 => 59,
    20327 => 59,
    20328 => 59,
    20329 => 59,
    20330 => 59,
    20331 => 59,
    20332 => 59,
    20333 => 59,
    20334 => 59,
    20335 => 59,
    20336 => 59,
    20337 => 59,
    20338 => 59,
    20339 => 59,
    20340 => 59,
    20341 => 59,
    20342 => 59,
    20343 => 59,
    20344 => 59,
    20345 => 59,
    20346 => 59,
    20347 => 59,
    20348 => 59,
    20349 => 59,
    20350 => 59,
    20351 => 58,
    20352 => 58,
    20353 => 58,
    20354 => 58,
    20355 => 58,
    20356 => 58,
    20357 => 58,
    20358 => 58,
    20359 => 58,
    20360 => 58,
    20361 => 58,
    20362 => 58,
    20363 => 58,
    20364 => 58,
    20365 => 58,
    20366 => 58,
    20367 => 58,
    20368 => 58,
    20369 => 58,
    20370 => 58,
    20371 => 58,
    20372 => 58,
    20373 => 58,
    20374 => 58,
    20375 => 58,
    20376 => 58,
    20377 => 58,
    20378 => 58,
    20379 => 58,
    20380 => 58,
    20381 => 58,
    20382 => 58,
    20383 => 58,
    20384 => 58,
    20385 => 58,
    20386 => 58,
    20387 => 58,
    20388 => 58,
    20389 => 58,
    20390 => 58,
    20391 => 58,
    20392 => 58,
    20393 => 58,
    20394 => 58,
    20395 => 58,
    20396 => 58,
    20397 => 58,
    20398 => 58,
    20399 => 58,
    20400 => 58,
    20401 => 58,
    20402 => 58,
    20403 => 58,
    20404 => 58,
    20405 => 58,
    20406 => 58,
    20407 => 58,
    20408 => 58,
    20409 => 58,
    20410 => 58,
    20411 => 58,
    20412 => 58,
    20413 => 58,
    20414 => 58,
    20415 => 58,
    20416 => 58,
    20417 => 58,
    20418 => 58,
    20419 => 58,
    20420 => 58,
    20421 => 58,
    20422 => 58,
    20423 => 58,
    20424 => 58,
    20425 => 58,
    20426 => 58,
    20427 => 58,
    20428 => 58,
    20429 => 58,
    20430 => 58,
    20431 => 58,
    20432 => 58,
    20433 => 58,
    20434 => 58,
    20435 => 58,
    20436 => 58,
    20437 => 58,
    20438 => 58,
    20439 => 58,
    20440 => 58,
    20441 => 58,
    20442 => 58,
    20443 => 58,
    20444 => 58,
    20445 => 58,
    20446 => 58,
    20447 => 58,
    20448 => 58,
    20449 => 58,
    20450 => 58,
    20451 => 58,
    20452 => 58,
    20453 => 58,
    20454 => 58,
    20455 => 58,
    20456 => 58,
    20457 => 58,
    20458 => 58,
    20459 => 58,
    20460 => 58,
    20461 => 58,
    20462 => 58,
    20463 => 58,
    20464 => 58,
    20465 => 58,
    20466 => 58,
    20467 => 58,
    20468 => 58,
    20469 => 58,
    20470 => 58,
    20471 => 58,
    20472 => 58,
    20473 => 58,
    20474 => 58,
    20475 => 58,
    20476 => 58,
    20477 => 58,
    20478 => 58,
    20479 => 58,
    20480 => 58,
    20481 => 58,
    20482 => 58,
    20483 => 58,
    20484 => 58,
    20485 => 58,
    20486 => 58,
    20487 => 58,
    20488 => 58,
    20489 => 58,
    20490 => 58,
    20491 => 58,
    20492 => 58,
    20493 => 58,
    20494 => 58,
    20495 => 58,
    20496 => 58,
    20497 => 58,
    20498 => 58,
    20499 => 58,
    20500 => 58,
    20501 => 58,
    20502 => 58,
    20503 => 58,
    20504 => 58,
    20505 => 58,
    20506 => 58,
    20507 => 58,
    20508 => 58,
    20509 => 58,
    20510 => 58,
    20511 => 58,
    20512 => 58,
    20513 => 58,
    20514 => 58,
    20515 => 58,
    20516 => 58,
    20517 => 58,
    20518 => 58,
    20519 => 58,
    20520 => 58,
    20521 => 58,
    20522 => 58,
    20523 => 58,
    20524 => 58,
    20525 => 58,
    20526 => 58,
    20527 => 58,
    20528 => 58,
    20529 => 58,
    20530 => 58,
    20531 => 58,
    20532 => 58,
    20533 => 58,
    20534 => 58,
    20535 => 58,
    20536 => 58,
    20537 => 58,
    20538 => 58,
    20539 => 58,
    20540 => 58,
    20541 => 58,
    20542 => 58,
    20543 => 58,
    20544 => 58,
    20545 => 58,
    20546 => 58,
    20547 => 58,
    20548 => 58,
    20549 => 58,
    20550 => 58,
    20551 => 58,
    20552 => 58,
    20553 => 58,
    20554 => 58,
    20555 => 58,
    20556 => 58,
    20557 => 58,
    20558 => 58,
    20559 => 58,
    20560 => 58,
    20561 => 58,
    20562 => 58,
    20563 => 58,
    20564 => 58,
    20565 => 58,
    20566 => 58,
    20567 => 58,
    20568 => 58,
    20569 => 58,
    20570 => 58,
    20571 => 58,
    20572 => 58,
    20573 => 58,
    20574 => 58,
    20575 => 58,
    20576 => 58,
    20577 => 58,
    20578 => 58,
    20579 => 58,
    20580 => 58,
    20581 => 58,
    20582 => 58,
    20583 => 58,
    20584 => 58,
    20585 => 58,
    20586 => 58,
    20587 => 58,
    20588 => 58,
    20589 => 58,
    20590 => 58,
    20591 => 58,
    20592 => 58,
    20593 => 58,
    20594 => 58,
    20595 => 58,
    20596 => 58,
    20597 => 58,
    20598 => 58,
    20599 => 58,
    20600 => 58,
    20601 => 58,
    20602 => 58,
    20603 => 58,
    20604 => 58,
    20605 => 58,
    20606 => 58,
    20607 => 58,
    20608 => 58,
    20609 => 58,
    20610 => 58,
    20611 => 58,
    20612 => 58,
    20613 => 58,
    20614 => 58,
    20615 => 58,
    20616 => 58,
    20617 => 58,
    20618 => 58,
    20619 => 58,
    20620 => 58,
    20621 => 58,
    20622 => 58,
    20623 => 58,
    20624 => 58,
    20625 => 58,
    20626 => 58,
    20627 => 58,
    20628 => 58,
    20629 => 58,
    20630 => 58,
    20631 => 58,
    20632 => 58,
    20633 => 58,
    20634 => 58,
    20635 => 58,
    20636 => 58,
    20637 => 58,
    20638 => 58,
    20639 => 58,
    20640 => 58,
    20641 => 58,
    20642 => 58,
    20643 => 58,
    20644 => 58,
    20645 => 58,
    20646 => 58,
    20647 => 58,
    20648 => 58,
    20649 => 58,
    20650 => 58,
    20651 => 58,
    20652 => 58,
    20653 => 58,
    20654 => 58,
    20655 => 58,
    20656 => 58,
    20657 => 58,
    20658 => 58,
    20659 => 58,
    20660 => 58,
    20661 => 58,
    20662 => 58,
    20663 => 58,
    20664 => 58,
    20665 => 58,
    20666 => 58,
    20667 => 58,
    20668 => 58,
    20669 => 58,
    20670 => 58,
    20671 => 58,
    20672 => 58,
    20673 => 58,
    20674 => 58,
    20675 => 58,
    20676 => 58,
    20677 => 58,
    20678 => 58,
    20679 => 58,
    20680 => 58,
    20681 => 58,
    20682 => 58,
    20683 => 58,
    20684 => 58,
    20685 => 58,
    20686 => 58,
    20687 => 58,
    20688 => 58,
    20689 => 58,
    20690 => 58,
    20691 => 58,
    20692 => 58,
    20693 => 58,
    20694 => 58,
    20695 => 58,
    20696 => 58,
    20697 => 58,
    20698 => 58,
    20699 => 58,
    20700 => 58,
    20701 => 58,
    20702 => 58,
    20703 => 58,
    20704 => 58,
    20705 => 58,
    20706 => 58,
    20707 => 58,
    20708 => 58,
    20709 => 58,
    20710 => 58,
    20711 => 58,
    20712 => 58,
    20713 => 58,
    20714 => 58,
    20715 => 58,
    20716 => 58,
    20717 => 58,
    20718 => 58,
    20719 => 58,
    20720 => 58,
    20721 => 58,
    20722 => 58,
    20723 => 58,
    20724 => 58,
    20725 => 58,
    20726 => 58,
    20727 => 58,
    20728 => 58,
    20729 => 58,
    20730 => 58,
    20731 => 58,
    20732 => 58,
    20733 => 58,
    20734 => 58,
    20735 => 58,
    20736 => 58,
    20737 => 58,
    20738 => 58,
    20739 => 58,
    20740 => 58,
    20741 => 58,
    20742 => 58,
    20743 => 58,
    20744 => 58,
    20745 => 58,
    20746 => 58,
    20747 => 58,
    20748 => 58,
    20749 => 58,
    20750 => 58,
    20751 => 58,
    20752 => 58,
    20753 => 58,
    20754 => 58,
    20755 => 58,
    20756 => 58,
    20757 => 58,
    20758 => 58,
    20759 => 58,
    20760 => 58,
    20761 => 58,
    20762 => 58,
    20763 => 58,
    20764 => 58,
    20765 => 58,
    20766 => 58,
    20767 => 58,
    20768 => 58,
    20769 => 58,
    20770 => 58,
    20771 => 58,
    20772 => 58,
    20773 => 58,
    20774 => 58,
    20775 => 57,
    20776 => 57,
    20777 => 57,
    20778 => 57,
    20779 => 57,
    20780 => 57,
    20781 => 57,
    20782 => 57,
    20783 => 57,
    20784 => 57,
    20785 => 57,
    20786 => 57,
    20787 => 57,
    20788 => 57,
    20789 => 57,
    20790 => 57,
    20791 => 57,
    20792 => 57,
    20793 => 57,
    20794 => 57,
    20795 => 57,
    20796 => 57,
    20797 => 57,
    20798 => 57,
    20799 => 57,
    20800 => 57,
    20801 => 57,
    20802 => 57,
    20803 => 57,
    20804 => 57,
    20805 => 57,
    20806 => 57,
    20807 => 57,
    20808 => 57,
    20809 => 57,
    20810 => 57,
    20811 => 57,
    20812 => 57,
    20813 => 57,
    20814 => 57,
    20815 => 57,
    20816 => 57,
    20817 => 57,
    20818 => 57,
    20819 => 57,
    20820 => 57,
    20821 => 57,
    20822 => 57,
    20823 => 57,
    20824 => 57,
    20825 => 57,
    20826 => 57,
    20827 => 57,
    20828 => 57,
    20829 => 57,
    20830 => 57,
    20831 => 57,
    20832 => 57,
    20833 => 57,
    20834 => 57,
    20835 => 57,
    20836 => 57,
    20837 => 57,
    20838 => 57,
    20839 => 57,
    20840 => 57,
    20841 => 57,
    20842 => 57,
    20843 => 57,
    20844 => 57,
    20845 => 57,
    20846 => 57,
    20847 => 57,
    20848 => 57,
    20849 => 57,
    20850 => 57,
    20851 => 57,
    20852 => 57,
    20853 => 57,
    20854 => 57,
    20855 => 57,
    20856 => 57,
    20857 => 57,
    20858 => 57,
    20859 => 57,
    20860 => 57,
    20861 => 57,
    20862 => 57,
    20863 => 57,
    20864 => 57,
    20865 => 57,
    20866 => 57,
    20867 => 57,
    20868 => 57,
    20869 => 57,
    20870 => 57,
    20871 => 57,
    20872 => 57,
    20873 => 57,
    20874 => 57,
    20875 => 57,
    20876 => 57,
    20877 => 57,
    20878 => 57,
    20879 => 57,
    20880 => 57,
    20881 => 57,
    20882 => 57,
    20883 => 57,
    20884 => 57,
    20885 => 57,
    20886 => 57,
    20887 => 57,
    20888 => 57,
    20889 => 57,
    20890 => 57,
    20891 => 57,
    20892 => 57,
    20893 => 57,
    20894 => 57,
    20895 => 57,
    20896 => 57,
    20897 => 57,
    20898 => 57,
    20899 => 57,
    20900 => 57,
    20901 => 57,
    20902 => 57,
    20903 => 57,
    20904 => 57,
    20905 => 57,
    20906 => 57,
    20907 => 57,
    20908 => 57,
    20909 => 57,
    20910 => 57,
    20911 => 57,
    20912 => 57,
    20913 => 57,
    20914 => 57,
    20915 => 57,
    20916 => 57,
    20917 => 57,
    20918 => 57,
    20919 => 57,
    20920 => 57,
    20921 => 57,
    20922 => 57,
    20923 => 57,
    20924 => 57,
    20925 => 57,
    20926 => 57,
    20927 => 57,
    20928 => 57,
    20929 => 57,
    20930 => 57,
    20931 => 57,
    20932 => 57,
    20933 => 57,
    20934 => 57,
    20935 => 57,
    20936 => 57,
    20937 => 57,
    20938 => 57,
    20939 => 57,
    20940 => 57,
    20941 => 57,
    20942 => 57,
    20943 => 57,
    20944 => 57,
    20945 => 57,
    20946 => 57,
    20947 => 57,
    20948 => 57,
    20949 => 57,
    20950 => 57,
    20951 => 57,
    20952 => 57,
    20953 => 57,
    20954 => 57,
    20955 => 57,
    20956 => 57,
    20957 => 57,
    20958 => 57,
    20959 => 57,
    20960 => 57,
    20961 => 57,
    20962 => 57,
    20963 => 57,
    20964 => 57,
    20965 => 57,
    20966 => 57,
    20967 => 57,
    20968 => 57,
    20969 => 57,
    20970 => 57,
    20971 => 57,
    20972 => 57,
    20973 => 57,
    20974 => 57,
    20975 => 57,
    20976 => 57,
    20977 => 57,
    20978 => 57,
    20979 => 57,
    20980 => 57,
    20981 => 57,
    20982 => 57,
    20983 => 57,
    20984 => 57,
    20985 => 57,
    20986 => 57,
    20987 => 57,
    20988 => 57,
    20989 => 57,
    20990 => 57,
    20991 => 57,
    20992 => 57,
    20993 => 57,
    20994 => 57,
    20995 => 57,
    20996 => 57,
    20997 => 57,
    20998 => 57,
    20999 => 57,
    21000 => 57,
    21001 => 57,
    21002 => 57,
    21003 => 57,
    21004 => 57,
    21005 => 57,
    21006 => 57,
    21007 => 57,
    21008 => 57,
    21009 => 57,
    21010 => 57,
    21011 => 57,
    21012 => 57,
    21013 => 57,
    21014 => 57,
    21015 => 57,
    21016 => 57,
    21017 => 57,
    21018 => 57,
    21019 => 57,
    21020 => 57,
    21021 => 57,
    21022 => 57,
    21023 => 57,
    21024 => 57,
    21025 => 57,
    21026 => 57,
    21027 => 57,
    21028 => 57,
    21029 => 57,
    21030 => 57,
    21031 => 57,
    21032 => 57,
    21033 => 57,
    21034 => 57,
    21035 => 57,
    21036 => 57,
    21037 => 57,
    21038 => 57,
    21039 => 57,
    21040 => 57,
    21041 => 57,
    21042 => 57,
    21043 => 57,
    21044 => 57,
    21045 => 57,
    21046 => 57,
    21047 => 57,
    21048 => 57,
    21049 => 57,
    21050 => 57,
    21051 => 57,
    21052 => 57,
    21053 => 57,
    21054 => 57,
    21055 => 57,
    21056 => 57,
    21057 => 57,
    21058 => 57,
    21059 => 57,
    21060 => 57,
    21061 => 57,
    21062 => 57,
    21063 => 57,
    21064 => 57,
    21065 => 57,
    21066 => 57,
    21067 => 57,
    21068 => 57,
    21069 => 57,
    21070 => 57,
    21071 => 57,
    21072 => 57,
    21073 => 57,
    21074 => 57,
    21075 => 57,
    21076 => 57,
    21077 => 57,
    21078 => 57,
    21079 => 57,
    21080 => 57,
    21081 => 57,
    21082 => 57,
    21083 => 57,
    21084 => 57,
    21085 => 57,
    21086 => 57,
    21087 => 57,
    21088 => 57,
    21089 => 57,
    21090 => 57,
    21091 => 57,
    21092 => 57,
    21093 => 57,
    21094 => 57,
    21095 => 57,
    21096 => 57,
    21097 => 57,
    21098 => 57,
    21099 => 57,
    21100 => 57,
    21101 => 57,
    21102 => 57,
    21103 => 57,
    21104 => 57,
    21105 => 57,
    21106 => 57,
    21107 => 57,
    21108 => 57,
    21109 => 57,
    21110 => 57,
    21111 => 57,
    21112 => 57,
    21113 => 57,
    21114 => 57,
    21115 => 57,
    21116 => 57,
    21117 => 57,
    21118 => 57,
    21119 => 57,
    21120 => 57,
    21121 => 57,
    21122 => 57,
    21123 => 57,
    21124 => 57,
    21125 => 57,
    21126 => 57,
    21127 => 57,
    21128 => 57,
    21129 => 57,
    21130 => 57,
    21131 => 57,
    21132 => 57,
    21133 => 57,
    21134 => 57,
    21135 => 57,
    21136 => 57,
    21137 => 57,
    21138 => 57,
    21139 => 57,
    21140 => 57,
    21141 => 57,
    21142 => 57,
    21143 => 57,
    21144 => 57,
    21145 => 57,
    21146 => 57,
    21147 => 57,
    21148 => 57,
    21149 => 57,
    21150 => 57,
    21151 => 57,
    21152 => 57,
    21153 => 57,
    21154 => 57,
    21155 => 57,
    21156 => 57,
    21157 => 57,
    21158 => 57,
    21159 => 57,
    21160 => 57,
    21161 => 57,
    21162 => 57,
    21163 => 57,
    21164 => 56,
    21165 => 56,
    21166 => 56,
    21167 => 56,
    21168 => 56,
    21169 => 56,
    21170 => 56,
    21171 => 56,
    21172 => 56,
    21173 => 56,
    21174 => 56,
    21175 => 56,
    21176 => 56,
    21177 => 56,
    21178 => 56,
    21179 => 56,
    21180 => 56,
    21181 => 56,
    21182 => 56,
    21183 => 56,
    21184 => 56,
    21185 => 56,
    21186 => 56,
    21187 => 56,
    21188 => 56,
    21189 => 56,
    21190 => 56,
    21191 => 56,
    21192 => 56,
    21193 => 56,
    21194 => 56,
    21195 => 56,
    21196 => 56,
    21197 => 56,
    21198 => 56,
    21199 => 56,
    21200 => 56,
    21201 => 56,
    21202 => 56,
    21203 => 56,
    21204 => 56,
    21205 => 56,
    21206 => 56,
    21207 => 56,
    21208 => 56,
    21209 => 56,
    21210 => 56,
    21211 => 56,
    21212 => 56,
    21213 => 56,
    21214 => 56,
    21215 => 56,
    21216 => 56,
    21217 => 56,
    21218 => 56,
    21219 => 56,
    21220 => 56,
    21221 => 56,
    21222 => 56,
    21223 => 56,
    21224 => 56,
    21225 => 56,
    21226 => 56,
    21227 => 56,
    21228 => 56,
    21229 => 56,
    21230 => 56,
    21231 => 56,
    21232 => 56,
    21233 => 56,
    21234 => 56,
    21235 => 56,
    21236 => 56,
    21237 => 56,
    21238 => 56,
    21239 => 56,
    21240 => 56,
    21241 => 56,
    21242 => 56,
    21243 => 56,
    21244 => 56,
    21245 => 56,
    21246 => 56,
    21247 => 56,
    21248 => 56,
    21249 => 56,
    21250 => 56,
    21251 => 56,
    21252 => 56,
    21253 => 56,
    21254 => 56,
    21255 => 56,
    21256 => 56,
    21257 => 56,
    21258 => 56,
    21259 => 56,
    21260 => 56,
    21261 => 56,
    21262 => 56,
    21263 => 56,
    21264 => 56,
    21265 => 56,
    21266 => 56,
    21267 => 56,
    21268 => 56,
    21269 => 56,
    21270 => 56,
    21271 => 56,
    21272 => 56,
    21273 => 56,
    21274 => 56,
    21275 => 56,
    21276 => 56,
    21277 => 56,
    21278 => 56,
    21279 => 56,
    21280 => 56,
    21281 => 56,
    21282 => 56,
    21283 => 56,
    21284 => 56,
    21285 => 56,
    21286 => 56,
    21287 => 56,
    21288 => 56,
    21289 => 56,
    21290 => 56,
    21291 => 56,
    21292 => 56,
    21293 => 56,
    21294 => 56,
    21295 => 56,
    21296 => 56,
    21297 => 56,
    21298 => 56,
    21299 => 56,
    21300 => 56,
    21301 => 56,
    21302 => 56,
    21303 => 56,
    21304 => 56,
    21305 => 56,
    21306 => 56,
    21307 => 56,
    21308 => 56,
    21309 => 56,
    21310 => 56,
    21311 => 56,
    21312 => 56,
    21313 => 56,
    21314 => 56,
    21315 => 56,
    21316 => 56,
    21317 => 56,
    21318 => 56,
    21319 => 56,
    21320 => 56,
    21321 => 56,
    21322 => 56,
    21323 => 56,
    21324 => 56,
    21325 => 56,
    21326 => 56,
    21327 => 56,
    21328 => 56,
    21329 => 56,
    21330 => 56,
    21331 => 56,
    21332 => 56,
    21333 => 56,
    21334 => 56,
    21335 => 56,
    21336 => 56,
    21337 => 56,
    21338 => 56,
    21339 => 56,
    21340 => 56,
    21341 => 56,
    21342 => 56,
    21343 => 56,
    21344 => 56,
    21345 => 56,
    21346 => 56,
    21347 => 56,
    21348 => 56,
    21349 => 56,
    21350 => 56,
    21351 => 56,
    21352 => 56,
    21353 => 56,
    21354 => 56,
    21355 => 56,
    21356 => 56,
    21357 => 56,
    21358 => 56,
    21359 => 56,
    21360 => 56,
    21361 => 56,
    21362 => 56,
    21363 => 56,
    21364 => 56,
    21365 => 56,
    21366 => 56,
    21367 => 56,
    21368 => 56,
    21369 => 56,
    21370 => 56,
    21371 => 56,
    21372 => 56,
    21373 => 56,
    21374 => 56,
    21375 => 56,
    21376 => 56,
    21377 => 56,
    21378 => 56,
    21379 => 56,
    21380 => 56,
    21381 => 56,
    21382 => 56,
    21383 => 56,
    21384 => 56,
    21385 => 56,
    21386 => 56,
    21387 => 56,
    21388 => 56,
    21389 => 56,
    21390 => 56,
    21391 => 56,
    21392 => 56,
    21393 => 56,
    21394 => 56,
    21395 => 56,
    21396 => 56,
    21397 => 56,
    21398 => 56,
    21399 => 56,
    21400 => 56,
    21401 => 56,
    21402 => 56,
    21403 => 56,
    21404 => 56,
    21405 => 56,
    21406 => 56,
    21407 => 56,
    21408 => 56,
    21409 => 56,
    21410 => 56,
    21411 => 56,
    21412 => 56,
    21413 => 56,
    21414 => 56,
    21415 => 56,
    21416 => 56,
    21417 => 56,
    21418 => 56,
    21419 => 56,
    21420 => 56,
    21421 => 56,
    21422 => 56,
    21423 => 56,
    21424 => 56,
    21425 => 56,
    21426 => 56,
    21427 => 56,
    21428 => 56,
    21429 => 56,
    21430 => 56,
    21431 => 56,
    21432 => 56,
    21433 => 56,
    21434 => 56,
    21435 => 56,
    21436 => 56,
    21437 => 56,
    21438 => 56,
    21439 => 56,
    21440 => 56,
    21441 => 56,
    21442 => 56,
    21443 => 56,
    21444 => 56,
    21445 => 56,
    21446 => 56,
    21447 => 56,
    21448 => 56,
    21449 => 56,
    21450 => 56,
    21451 => 56,
    21452 => 56,
    21453 => 56,
    21454 => 56,
    21455 => 56,
    21456 => 56,
    21457 => 56,
    21458 => 56,
    21459 => 56,
    21460 => 56,
    21461 => 56,
    21462 => 56,
    21463 => 56,
    21464 => 56,
    21465 => 56,
    21466 => 56,
    21467 => 56,
    21468 => 56,
    21469 => 56,
    21470 => 56,
    21471 => 56,
    21472 => 56,
    21473 => 56,
    21474 => 56,
    21475 => 56,
    21476 => 56,
    21477 => 56,
    21478 => 56,
    21479 => 56,
    21480 => 56,
    21481 => 56,
    21482 => 56,
    21483 => 56,
    21484 => 56,
    21485 => 56,
    21486 => 56,
    21487 => 56,
    21488 => 56,
    21489 => 56,
    21490 => 56,
    21491 => 56,
    21492 => 56,
    21493 => 56,
    21494 => 56,
    21495 => 56,
    21496 => 56,
    21497 => 56,
    21498 => 56,
    21499 => 56,
    21500 => 56,
    21501 => 56,
    21502 => 56,
    21503 => 56,
    21504 => 56,
    21505 => 56,
    21506 => 56,
    21507 => 56,
    21508 => 56,
    21509 => 56,
    21510 => 56,
    21511 => 56,
    21512 => 56,
    21513 => 56,
    21514 => 56,
    21515 => 56,
    21516 => 56,
    21517 => 56,
    21518 => 56,
    21519 => 56,
    21520 => 56,
    21521 => 56,
    21522 => 56,
    21523 => 56,
    21524 => 56,
    21525 => 56,
    21526 => 55,
    21527 => 55,
    21528 => 55,
    21529 => 55,
    21530 => 55,
    21531 => 55,
    21532 => 55,
    21533 => 55,
    21534 => 55,
    21535 => 55,
    21536 => 55,
    21537 => 55,
    21538 => 55,
    21539 => 55,
    21540 => 55,
    21541 => 55,
    21542 => 55,
    21543 => 55,
    21544 => 55,
    21545 => 55,
    21546 => 55,
    21547 => 55,
    21548 => 55,
    21549 => 55,
    21550 => 55,
    21551 => 55,
    21552 => 55,
    21553 => 55,
    21554 => 55,
    21555 => 55,
    21556 => 55,
    21557 => 55,
    21558 => 55,
    21559 => 55,
    21560 => 55,
    21561 => 55,
    21562 => 55,
    21563 => 55,
    21564 => 55,
    21565 => 55,
    21566 => 55,
    21567 => 55,
    21568 => 55,
    21569 => 55,
    21570 => 55,
    21571 => 55,
    21572 => 55,
    21573 => 55,
    21574 => 55,
    21575 => 55,
    21576 => 55,
    21577 => 55,
    21578 => 55,
    21579 => 55,
    21580 => 55,
    21581 => 55,
    21582 => 55,
    21583 => 55,
    21584 => 55,
    21585 => 55,
    21586 => 55,
    21587 => 55,
    21588 => 55,
    21589 => 55,
    21590 => 55,
    21591 => 55,
    21592 => 55,
    21593 => 55,
    21594 => 55,
    21595 => 55,
    21596 => 55,
    21597 => 55,
    21598 => 55,
    21599 => 55,
    21600 => 55,
    21601 => 55,
    21602 => 55,
    21603 => 55,
    21604 => 55,
    21605 => 55,
    21606 => 55,
    21607 => 55,
    21608 => 55,
    21609 => 55,
    21610 => 55,
    21611 => 55,
    21612 => 55,
    21613 => 55,
    21614 => 55,
    21615 => 55,
    21616 => 55,
    21617 => 55,
    21618 => 55,
    21619 => 55,
    21620 => 55,
    21621 => 55,
    21622 => 55,
    21623 => 55,
    21624 => 55,
    21625 => 55,
    21626 => 55,
    21627 => 55,
    21628 => 55,
    21629 => 55,
    21630 => 55,
    21631 => 55,
    21632 => 55,
    21633 => 55,
    21634 => 55,
    21635 => 55,
    21636 => 55,
    21637 => 55,
    21638 => 55,
    21639 => 55,
    21640 => 55,
    21641 => 55,
    21642 => 55,
    21643 => 55,
    21644 => 55,
    21645 => 55,
    21646 => 55,
    21647 => 55,
    21648 => 55,
    21649 => 55,
    21650 => 55,
    21651 => 55,
    21652 => 55,
    21653 => 55,
    21654 => 55,
    21655 => 55,
    21656 => 55,
    21657 => 55,
    21658 => 55,
    21659 => 55,
    21660 => 55,
    21661 => 55,
    21662 => 55,
    21663 => 55,
    21664 => 55,
    21665 => 55,
    21666 => 55,
    21667 => 55,
    21668 => 55,
    21669 => 55,
    21670 => 55,
    21671 => 55,
    21672 => 55,
    21673 => 55,
    21674 => 55,
    21675 => 55,
    21676 => 55,
    21677 => 55,
    21678 => 55,
    21679 => 55,
    21680 => 55,
    21681 => 55,
    21682 => 55,
    21683 => 55,
    21684 => 55,
    21685 => 55,
    21686 => 55,
    21687 => 55,
    21688 => 55,
    21689 => 55,
    21690 => 55,
    21691 => 55,
    21692 => 55,
    21693 => 55,
    21694 => 55,
    21695 => 55,
    21696 => 55,
    21697 => 55,
    21698 => 55,
    21699 => 55,
    21700 => 55,
    21701 => 55,
    21702 => 55,
    21703 => 55,
    21704 => 55,
    21705 => 55,
    21706 => 55,
    21707 => 55,
    21708 => 55,
    21709 => 55,
    21710 => 55,
    21711 => 55,
    21712 => 55,
    21713 => 55,
    21714 => 55,
    21715 => 55,
    21716 => 55,
    21717 => 55,
    21718 => 55,
    21719 => 55,
    21720 => 55,
    21721 => 55,
    21722 => 55,
    21723 => 55,
    21724 => 55,
    21725 => 55,
    21726 => 55,
    21727 => 55,
    21728 => 55,
    21729 => 55,
    21730 => 55,
    21731 => 55,
    21732 => 55,
    21733 => 55,
    21734 => 55,
    21735 => 55,
    21736 => 55,
    21737 => 55,
    21738 => 55,
    21739 => 55,
    21740 => 55,
    21741 => 55,
    21742 => 55,
    21743 => 55,
    21744 => 55,
    21745 => 55,
    21746 => 55,
    21747 => 55,
    21748 => 55,
    21749 => 55,
    21750 => 55,
    21751 => 55,
    21752 => 55,
    21753 => 55,
    21754 => 55,
    21755 => 55,
    21756 => 55,
    21757 => 55,
    21758 => 55,
    21759 => 55,
    21760 => 55,
    21761 => 55,
    21762 => 55,
    21763 => 55,
    21764 => 55,
    21765 => 55,
    21766 => 55,
    21767 => 55,
    21768 => 55,
    21769 => 55,
    21770 => 55,
    21771 => 55,
    21772 => 55,
    21773 => 55,
    21774 => 55,
    21775 => 55,
    21776 => 55,
    21777 => 55,
    21778 => 55,
    21779 => 55,
    21780 => 55,
    21781 => 55,
    21782 => 55,
    21783 => 55,
    21784 => 55,
    21785 => 55,
    21786 => 55,
    21787 => 55,
    21788 => 55,
    21789 => 55,
    21790 => 55,
    21791 => 55,
    21792 => 55,
    21793 => 55,
    21794 => 55,
    21795 => 55,
    21796 => 55,
    21797 => 55,
    21798 => 55,
    21799 => 55,
    21800 => 55,
    21801 => 55,
    21802 => 55,
    21803 => 55,
    21804 => 55,
    21805 => 55,
    21806 => 55,
    21807 => 55,
    21808 => 55,
    21809 => 55,
    21810 => 55,
    21811 => 55,
    21812 => 55,
    21813 => 55,
    21814 => 55,
    21815 => 55,
    21816 => 55,
    21817 => 55,
    21818 => 55,
    21819 => 55,
    21820 => 55,
    21821 => 55,
    21822 => 55,
    21823 => 55,
    21824 => 55,
    21825 => 55,
    21826 => 55,
    21827 => 55,
    21828 => 55,
    21829 => 55,
    21830 => 55,
    21831 => 55,
    21832 => 55,
    21833 => 55,
    21834 => 55,
    21835 => 55,
    21836 => 55,
    21837 => 55,
    21838 => 55,
    21839 => 55,
    21840 => 55,
    21841 => 55,
    21842 => 55,
    21843 => 55,
    21844 => 55,
    21845 => 55,
    21846 => 55,
    21847 => 55,
    21848 => 55,
    21849 => 55,
    21850 => 55,
    21851 => 55,
    21852 => 55,
    21853 => 55,
    21854 => 55,
    21855 => 55,
    21856 => 55,
    21857 => 55,
    21858 => 55,
    21859 => 55,
    21860 => 55,
    21861 => 55,
    21862 => 55,
    21863 => 55,
    21864 => 55,
    21865 => 55,
    21866 => 54,
    21867 => 54,
    21868 => 54,
    21869 => 54,
    21870 => 54,
    21871 => 54,
    21872 => 54,
    21873 => 54,
    21874 => 54,
    21875 => 54,
    21876 => 54,
    21877 => 54,
    21878 => 54,
    21879 => 54,
    21880 => 54,
    21881 => 54,
    21882 => 54,
    21883 => 54,
    21884 => 54,
    21885 => 54,
    21886 => 54,
    21887 => 54,
    21888 => 54,
    21889 => 54,
    21890 => 54,
    21891 => 54,
    21892 => 54,
    21893 => 54,
    21894 => 54,
    21895 => 54,
    21896 => 54,
    21897 => 54,
    21898 => 54,
    21899 => 54,
    21900 => 54,
    21901 => 54,
    21902 => 54,
    21903 => 54,
    21904 => 54,
    21905 => 54,
    21906 => 54,
    21907 => 54,
    21908 => 54,
    21909 => 54,
    21910 => 54,
    21911 => 54,
    21912 => 54,
    21913 => 54,
    21914 => 54,
    21915 => 54,
    21916 => 54,
    21917 => 54,
    21918 => 54,
    21919 => 54,
    21920 => 54,
    21921 => 54,
    21922 => 54,
    21923 => 54,
    21924 => 54,
    21925 => 54,
    21926 => 54,
    21927 => 54,
    21928 => 54,
    21929 => 54,
    21930 => 54,
    21931 => 54,
    21932 => 54,
    21933 => 54,
    21934 => 54,
    21935 => 54,
    21936 => 54,
    21937 => 54,
    21938 => 54,
    21939 => 54,
    21940 => 54,
    21941 => 54,
    21942 => 54,
    21943 => 54,
    21944 => 54,
    21945 => 54,
    21946 => 54,
    21947 => 54,
    21948 => 54,
    21949 => 54,
    21950 => 54,
    21951 => 54,
    21952 => 54,
    21953 => 54,
    21954 => 54,
    21955 => 54,
    21956 => 54,
    21957 => 54,
    21958 => 54,
    21959 => 54,
    21960 => 54,
    21961 => 54,
    21962 => 54,
    21963 => 54,
    21964 => 54,
    21965 => 54,
    21966 => 54,
    21967 => 54,
    21968 => 54,
    21969 => 54,
    21970 => 54,
    21971 => 54,
    21972 => 54,
    21973 => 54,
    21974 => 54,
    21975 => 54,
    21976 => 54,
    21977 => 54,
    21978 => 54,
    21979 => 54,
    21980 => 54,
    21981 => 54,
    21982 => 54,
    21983 => 54,
    21984 => 54,
    21985 => 54,
    21986 => 54,
    21987 => 54,
    21988 => 54,
    21989 => 54,
    21990 => 54,
    21991 => 54,
    21992 => 54,
    21993 => 54,
    21994 => 54,
    21995 => 54,
    21996 => 54,
    21997 => 54,
    21998 => 54,
    21999 => 54,
    22000 => 54,
    22001 => 54,
    22002 => 54,
    22003 => 54,
    22004 => 54,
    22005 => 54,
    22006 => 54,
    22007 => 54,
    22008 => 54,
    22009 => 54,
    22010 => 54,
    22011 => 54,
    22012 => 54,
    22013 => 54,
    22014 => 54,
    22015 => 54,
    22016 => 54,
    22017 => 54,
    22018 => 54,
    22019 => 54,
    22020 => 54,
    22021 => 54,
    22022 => 54,
    22023 => 54,
    22024 => 54,
    22025 => 54,
    22026 => 54,
    22027 => 54,
    22028 => 54,
    22029 => 54,
    22030 => 54,
    22031 => 54,
    22032 => 54,
    22033 => 54,
    22034 => 54,
    22035 => 54,
    22036 => 54,
    22037 => 54,
    22038 => 54,
    22039 => 54,
    22040 => 54,
    22041 => 54,
    22042 => 54,
    22043 => 54,
    22044 => 54,
    22045 => 54,
    22046 => 54,
    22047 => 54,
    22048 => 54,
    22049 => 54,
    22050 => 54,
    22051 => 54,
    22052 => 54,
    22053 => 54,
    22054 => 54,
    22055 => 54,
    22056 => 54,
    22057 => 54,
    22058 => 54,
    22059 => 54,
    22060 => 54,
    22061 => 54,
    22062 => 54,
    22063 => 54,
    22064 => 54,
    22065 => 54,
    22066 => 54,
    22067 => 54,
    22068 => 54,
    22069 => 54,
    22070 => 54,
    22071 => 54,
    22072 => 54,
    22073 => 54,
    22074 => 54,
    22075 => 54,
    22076 => 54,
    22077 => 54,
    22078 => 54,
    22079 => 54,
    22080 => 54,
    22081 => 54,
    22082 => 54,
    22083 => 54,
    22084 => 54,
    22085 => 54,
    22086 => 54,
    22087 => 54,
    22088 => 54,
    22089 => 54,
    22090 => 54,
    22091 => 54,
    22092 => 54,
    22093 => 54,
    22094 => 54,
    22095 => 54,
    22096 => 54,
    22097 => 54,
    22098 => 54,
    22099 => 54,
    22100 => 54,
    22101 => 54,
    22102 => 54,
    22103 => 54,
    22104 => 54,
    22105 => 54,
    22106 => 54,
    22107 => 54,
    22108 => 54,
    22109 => 54,
    22110 => 54,
    22111 => 54,
    22112 => 54,
    22113 => 54,
    22114 => 54,
    22115 => 54,
    22116 => 54,
    22117 => 54,
    22118 => 54,
    22119 => 54,
    22120 => 54,
    22121 => 54,
    22122 => 54,
    22123 => 54,
    22124 => 54,
    22125 => 54,
    22126 => 54,
    22127 => 54,
    22128 => 54,
    22129 => 54,
    22130 => 54,
    22131 => 54,
    22132 => 54,
    22133 => 54,
    22134 => 54,
    22135 => 54,
    22136 => 54,
    22137 => 54,
    22138 => 54,
    22139 => 54,
    22140 => 54,
    22141 => 54,
    22142 => 54,
    22143 => 54,
    22144 => 54,
    22145 => 54,
    22146 => 54,
    22147 => 54,
    22148 => 54,
    22149 => 54,
    22150 => 54,
    22151 => 54,
    22152 => 54,
    22153 => 54,
    22154 => 54,
    22155 => 54,
    22156 => 54,
    22157 => 54,
    22158 => 54,
    22159 => 54,
    22160 => 54,
    22161 => 54,
    22162 => 54,
    22163 => 54,
    22164 => 54,
    22165 => 54,
    22166 => 54,
    22167 => 54,
    22168 => 54,
    22169 => 54,
    22170 => 54,
    22171 => 54,
    22172 => 54,
    22173 => 54,
    22174 => 54,
    22175 => 54,
    22176 => 54,
    22177 => 54,
    22178 => 54,
    22179 => 54,
    22180 => 54,
    22181 => 54,
    22182 => 54,
    22183 => 54,
    22184 => 54,
    22185 => 54,
    22186 => 54,
    22187 => 53,
    22188 => 53,
    22189 => 53,
    22190 => 53,
    22191 => 53,
    22192 => 53,
    22193 => 53,
    22194 => 53,
    22195 => 53,
    22196 => 53,
    22197 => 53,
    22198 => 53,
    22199 => 53,
    22200 => 53,
    22201 => 53,
    22202 => 53,
    22203 => 53,
    22204 => 53,
    22205 => 53,
    22206 => 53,
    22207 => 53,
    22208 => 53,
    22209 => 53,
    22210 => 53,
    22211 => 53,
    22212 => 53,
    22213 => 53,
    22214 => 53,
    22215 => 53,
    22216 => 53,
    22217 => 53,
    22218 => 53,
    22219 => 53,
    22220 => 53,
    22221 => 53,
    22222 => 53,
    22223 => 53,
    22224 => 53,
    22225 => 53,
    22226 => 53,
    22227 => 53,
    22228 => 53,
    22229 => 53,
    22230 => 53,
    22231 => 53,
    22232 => 53,
    22233 => 53,
    22234 => 53,
    22235 => 53,
    22236 => 53,
    22237 => 53,
    22238 => 53,
    22239 => 53,
    22240 => 53,
    22241 => 53,
    22242 => 53,
    22243 => 53,
    22244 => 53,
    22245 => 53,
    22246 => 53,
    22247 => 53,
    22248 => 53,
    22249 => 53,
    22250 => 53,
    22251 => 53,
    22252 => 53,
    22253 => 53,
    22254 => 53,
    22255 => 53,
    22256 => 53,
    22257 => 53,
    22258 => 53,
    22259 => 53,
    22260 => 53,
    22261 => 53,
    22262 => 53,
    22263 => 53,
    22264 => 53,
    22265 => 53,
    22266 => 53,
    22267 => 53,
    22268 => 53,
    22269 => 53,
    22270 => 53,
    22271 => 53,
    22272 => 53,
    22273 => 53,
    22274 => 53,
    22275 => 53,
    22276 => 53,
    22277 => 53,
    22278 => 53,
    22279 => 53,
    22280 => 53,
    22281 => 53,
    22282 => 53,
    22283 => 53,
    22284 => 53,
    22285 => 53,
    22286 => 53,
    22287 => 53,
    22288 => 53,
    22289 => 53,
    22290 => 53,
    22291 => 53,
    22292 => 53,
    22293 => 53,
    22294 => 53,
    22295 => 53,
    22296 => 53,
    22297 => 53,
    22298 => 53,
    22299 => 53,
    22300 => 53,
    22301 => 53,
    22302 => 53,
    22303 => 53,
    22304 => 53,
    22305 => 53,
    22306 => 53,
    22307 => 53,
    22308 => 53,
    22309 => 53,
    22310 => 53,
    22311 => 53,
    22312 => 53,
    22313 => 53,
    22314 => 53,
    22315 => 53,
    22316 => 53,
    22317 => 53,
    22318 => 53,
    22319 => 53,
    22320 => 53,
    22321 => 53,
    22322 => 53,
    22323 => 53,
    22324 => 53,
    22325 => 53,
    22326 => 53,
    22327 => 53,
    22328 => 53,
    22329 => 53,
    22330 => 53,
    22331 => 53,
    22332 => 53,
    22333 => 53,
    22334 => 53,
    22335 => 53,
    22336 => 53,
    22337 => 53,
    22338 => 53,
    22339 => 53,
    22340 => 53,
    22341 => 53,
    22342 => 53,
    22343 => 53,
    22344 => 53,
    22345 => 53,
    22346 => 53,
    22347 => 53,
    22348 => 53,
    22349 => 53,
    22350 => 53,
    22351 => 53,
    22352 => 53,
    22353 => 53,
    22354 => 53,
    22355 => 53,
    22356 => 53,
    22357 => 53,
    22358 => 53,
    22359 => 53,
    22360 => 53,
    22361 => 53,
    22362 => 53,
    22363 => 53,
    22364 => 53,
    22365 => 53,
    22366 => 53,
    22367 => 53,
    22368 => 53,
    22369 => 53,
    22370 => 53,
    22371 => 53,
    22372 => 53,
    22373 => 53,
    22374 => 53,
    22375 => 53,
    22376 => 53,
    22377 => 53,
    22378 => 53,
    22379 => 53,
    22380 => 53,
    22381 => 53,
    22382 => 53,
    22383 => 53,
    22384 => 53,
    22385 => 53,
    22386 => 53,
    22387 => 53,
    22388 => 53,
    22389 => 53,
    22390 => 53,
    22391 => 53,
    22392 => 53,
    22393 => 53,
    22394 => 53,
    22395 => 53,
    22396 => 53,
    22397 => 53,
    22398 => 53,
    22399 => 53,
    22400 => 53,
    22401 => 53,
    22402 => 53,
    22403 => 53,
    22404 => 53,
    22405 => 53,
    22406 => 53,
    22407 => 53,
    22408 => 53,
    22409 => 53,
    22410 => 53,
    22411 => 53,
    22412 => 53,
    22413 => 53,
    22414 => 53,
    22415 => 53,
    22416 => 53,
    22417 => 53,
    22418 => 53,
    22419 => 53,
    22420 => 53,
    22421 => 53,
    22422 => 53,
    22423 => 53,
    22424 => 53,
    22425 => 53,
    22426 => 53,
    22427 => 53,
    22428 => 53,
    22429 => 53,
    22430 => 53,
    22431 => 53,
    22432 => 53,
    22433 => 53,
    22434 => 53,
    22435 => 53,
    22436 => 53,
    22437 => 53,
    22438 => 53,
    22439 => 53,
    22440 => 53,
    22441 => 53,
    22442 => 53,
    22443 => 53,
    22444 => 53,
    22445 => 53,
    22446 => 53,
    22447 => 53,
    22448 => 53,
    22449 => 53,
    22450 => 53,
    22451 => 53,
    22452 => 53,
    22453 => 53,
    22454 => 53,
    22455 => 53,
    22456 => 53,
    22457 => 53,
    22458 => 53,
    22459 => 53,
    22460 => 53,
    22461 => 53,
    22462 => 53,
    22463 => 53,
    22464 => 53,
    22465 => 53,
    22466 => 53,
    22467 => 53,
    22468 => 53,
    22469 => 53,
    22470 => 53,
    22471 => 53,
    22472 => 53,
    22473 => 53,
    22474 => 53,
    22475 => 53,
    22476 => 53,
    22477 => 53,
    22478 => 53,
    22479 => 53,
    22480 => 53,
    22481 => 53,
    22482 => 53,
    22483 => 53,
    22484 => 53,
    22485 => 53,
    22486 => 53,
    22487 => 53,
    22488 => 53,
    22489 => 53,
    22490 => 53,
    22491 => 53,
    22492 => 53,
    22493 => 52,
    22494 => 52,
    22495 => 52,
    22496 => 52,
    22497 => 52,
    22498 => 52,
    22499 => 52,
    22500 => 52,
    22501 => 52,
    22502 => 52,
    22503 => 52,
    22504 => 52,
    22505 => 52,
    22506 => 52,
    22507 => 52,
    22508 => 52,
    22509 => 52,
    22510 => 52,
    22511 => 52,
    22512 => 52,
    22513 => 52,
    22514 => 52,
    22515 => 52,
    22516 => 52,
    22517 => 52,
    22518 => 52,
    22519 => 52,
    22520 => 52,
    22521 => 52,
    22522 => 52,
    22523 => 52,
    22524 => 52,
    22525 => 52,
    22526 => 52,
    22527 => 52,
    22528 => 52,
    22529 => 52,
    22530 => 52,
    22531 => 52,
    22532 => 52,
    22533 => 52,
    22534 => 52,
    22535 => 52,
    22536 => 52,
    22537 => 52,
    22538 => 52,
    22539 => 52,
    22540 => 52,
    22541 => 52,
    22542 => 52,
    22543 => 52,
    22544 => 52,
    22545 => 52,
    22546 => 52,
    22547 => 52,
    22548 => 52,
    22549 => 52,
    22550 => 52,
    22551 => 52,
    22552 => 52,
    22553 => 52,
    22554 => 52,
    22555 => 52,
    22556 => 52,
    22557 => 52,
    22558 => 52,
    22559 => 52,
    22560 => 52,
    22561 => 52,
    22562 => 52,
    22563 => 52,
    22564 => 52,
    22565 => 52,
    22566 => 52,
    22567 => 52,
    22568 => 52,
    22569 => 52,
    22570 => 52,
    22571 => 52,
    22572 => 52,
    22573 => 52,
    22574 => 52,
    22575 => 52,
    22576 => 52,
    22577 => 52,
    22578 => 52,
    22579 => 52,
    22580 => 52,
    22581 => 52,
    22582 => 52,
    22583 => 52,
    22584 => 52,
    22585 => 52,
    22586 => 52,
    22587 => 52,
    22588 => 52,
    22589 => 52,
    22590 => 52,
    22591 => 52,
    22592 => 52,
    22593 => 52,
    22594 => 52,
    22595 => 52,
    22596 => 52,
    22597 => 52,
    22598 => 52,
    22599 => 52,
    22600 => 52,
    22601 => 52,
    22602 => 52,
    22603 => 52,
    22604 => 52,
    22605 => 52,
    22606 => 52,
    22607 => 52,
    22608 => 52,
    22609 => 52,
    22610 => 52,
    22611 => 52,
    22612 => 52,
    22613 => 52,
    22614 => 52,
    22615 => 52,
    22616 => 52,
    22617 => 52,
    22618 => 52,
    22619 => 52,
    22620 => 52,
    22621 => 52,
    22622 => 52,
    22623 => 52,
    22624 => 52,
    22625 => 52,
    22626 => 52,
    22627 => 52,
    22628 => 52,
    22629 => 52,
    22630 => 52,
    22631 => 52,
    22632 => 52,
    22633 => 52,
    22634 => 52,
    22635 => 52,
    22636 => 52,
    22637 => 52,
    22638 => 52,
    22639 => 52,
    22640 => 52,
    22641 => 52,
    22642 => 52,
    22643 => 52,
    22644 => 52,
    22645 => 52,
    22646 => 52,
    22647 => 52,
    22648 => 52,
    22649 => 52,
    22650 => 52,
    22651 => 52,
    22652 => 52,
    22653 => 52,
    22654 => 52,
    22655 => 52,
    22656 => 52,
    22657 => 52,
    22658 => 52,
    22659 => 52,
    22660 => 52,
    22661 => 52,
    22662 => 52,
    22663 => 52,
    22664 => 52,
    22665 => 52,
    22666 => 52,
    22667 => 52,
    22668 => 52,
    22669 => 52,
    22670 => 52,
    22671 => 52,
    22672 => 52,
    22673 => 52,
    22674 => 52,
    22675 => 52,
    22676 => 52,
    22677 => 52,
    22678 => 52,
    22679 => 52,
    22680 => 52,
    22681 => 52,
    22682 => 52,
    22683 => 52,
    22684 => 52,
    22685 => 52,
    22686 => 52,
    22687 => 52,
    22688 => 52,
    22689 => 52,
    22690 => 52,
    22691 => 52,
    22692 => 52,
    22693 => 52,
    22694 => 52,
    22695 => 52,
    22696 => 52,
    22697 => 52,
    22698 => 52,
    22699 => 52,
    22700 => 52,
    22701 => 52,
    22702 => 52,
    22703 => 52,
    22704 => 52,
    22705 => 52,
    22706 => 52,
    22707 => 52,
    22708 => 52,
    22709 => 52,
    22710 => 52,
    22711 => 52,
    22712 => 52,
    22713 => 52,
    22714 => 52,
    22715 => 52,
    22716 => 52,
    22717 => 52,
    22718 => 52,
    22719 => 52,
    22720 => 52,
    22721 => 52,
    22722 => 52,
    22723 => 52,
    22724 => 52,
    22725 => 52,
    22726 => 52,
    22727 => 52,
    22728 => 52,
    22729 => 52,
    22730 => 52,
    22731 => 52,
    22732 => 52,
    22733 => 52,
    22734 => 52,
    22735 => 52,
    22736 => 52,
    22737 => 52,
    22738 => 52,
    22739 => 52,
    22740 => 52,
    22741 => 52,
    22742 => 52,
    22743 => 52,
    22744 => 52,
    22745 => 52,
    22746 => 52,
    22747 => 52,
    22748 => 52,
    22749 => 52,
    22750 => 52,
    22751 => 52,
    22752 => 52,
    22753 => 52,
    22754 => 52,
    22755 => 52,
    22756 => 52,
    22757 => 52,
    22758 => 52,
    22759 => 52,
    22760 => 52,
    22761 => 52,
    22762 => 52,
    22763 => 52,
    22764 => 52,
    22765 => 52,
    22766 => 52,
    22767 => 52,
    22768 => 52,
    22769 => 52,
    22770 => 52,
    22771 => 52,
    22772 => 52,
    22773 => 52,
    22774 => 52,
    22775 => 52,
    22776 => 52,
    22777 => 52,
    22778 => 52,
    22779 => 52,
    22780 => 52,
    22781 => 52,
    22782 => 52,
    22783 => 52,
    22784 => 52,
    22785 => 52,
    22786 => 52,
    22787 => 51,
    22788 => 51,
    22789 => 51,
    22790 => 51,
    22791 => 51,
    22792 => 51,
    22793 => 51,
    22794 => 51,
    22795 => 51,
    22796 => 51,
    22797 => 51,
    22798 => 51,
    22799 => 51,
    22800 => 51,
    22801 => 51,
    22802 => 51,
    22803 => 51,
    22804 => 51,
    22805 => 51,
    22806 => 51,
    22807 => 51,
    22808 => 51,
    22809 => 51,
    22810 => 51,
    22811 => 51,
    22812 => 51,
    22813 => 51,
    22814 => 51,
    22815 => 51,
    22816 => 51,
    22817 => 51,
    22818 => 51,
    22819 => 51,
    22820 => 51,
    22821 => 51,
    22822 => 51,
    22823 => 51,
    22824 => 51,
    22825 => 51,
    22826 => 51,
    22827 => 51,
    22828 => 51,
    22829 => 51,
    22830 => 51,
    22831 => 51,
    22832 => 51,
    22833 => 51,
    22834 => 51,
    22835 => 51,
    22836 => 51,
    22837 => 51,
    22838 => 51,
    22839 => 51,
    22840 => 51,
    22841 => 51,
    22842 => 51,
    22843 => 51,
    22844 => 51,
    22845 => 51,
    22846 => 51,
    22847 => 51,
    22848 => 51,
    22849 => 51,
    22850 => 51,
    22851 => 51,
    22852 => 51,
    22853 => 51,
    22854 => 51,
    22855 => 51,
    22856 => 51,
    22857 => 51,
    22858 => 51,
    22859 => 51,
    22860 => 51,
    22861 => 51,
    22862 => 51,
    22863 => 51,
    22864 => 51,
    22865 => 51,
    22866 => 51,
    22867 => 51,
    22868 => 51,
    22869 => 51,
    22870 => 51,
    22871 => 51,
    22872 => 51,
    22873 => 51,
    22874 => 51,
    22875 => 51,
    22876 => 51,
    22877 => 51,
    22878 => 51,
    22879 => 51,
    22880 => 51,
    22881 => 51,
    22882 => 51,
    22883 => 51,
    22884 => 51,
    22885 => 51,
    22886 => 51,
    22887 => 51,
    22888 => 51,
    22889 => 51,
    22890 => 51,
    22891 => 51,
    22892 => 51,
    22893 => 51,
    22894 => 51,
    22895 => 51,
    22896 => 51,
    22897 => 51,
    22898 => 51,
    22899 => 51,
    22900 => 51,
    22901 => 51,
    22902 => 51,
    22903 => 51,
    22904 => 51,
    22905 => 51,
    22906 => 51,
    22907 => 51,
    22908 => 51,
    22909 => 51,
    22910 => 51,
    22911 => 51,
    22912 => 51,
    22913 => 51,
    22914 => 51,
    22915 => 51,
    22916 => 51,
    22917 => 51,
    22918 => 51,
    22919 => 51,
    22920 => 51,
    22921 => 51,
    22922 => 51,
    22923 => 51,
    22924 => 51,
    22925 => 51,
    22926 => 51,
    22927 => 51,
    22928 => 51,
    22929 => 51,
    22930 => 51,
    22931 => 51,
    22932 => 51,
    22933 => 51,
    22934 => 51,
    22935 => 51,
    22936 => 51,
    22937 => 51,
    22938 => 51,
    22939 => 51,
    22940 => 51,
    22941 => 51,
    22942 => 51,
    22943 => 51,
    22944 => 51,
    22945 => 51,
    22946 => 51,
    22947 => 51,
    22948 => 51,
    22949 => 51,
    22950 => 51,
    22951 => 51,
    22952 => 51,
    22953 => 51,
    22954 => 51,
    22955 => 51,
    22956 => 51,
    22957 => 51,
    22958 => 51,
    22959 => 51,
    22960 => 51,
    22961 => 51,
    22962 => 51,
    22963 => 51,
    22964 => 51,
    22965 => 51,
    22966 => 51,
    22967 => 51,
    22968 => 51,
    22969 => 51,
    22970 => 51,
    22971 => 51,
    22972 => 51,
    22973 => 51,
    22974 => 51,
    22975 => 51,
    22976 => 51,
    22977 => 51,
    22978 => 51,
    22979 => 51,
    22980 => 51,
    22981 => 51,
    22982 => 51,
    22983 => 51,
    22984 => 51,
    22985 => 51,
    22986 => 51,
    22987 => 51,
    22988 => 51,
    22989 => 51,
    22990 => 51,
    22991 => 51,
    22992 => 51,
    22993 => 51,
    22994 => 51,
    22995 => 51,
    22996 => 51,
    22997 => 51,
    22998 => 51,
    22999 => 51,
    23000 => 51,
    23001 => 51,
    23002 => 51,
    23003 => 51,
    23004 => 51,
    23005 => 51,
    23006 => 51,
    23007 => 51,
    23008 => 51,
    23009 => 51,
    23010 => 51,
    23011 => 51,
    23012 => 51,
    23013 => 51,
    23014 => 51,
    23015 => 51,
    23016 => 51,
    23017 => 51,
    23018 => 51,
    23019 => 51,
    23020 => 51,
    23021 => 51,
    23022 => 51,
    23023 => 51,
    23024 => 51,
    23025 => 51,
    23026 => 51,
    23027 => 51,
    23028 => 51,
    23029 => 51,
    23030 => 51,
    23031 => 51,
    23032 => 51,
    23033 => 51,
    23034 => 51,
    23035 => 51,
    23036 => 51,
    23037 => 51,
    23038 => 51,
    23039 => 51,
    23040 => 51,
    23041 => 51,
    23042 => 51,
    23043 => 51,
    23044 => 51,
    23045 => 51,
    23046 => 51,
    23047 => 51,
    23048 => 51,
    23049 => 51,
    23050 => 51,
    23051 => 51,
    23052 => 51,
    23053 => 51,
    23054 => 51,
    23055 => 51,
    23056 => 51,
    23057 => 51,
    23058 => 51,
    23059 => 51,
    23060 => 51,
    23061 => 51,
    23062 => 51,
    23063 => 51,
    23064 => 51,
    23065 => 51,
    23066 => 51,
    23067 => 51,
    23068 => 51,
    23069 => 50,
    23070 => 50,
    23071 => 50,
    23072 => 50,
    23073 => 50,
    23074 => 50,
    23075 => 50,
    23076 => 50,
    23077 => 50,
    23078 => 50,
    23079 => 50,
    23080 => 50,
    23081 => 50,
    23082 => 50,
    23083 => 50,
    23084 => 50,
    23085 => 50,
    23086 => 50,
    23087 => 50,
    23088 => 50,
    23089 => 50,
    23090 => 50,
    23091 => 50,
    23092 => 50,
    23093 => 50,
    23094 => 50,
    23095 => 50,
    23096 => 50,
    23097 => 50,
    23098 => 50,
    23099 => 50,
    23100 => 50,
    23101 => 50,
    23102 => 50,
    23103 => 50,
    23104 => 50,
    23105 => 50,
    23106 => 50,
    23107 => 50,
    23108 => 50,
    23109 => 50,
    23110 => 50,
    23111 => 50,
    23112 => 50,
    23113 => 50,
    23114 => 50,
    23115 => 50,
    23116 => 50,
    23117 => 50,
    23118 => 50,
    23119 => 50,
    23120 => 50,
    23121 => 50,
    23122 => 50,
    23123 => 50,
    23124 => 50,
    23125 => 50,
    23126 => 50,
    23127 => 50,
    23128 => 50,
    23129 => 50,
    23130 => 50,
    23131 => 50,
    23132 => 50,
    23133 => 50,
    23134 => 50,
    23135 => 50,
    23136 => 50,
    23137 => 50,
    23138 => 50,
    23139 => 50,
    23140 => 50,
    23141 => 50,
    23142 => 50,
    23143 => 50,
    23144 => 50,
    23145 => 50,
    23146 => 50,
    23147 => 50,
    23148 => 50,
    23149 => 50,
    23150 => 50,
    23151 => 50,
    23152 => 50,
    23153 => 50,
    23154 => 50,
    23155 => 50,
    23156 => 50,
    23157 => 50,
    23158 => 50,
    23159 => 50,
    23160 => 50,
    23161 => 50,
    23162 => 50,
    23163 => 50,
    23164 => 50,
    23165 => 50,
    23166 => 50,
    23167 => 50,
    23168 => 50,
    23169 => 50,
    23170 => 50,
    23171 => 50,
    23172 => 50,
    23173 => 50,
    23174 => 50,
    23175 => 50,
    23176 => 50,
    23177 => 50,
    23178 => 50,
    23179 => 50,
    23180 => 50,
    23181 => 50,
    23182 => 50,
    23183 => 50,
    23184 => 50,
    23185 => 50,
    23186 => 50,
    23187 => 50,
    23188 => 50,
    23189 => 50,
    23190 => 50,
    23191 => 50,
    23192 => 50,
    23193 => 50,
    23194 => 50,
    23195 => 50,
    23196 => 50,
    23197 => 50,
    23198 => 50,
    23199 => 50,
    23200 => 50,
    23201 => 50,
    23202 => 50,
    23203 => 50,
    23204 => 50,
    23205 => 50,
    23206 => 50,
    23207 => 50,
    23208 => 50,
    23209 => 50,
    23210 => 50,
    23211 => 50,
    23212 => 50,
    23213 => 50,
    23214 => 50,
    23215 => 50,
    23216 => 50,
    23217 => 50,
    23218 => 50,
    23219 => 50,
    23220 => 50,
    23221 => 50,
    23222 => 50,
    23223 => 50,
    23224 => 50,
    23225 => 50,
    23226 => 50,
    23227 => 50,
    23228 => 50,
    23229 => 50,
    23230 => 50,
    23231 => 50,
    23232 => 50,
    23233 => 50,
    23234 => 50,
    23235 => 50,
    23236 => 50,
    23237 => 50,
    23238 => 50,
    23239 => 50,
    23240 => 50,
    23241 => 50,
    23242 => 50,
    23243 => 50,
    23244 => 50,
    23245 => 50,
    23246 => 50,
    23247 => 50,
    23248 => 50,
    23249 => 50,
    23250 => 50,
    23251 => 50,
    23252 => 50,
    23253 => 50,
    23254 => 50,
    23255 => 50,
    23256 => 50,
    23257 => 50,
    23258 => 50,
    23259 => 50,
    23260 => 50,
    23261 => 50,
    23262 => 50,
    23263 => 50,
    23264 => 50,
    23265 => 50,
    23266 => 50,
    23267 => 50,
    23268 => 50,
    23269 => 50,
    23270 => 50,
    23271 => 50,
    23272 => 50,
    23273 => 50,
    23274 => 50,
    23275 => 50,
    23276 => 50,
    23277 => 50,
    23278 => 50,
    23279 => 50,
    23280 => 50,
    23281 => 50,
    23282 => 50,
    23283 => 50,
    23284 => 50,
    23285 => 50,
    23286 => 50,
    23287 => 50,
    23288 => 50,
    23289 => 50,
    23290 => 50,
    23291 => 50,
    23292 => 50,
    23293 => 50,
    23294 => 50,
    23295 => 50,
    23296 => 50,
    23297 => 50,
    23298 => 50,
    23299 => 50,
    23300 => 50,
    23301 => 50,
    23302 => 50,
    23303 => 50,
    23304 => 50,
    23305 => 50,
    23306 => 50,
    23307 => 50,
    23308 => 50,
    23309 => 50,
    23310 => 50,
    23311 => 50,
    23312 => 50,
    23313 => 50,
    23314 => 50,
    23315 => 50,
    23316 => 50,
    23317 => 50,
    23318 => 50,
    23319 => 50,
    23320 => 50,
    23321 => 50,
    23322 => 50,
    23323 => 50,
    23324 => 50,
    23325 => 50,
    23326 => 50,
    23327 => 50,
    23328 => 50,
    23329 => 50,
    23330 => 50,
    23331 => 50,
    23332 => 50,
    23333 => 50,
    23334 => 50,
    23335 => 50,
    23336 => 50,
    23337 => 50,
    23338 => 50,
    23339 => 50,
    23340 => 50,
    23341 => 49,
    23342 => 49,
    23343 => 49,
    23344 => 49,
    23345 => 49,
    23346 => 49,
    23347 => 49,
    23348 => 49,
    23349 => 49,
    23350 => 49,
    23351 => 49,
    23352 => 49,
    23353 => 49,
    23354 => 49,
    23355 => 49,
    23356 => 49,
    23357 => 49,
    23358 => 49,
    23359 => 49,
    23360 => 49,
    23361 => 49,
    23362 => 49,
    23363 => 49,
    23364 => 49,
    23365 => 49,
    23366 => 49,
    23367 => 49,
    23368 => 49,
    23369 => 49,
    23370 => 49,
    23371 => 49,
    23372 => 49,
    23373 => 49,
    23374 => 49,
    23375 => 49,
    23376 => 49,
    23377 => 49,
    23378 => 49,
    23379 => 49,
    23380 => 49,
    23381 => 49,
    23382 => 49,
    23383 => 49,
    23384 => 49,
    23385 => 49,
    23386 => 49,
    23387 => 49,
    23388 => 49,
    23389 => 49,
    23390 => 49,
    23391 => 49,
    23392 => 49,
    23393 => 49,
    23394 => 49,
    23395 => 49,
    23396 => 49,
    23397 => 49,
    23398 => 49,
    23399 => 49,
    23400 => 49,
    23401 => 49,
    23402 => 49,
    23403 => 49,
    23404 => 49,
    23405 => 49,
    23406 => 49,
    23407 => 49,
    23408 => 49,
    23409 => 49,
    23410 => 49,
    23411 => 49,
    23412 => 49,
    23413 => 49,
    23414 => 49,
    23415 => 49,
    23416 => 49,
    23417 => 49,
    23418 => 49,
    23419 => 49,
    23420 => 49,
    23421 => 49,
    23422 => 49,
    23423 => 49,
    23424 => 49,
    23425 => 49,
    23426 => 49,
    23427 => 49,
    23428 => 49,
    23429 => 49,
    23430 => 49,
    23431 => 49,
    23432 => 49,
    23433 => 49,
    23434 => 49,
    23435 => 49,
    23436 => 49,
    23437 => 49,
    23438 => 49,
    23439 => 49,
    23440 => 49,
    23441 => 49,
    23442 => 49,
    23443 => 49,
    23444 => 49,
    23445 => 49,
    23446 => 49,
    23447 => 49,
    23448 => 49,
    23449 => 49,
    23450 => 49,
    23451 => 49,
    23452 => 49,
    23453 => 49,
    23454 => 49,
    23455 => 49,
    23456 => 49,
    23457 => 49,
    23458 => 49,
    23459 => 49,
    23460 => 49,
    23461 => 49,
    23462 => 49,
    23463 => 49,
    23464 => 49,
    23465 => 49,
    23466 => 49,
    23467 => 49,
    23468 => 49,
    23469 => 49,
    23470 => 49,
    23471 => 49,
    23472 => 49,
    23473 => 49,
    23474 => 49,
    23475 => 49,
    23476 => 49,
    23477 => 49,
    23478 => 49,
    23479 => 49,
    23480 => 49,
    23481 => 49,
    23482 => 49,
    23483 => 49,
    23484 => 49,
    23485 => 49,
    23486 => 49,
    23487 => 49,
    23488 => 49,
    23489 => 49,
    23490 => 49,
    23491 => 49,
    23492 => 49,
    23493 => 49,
    23494 => 49,
    23495 => 49,
    23496 => 49,
    23497 => 49,
    23498 => 49,
    23499 => 49,
    23500 => 49,
    23501 => 49,
    23502 => 49,
    23503 => 49,
    23504 => 49,
    23505 => 49,
    23506 => 49,
    23507 => 49,
    23508 => 49,
    23509 => 49,
    23510 => 49,
    23511 => 49,
    23512 => 49,
    23513 => 49,
    23514 => 49,
    23515 => 49,
    23516 => 49,
    23517 => 49,
    23518 => 49,
    23519 => 49,
    23520 => 49,
    23521 => 49,
    23522 => 49,
    23523 => 49,
    23524 => 49,
    23525 => 49,
    23526 => 49,
    23527 => 49,
    23528 => 49,
    23529 => 49,
    23530 => 49,
    23531 => 49,
    23532 => 49,
    23533 => 49,
    23534 => 49,
    23535 => 49,
    23536 => 49,
    23537 => 49,
    23538 => 49,
    23539 => 49,
    23540 => 49,
    23541 => 49,
    23542 => 49,
    23543 => 49,
    23544 => 49,
    23545 => 49,
    23546 => 49,
    23547 => 49,
    23548 => 49,
    23549 => 49,
    23550 => 49,
    23551 => 49,
    23552 => 49,
    23553 => 49,
    23554 => 49,
    23555 => 49,
    23556 => 49,
    23557 => 49,
    23558 => 49,
    23559 => 49,
    23560 => 49,
    23561 => 49,
    23562 => 49,
    23563 => 49,
    23564 => 49,
    23565 => 49,
    23566 => 49,
    23567 => 49,
    23568 => 49,
    23569 => 49,
    23570 => 49,
    23571 => 49,
    23572 => 49,
    23573 => 49,
    23574 => 49,
    23575 => 49,
    23576 => 49,
    23577 => 49,
    23578 => 49,
    23579 => 49,
    23580 => 49,
    23581 => 49,
    23582 => 49,
    23583 => 49,
    23584 => 49,
    23585 => 49,
    23586 => 49,
    23587 => 49,
    23588 => 49,
    23589 => 49,
    23590 => 49,
    23591 => 49,
    23592 => 49,
    23593 => 49,
    23594 => 49,
    23595 => 49,
    23596 => 49,
    23597 => 49,
    23598 => 49,
    23599 => 49,
    23600 => 49,
    23601 => 49,
    23602 => 49,
    23603 => 49,
    23604 => 48,
    23605 => 48,
    23606 => 48,
    23607 => 48,
    23608 => 48,
    23609 => 48,
    23610 => 48,
    23611 => 48,
    23612 => 48,
    23613 => 48,
    23614 => 48,
    23615 => 48,
    23616 => 48,
    23617 => 48,
    23618 => 48,
    23619 => 48,
    23620 => 48,
    23621 => 48,
    23622 => 48,
    23623 => 48,
    23624 => 48,
    23625 => 48,
    23626 => 48,
    23627 => 48,
    23628 => 48,
    23629 => 48,
    23630 => 48,
    23631 => 48,
    23632 => 48,
    23633 => 48,
    23634 => 48,
    23635 => 48,
    23636 => 48,
    23637 => 48,
    23638 => 48,
    23639 => 48,
    23640 => 48,
    23641 => 48,
    23642 => 48,
    23643 => 48,
    23644 => 48,
    23645 => 48,
    23646 => 48,
    23647 => 48,
    23648 => 48,
    23649 => 48,
    23650 => 48,
    23651 => 48,
    23652 => 48,
    23653 => 48,
    23654 => 48,
    23655 => 48,
    23656 => 48,
    23657 => 48,
    23658 => 48,
    23659 => 48,
    23660 => 48,
    23661 => 48,
    23662 => 48,
    23663 => 48,
    23664 => 48,
    23665 => 48,
    23666 => 48,
    23667 => 48,
    23668 => 48,
    23669 => 48,
    23670 => 48,
    23671 => 48,
    23672 => 48,
    23673 => 48,
    23674 => 48,
    23675 => 48,
    23676 => 48,
    23677 => 48,
    23678 => 48,
    23679 => 48,
    23680 => 48,
    23681 => 48,
    23682 => 48,
    23683 => 48,
    23684 => 48,
    23685 => 48,
    23686 => 48,
    23687 => 48,
    23688 => 48,
    23689 => 48,
    23690 => 48,
    23691 => 48,
    23692 => 48,
    23693 => 48,
    23694 => 48,
    23695 => 48,
    23696 => 48,
    23697 => 48,
    23698 => 48,
    23699 => 48,
    23700 => 48,
    23701 => 48,
    23702 => 48,
    23703 => 48,
    23704 => 48,
    23705 => 48,
    23706 => 48,
    23707 => 48,
    23708 => 48,
    23709 => 48,
    23710 => 48,
    23711 => 48,
    23712 => 48,
    23713 => 48,
    23714 => 48,
    23715 => 48,
    23716 => 48,
    23717 => 48,
    23718 => 48,
    23719 => 48,
    23720 => 48,
    23721 => 48,
    23722 => 48,
    23723 => 48,
    23724 => 48,
    23725 => 48,
    23726 => 48,
    23727 => 48,
    23728 => 48,
    23729 => 48,
    23730 => 48,
    23731 => 48,
    23732 => 48,
    23733 => 48,
    23734 => 48,
    23735 => 48,
    23736 => 48,
    23737 => 48,
    23738 => 48,
    23739 => 48,
    23740 => 48,
    23741 => 48,
    23742 => 48,
    23743 => 48,
    23744 => 48,
    23745 => 48,
    23746 => 48,
    23747 => 48,
    23748 => 48,
    23749 => 48,
    23750 => 48,
    23751 => 48,
    23752 => 48,
    23753 => 48,
    23754 => 48,
    23755 => 48,
    23756 => 48,
    23757 => 48,
    23758 => 48,
    23759 => 48,
    23760 => 48,
    23761 => 48,
    23762 => 48,
    23763 => 48,
    23764 => 48,
    23765 => 48,
    23766 => 48,
    23767 => 48,
    23768 => 48,
    23769 => 48,
    23770 => 48,
    23771 => 48,
    23772 => 48,
    23773 => 48,
    23774 => 48,
    23775 => 48,
    23776 => 48,
    23777 => 48,
    23778 => 48,
    23779 => 48,
    23780 => 48,
    23781 => 48,
    23782 => 48,
    23783 => 48,
    23784 => 48,
    23785 => 48,
    23786 => 48,
    23787 => 48,
    23788 => 48,
    23789 => 48,
    23790 => 48,
    23791 => 48,
    23792 => 48,
    23793 => 48,
    23794 => 48,
    23795 => 48,
    23796 => 48,
    23797 => 48,
    23798 => 48,
    23799 => 48,
    23800 => 48,
    23801 => 48,
    23802 => 48,
    23803 => 48,
    23804 => 48,
    23805 => 48,
    23806 => 48,
    23807 => 48,
    23808 => 48,
    23809 => 48,
    23810 => 48,
    23811 => 48,
    23812 => 48,
    23813 => 48,
    23814 => 48,
    23815 => 48,
    23816 => 48,
    23817 => 48,
    23818 => 48,
    23819 => 48,
    23820 => 48,
    23821 => 48,
    23822 => 48,
    23823 => 48,
    23824 => 48,
    23825 => 48,
    23826 => 48,
    23827 => 48,
    23828 => 48,
    23829 => 48,
    23830 => 48,
    23831 => 48,
    23832 => 48,
    23833 => 48,
    23834 => 48,
    23835 => 48,
    23836 => 48,
    23837 => 48,
    23838 => 48,
    23839 => 48,
    23840 => 48,
    23841 => 48,
    23842 => 48,
    23843 => 48,
    23844 => 48,
    23845 => 48,
    23846 => 48,
    23847 => 48,
    23848 => 48,
    23849 => 48,
    23850 => 48,
    23851 => 48,
    23852 => 48,
    23853 => 48,
    23854 => 48,
    23855 => 48,
    23856 => 48,
    23857 => 48,
    23858 => 48,
    23859 => 48,
    23860 => 47,
    23861 => 47,
    23862 => 47,
    23863 => 47,
    23864 => 47,
    23865 => 47,
    23866 => 47,
    23867 => 47,
    23868 => 47,
    23869 => 47,
    23870 => 47,
    23871 => 47,
    23872 => 47,
    23873 => 47,
    23874 => 47,
    23875 => 47,
    23876 => 47,
    23877 => 47,
    23878 => 47,
    23879 => 47,
    23880 => 47,
    23881 => 47,
    23882 => 47,
    23883 => 47,
    23884 => 47,
    23885 => 47,
    23886 => 47,
    23887 => 47,
    23888 => 47,
    23889 => 47,
    23890 => 47,
    23891 => 47,
    23892 => 47,
    23893 => 47,
    23894 => 47,
    23895 => 47,
    23896 => 47,
    23897 => 47,
    23898 => 47,
    23899 => 47,
    23900 => 47,
    23901 => 47,
    23902 => 47,
    23903 => 47,
    23904 => 47,
    23905 => 47,
    23906 => 47,
    23907 => 47,
    23908 => 47,
    23909 => 47,
    23910 => 47,
    23911 => 47,
    23912 => 47,
    23913 => 47,
    23914 => 47,
    23915 => 47,
    23916 => 47,
    23917 => 47,
    23918 => 47,
    23919 => 47,
    23920 => 47,
    23921 => 47,
    23922 => 47,
    23923 => 47,
    23924 => 47,
    23925 => 47,
    23926 => 47,
    23927 => 47,
    23928 => 47,
    23929 => 47,
    23930 => 47,
    23931 => 47,
    23932 => 47,
    23933 => 47,
    23934 => 47,
    23935 => 47,
    23936 => 47,
    23937 => 47,
    23938 => 47,
    23939 => 47,
    23940 => 47,
    23941 => 47,
    23942 => 47,
    23943 => 47,
    23944 => 47,
    23945 => 47,
    23946 => 47,
    23947 => 47,
    23948 => 47,
    23949 => 47,
    23950 => 47,
    23951 => 47,
    23952 => 47,
    23953 => 47,
    23954 => 47,
    23955 => 47,
    23956 => 47,
    23957 => 47,
    23958 => 47,
    23959 => 47,
    23960 => 47,
    23961 => 47,
    23962 => 47,
    23963 => 47,
    23964 => 47,
    23965 => 47,
    23966 => 47,
    23967 => 47,
    23968 => 47,
    23969 => 47,
    23970 => 47,
    23971 => 47,
    23972 => 47,
    23973 => 47,
    23974 => 47,
    23975 => 47,
    23976 => 47,
    23977 => 47,
    23978 => 47,
    23979 => 47,
    23980 => 47,
    23981 => 47,
    23982 => 47,
    23983 => 47,
    23984 => 47,
    23985 => 47,
    23986 => 47,
    23987 => 47,
    23988 => 47,
    23989 => 47,
    23990 => 47,
    23991 => 47,
    23992 => 47,
    23993 => 47,
    23994 => 47,
    23995 => 47,
    23996 => 47,
    23997 => 47,
    23998 => 47,
    23999 => 47,
    24000 => 47,
    24001 => 47,
    24002 => 47,
    24003 => 47,
    24004 => 47,
    24005 => 47,
    24006 => 47,
    24007 => 47,
    24008 => 47,
    24009 => 47,
    24010 => 47,
    24011 => 47,
    24012 => 47,
    24013 => 47,
    24014 => 47,
    24015 => 47,
    24016 => 47,
    24017 => 47,
    24018 => 47,
    24019 => 47,
    24020 => 47,
    24021 => 47,
    24022 => 47,
    24023 => 47,
    24024 => 47,
    24025 => 47,
    24026 => 47,
    24027 => 47,
    24028 => 47,
    24029 => 47,
    24030 => 47,
    24031 => 47,
    24032 => 47,
    24033 => 47,
    24034 => 47,
    24035 => 47,
    24036 => 47,
    24037 => 47,
    24038 => 47,
    24039 => 47,
    24040 => 47,
    24041 => 47,
    24042 => 47,
    24043 => 47,
    24044 => 47,
    24045 => 47,
    24046 => 47,
    24047 => 47,
    24048 => 47,
    24049 => 47,
    24050 => 47,
    24051 => 47,
    24052 => 47,
    24053 => 47,
    24054 => 47,
    24055 => 47,
    24056 => 47,
    24057 => 47,
    24058 => 47,
    24059 => 47,
    24060 => 47,
    24061 => 47,
    24062 => 47,
    24063 => 47,
    24064 => 47,
    24065 => 47,
    24066 => 47,
    24067 => 47,
    24068 => 47,
    24069 => 47,
    24070 => 47,
    24071 => 47,
    24072 => 47,
    24073 => 47,
    24074 => 47,
    24075 => 47,
    24076 => 47,
    24077 => 47,
    24078 => 47,
    24079 => 47,
    24080 => 47,
    24081 => 47,
    24082 => 47,
    24083 => 47,
    24084 => 47,
    24085 => 47,
    24086 => 47,
    24087 => 47,
    24088 => 47,
    24089 => 47,
    24090 => 47,
    24091 => 47,
    24092 => 47,
    24093 => 47,
    24094 => 47,
    24095 => 47,
    24096 => 47,
    24097 => 47,
    24098 => 47,
    24099 => 47,
    24100 => 47,
    24101 => 47,
    24102 => 47,
    24103 => 47,
    24104 => 47,
    24105 => 47,
    24106 => 47,
    24107 => 47,
    24108 => 47,
    24109 => 46,
    24110 => 46,
    24111 => 46,
    24112 => 46,
    24113 => 46,
    24114 => 46,
    24115 => 46,
    24116 => 46,
    24117 => 46,
    24118 => 46,
    24119 => 46,
    24120 => 46,
    24121 => 46,
    24122 => 46,
    24123 => 46,
    24124 => 46,
    24125 => 46,
    24126 => 46,
    24127 => 46,
    24128 => 46,
    24129 => 46,
    24130 => 46,
    24131 => 46,
    24132 => 46,
    24133 => 46,
    24134 => 46,
    24135 => 46,
    24136 => 46,
    24137 => 46,
    24138 => 46,
    24139 => 46,
    24140 => 46,
    24141 => 46,
    24142 => 46,
    24143 => 46,
    24144 => 46,
    24145 => 46,
    24146 => 46,
    24147 => 46,
    24148 => 46,
    24149 => 46,
    24150 => 46,
    24151 => 46,
    24152 => 46,
    24153 => 46,
    24154 => 46,
    24155 => 46,
    24156 => 46,
    24157 => 46,
    24158 => 46,
    24159 => 46,
    24160 => 46,
    24161 => 46,
    24162 => 46,
    24163 => 46,
    24164 => 46,
    24165 => 46,
    24166 => 46,
    24167 => 46,
    24168 => 46,
    24169 => 46,
    24170 => 46,
    24171 => 46,
    24172 => 46,
    24173 => 46,
    24174 => 46,
    24175 => 46,
    24176 => 46,
    24177 => 46,
    24178 => 46,
    24179 => 46,
    24180 => 46,
    24181 => 46,
    24182 => 46,
    24183 => 46,
    24184 => 46,
    24185 => 46,
    24186 => 46,
    24187 => 46,
    24188 => 46,
    24189 => 46,
    24190 => 46,
    24191 => 46,
    24192 => 46,
    24193 => 46,
    24194 => 46,
    24195 => 46,
    24196 => 46,
    24197 => 46,
    24198 => 46,
    24199 => 46,
    24200 => 46,
    24201 => 46,
    24202 => 46,
    24203 => 46,
    24204 => 46,
    24205 => 46,
    24206 => 46,
    24207 => 46,
    24208 => 46,
    24209 => 46,
    24210 => 46,
    24211 => 46,
    24212 => 46,
    24213 => 46,
    24214 => 46,
    24215 => 46,
    24216 => 46,
    24217 => 46,
    24218 => 46,
    24219 => 46,
    24220 => 46,
    24221 => 46,
    24222 => 46,
    24223 => 46,
    24224 => 46,
    24225 => 46,
    24226 => 46,
    24227 => 46,
    24228 => 46,
    24229 => 46,
    24230 => 46,
    24231 => 46,
    24232 => 46,
    24233 => 46,
    24234 => 46,
    24235 => 46,
    24236 => 46,
    24237 => 46,
    24238 => 46,
    24239 => 46,
    24240 => 46,
    24241 => 46,
    24242 => 46,
    24243 => 46,
    24244 => 46,
    24245 => 46,
    24246 => 46,
    24247 => 46,
    24248 => 46,
    24249 => 46,
    24250 => 46,
    24251 => 46,
    24252 => 46,
    24253 => 46,
    24254 => 46,
    24255 => 46,
    24256 => 46,
    24257 => 46,
    24258 => 46,
    24259 => 46,
    24260 => 46,
    24261 => 46,
    24262 => 46,
    24263 => 46,
    24264 => 46,
    24265 => 46,
    24266 => 46,
    24267 => 46,
    24268 => 46,
    24269 => 46,
    24270 => 46,
    24271 => 46,
    24272 => 46,
    24273 => 46,
    24274 => 46,
    24275 => 46,
    24276 => 46,
    24277 => 46,
    24278 => 46,
    24279 => 46,
    24280 => 46,
    24281 => 46,
    24282 => 46,
    24283 => 46,
    24284 => 46,
    24285 => 46,
    24286 => 46,
    24287 => 46,
    24288 => 46,
    24289 => 46,
    24290 => 46,
    24291 => 46,
    24292 => 46,
    24293 => 46,
    24294 => 46,
    24295 => 46,
    24296 => 46,
    24297 => 46,
    24298 => 46,
    24299 => 46,
    24300 => 46,
    24301 => 46,
    24302 => 46,
    24303 => 46,
    24304 => 46,
    24305 => 46,
    24306 => 46,
    24307 => 46,
    24308 => 46,
    24309 => 46,
    24310 => 46,
    24311 => 46,
    24312 => 46,
    24313 => 46,
    24314 => 46,
    24315 => 46,
    24316 => 46,
    24317 => 46,
    24318 => 46,
    24319 => 46,
    24320 => 46,
    24321 => 46,
    24322 => 46,
    24323 => 46,
    24324 => 46,
    24325 => 46,
    24326 => 46,
    24327 => 46,
    24328 => 46,
    24329 => 46,
    24330 => 46,
    24331 => 46,
    24332 => 46,
    24333 => 46,
    24334 => 46,
    24335 => 46,
    24336 => 46,
    24337 => 46,
    24338 => 46,
    24339 => 46,
    24340 => 46,
    24341 => 46,
    24342 => 46,
    24343 => 46,
    24344 => 46,
    24345 => 46,
    24346 => 46,
    24347 => 46,
    24348 => 46,
    24349 => 46,
    24350 => 46,
    24351 => 45,
    24352 => 45,
    24353 => 45,
    24354 => 45,
    24355 => 45,
    24356 => 45,
    24357 => 45,
    24358 => 45,
    24359 => 45,
    24360 => 45,
    24361 => 45,
    24362 => 45,
    24363 => 45,
    24364 => 45,
    24365 => 45,
    24366 => 45,
    24367 => 45,
    24368 => 45,
    24369 => 45,
    24370 => 45,
    24371 => 45,
    24372 => 45,
    24373 => 45,
    24374 => 45,
    24375 => 45,
    24376 => 45,
    24377 => 45,
    24378 => 45,
    24379 => 45,
    24380 => 45,
    24381 => 45,
    24382 => 45,
    24383 => 45,
    24384 => 45,
    24385 => 45,
    24386 => 45,
    24387 => 45,
    24388 => 45,
    24389 => 45,
    24390 => 45,
    24391 => 45,
    24392 => 45,
    24393 => 45,
    24394 => 45,
    24395 => 45,
    24396 => 45,
    24397 => 45,
    24398 => 45,
    24399 => 45,
    24400 => 45,
    24401 => 45,
    24402 => 45,
    24403 => 45,
    24404 => 45,
    24405 => 45,
    24406 => 45,
    24407 => 45,
    24408 => 45,
    24409 => 45,
    24410 => 45,
    24411 => 45,
    24412 => 45,
    24413 => 45,
    24414 => 45,
    24415 => 45,
    24416 => 45,
    24417 => 45,
    24418 => 45,
    24419 => 45,
    24420 => 45,
    24421 => 45,
    24422 => 45,
    24423 => 45,
    24424 => 45,
    24425 => 45,
    24426 => 45,
    24427 => 45,
    24428 => 45,
    24429 => 45,
    24430 => 45,
    24431 => 45,
    24432 => 45,
    24433 => 45,
    24434 => 45,
    24435 => 45,
    24436 => 45,
    24437 => 45,
    24438 => 45,
    24439 => 45,
    24440 => 45,
    24441 => 45,
    24442 => 45,
    24443 => 45,
    24444 => 45,
    24445 => 45,
    24446 => 45,
    24447 => 45,
    24448 => 45,
    24449 => 45,
    24450 => 45,
    24451 => 45,
    24452 => 45,
    24453 => 45,
    24454 => 45,
    24455 => 45,
    24456 => 45,
    24457 => 45,
    24458 => 45,
    24459 => 45,
    24460 => 45,
    24461 => 45,
    24462 => 45,
    24463 => 45,
    24464 => 45,
    24465 => 45,
    24466 => 45,
    24467 => 45,
    24468 => 45,
    24469 => 45,
    24470 => 45,
    24471 => 45,
    24472 => 45,
    24473 => 45,
    24474 => 45,
    24475 => 45,
    24476 => 45,
    24477 => 45,
    24478 => 45,
    24479 => 45,
    24480 => 45,
    24481 => 45,
    24482 => 45,
    24483 => 45,
    24484 => 45,
    24485 => 45,
    24486 => 45,
    24487 => 45,
    24488 => 45,
    24489 => 45,
    24490 => 45,
    24491 => 45,
    24492 => 45,
    24493 => 45,
    24494 => 45,
    24495 => 45,
    24496 => 45,
    24497 => 45,
    24498 => 45,
    24499 => 45,
    24500 => 45,
    24501 => 45,
    24502 => 45,
    24503 => 45,
    24504 => 45,
    24505 => 45,
    24506 => 45,
    24507 => 45,
    24508 => 45,
    24509 => 45,
    24510 => 45,
    24511 => 45,
    24512 => 45,
    24513 => 45,
    24514 => 45,
    24515 => 45,
    24516 => 45,
    24517 => 45,
    24518 => 45,
    24519 => 45,
    24520 => 45,
    24521 => 45,
    24522 => 45,
    24523 => 45,
    24524 => 45,
    24525 => 45,
    24526 => 45,
    24527 => 45,
    24528 => 45,
    24529 => 45,
    24530 => 45,
    24531 => 45,
    24532 => 45,
    24533 => 45,
    24534 => 45,
    24535 => 45,
    24536 => 45,
    24537 => 45,
    24538 => 45,
    24539 => 45,
    24540 => 45,
    24541 => 45,
    24542 => 45,
    24543 => 45,
    24544 => 45,
    24545 => 45,
    24546 => 45,
    24547 => 45,
    24548 => 45,
    24549 => 45,
    24550 => 45,
    24551 => 45,
    24552 => 45,
    24553 => 45,
    24554 => 45,
    24555 => 45,
    24556 => 45,
    24557 => 45,
    24558 => 45,
    24559 => 45,
    24560 => 45,
    24561 => 45,
    24562 => 45,
    24563 => 45,
    24564 => 45,
    24565 => 45,
    24566 => 45,
    24567 => 45,
    24568 => 45,
    24569 => 45,
    24570 => 45,
    24571 => 45,
    24572 => 45,
    24573 => 45,
    24574 => 45,
    24575 => 45,
    24576 => 45,
    24577 => 45,
    24578 => 45,
    24579 => 45,
    24580 => 45,
    24581 => 45,
    24582 => 45,
    24583 => 45,
    24584 => 45,
    24585 => 45,
    24586 => 45,
    24587 => 45,
    24588 => 44,
    24589 => 44,
    24590 => 44,
    24591 => 44,
    24592 => 44,
    24593 => 44,
    24594 => 44,
    24595 => 44,
    24596 => 44,
    24597 => 44,
    24598 => 44,
    24599 => 44,
    24600 => 44,
    24601 => 44,
    24602 => 44,
    24603 => 44,
    24604 => 44,
    24605 => 44,
    24606 => 44,
    24607 => 44,
    24608 => 44,
    24609 => 44,
    24610 => 44,
    24611 => 44,
    24612 => 44,
    24613 => 44,
    24614 => 44,
    24615 => 44,
    24616 => 44,
    24617 => 44,
    24618 => 44,
    24619 => 44,
    24620 => 44,
    24621 => 44,
    24622 => 44,
    24623 => 44,
    24624 => 44,
    24625 => 44,
    24626 => 44,
    24627 => 44,
    24628 => 44,
    24629 => 44,
    24630 => 44,
    24631 => 44,
    24632 => 44,
    24633 => 44,
    24634 => 44,
    24635 => 44,
    24636 => 44,
    24637 => 44,
    24638 => 44,
    24639 => 44,
    24640 => 44,
    24641 => 44,
    24642 => 44,
    24643 => 44,
    24644 => 44,
    24645 => 44,
    24646 => 44,
    24647 => 44,
    24648 => 44,
    24649 => 44,
    24650 => 44,
    24651 => 44,
    24652 => 44,
    24653 => 44,
    24654 => 44,
    24655 => 44,
    24656 => 44,
    24657 => 44,
    24658 => 44,
    24659 => 44,
    24660 => 44,
    24661 => 44,
    24662 => 44,
    24663 => 44,
    24664 => 44,
    24665 => 44,
    24666 => 44,
    24667 => 44,
    24668 => 44,
    24669 => 44,
    24670 => 44,
    24671 => 44,
    24672 => 44,
    24673 => 44,
    24674 => 44,
    24675 => 44,
    24676 => 44,
    24677 => 44,
    24678 => 44,
    24679 => 44,
    24680 => 44,
    24681 => 44,
    24682 => 44,
    24683 => 44,
    24684 => 44,
    24685 => 44,
    24686 => 44,
    24687 => 44,
    24688 => 44,
    24689 => 44,
    24690 => 44,
    24691 => 44,
    24692 => 44,
    24693 => 44,
    24694 => 44,
    24695 => 44,
    24696 => 44,
    24697 => 44,
    24698 => 44,
    24699 => 44,
    24700 => 44,
    24701 => 44,
    24702 => 44,
    24703 => 44,
    24704 => 44,
    24705 => 44,
    24706 => 44,
    24707 => 44,
    24708 => 44,
    24709 => 44,
    24710 => 44,
    24711 => 44,
    24712 => 44,
    24713 => 44,
    24714 => 44,
    24715 => 44,
    24716 => 44,
    24717 => 44,
    24718 => 44,
    24719 => 44,
    24720 => 44,
    24721 => 44,
    24722 => 44,
    24723 => 44,
    24724 => 44,
    24725 => 44,
    24726 => 44,
    24727 => 44,
    24728 => 44,
    24729 => 44,
    24730 => 44,
    24731 => 44,
    24732 => 44,
    24733 => 44,
    24734 => 44,
    24735 => 44,
    24736 => 44,
    24737 => 44,
    24738 => 44,
    24739 => 44,
    24740 => 44,
    24741 => 44,
    24742 => 44,
    24743 => 44,
    24744 => 44,
    24745 => 44,
    24746 => 44,
    24747 => 44,
    24748 => 44,
    24749 => 44,
    24750 => 44,
    24751 => 44,
    24752 => 44,
    24753 => 44,
    24754 => 44,
    24755 => 44,
    24756 => 44,
    24757 => 44,
    24758 => 44,
    24759 => 44,
    24760 => 44,
    24761 => 44,
    24762 => 44,
    24763 => 44,
    24764 => 44,
    24765 => 44,
    24766 => 44,
    24767 => 44,
    24768 => 44,
    24769 => 44,
    24770 => 44,
    24771 => 44,
    24772 => 44,
    24773 => 44,
    24774 => 44,
    24775 => 44,
    24776 => 44,
    24777 => 44,
    24778 => 44,
    24779 => 44,
    24780 => 44,
    24781 => 44,
    24782 => 44,
    24783 => 44,
    24784 => 44,
    24785 => 44,
    24786 => 44,
    24787 => 44,
    24788 => 44,
    24789 => 44,
    24790 => 44,
    24791 => 44,
    24792 => 44,
    24793 => 44,
    24794 => 44,
    24795 => 44,
    24796 => 44,
    24797 => 44,
    24798 => 44,
    24799 => 44,
    24800 => 44,
    24801 => 44,
    24802 => 44,
    24803 => 44,
    24804 => 44,
    24805 => 44,
    24806 => 44,
    24807 => 44,
    24808 => 44,
    24809 => 44,
    24810 => 44,
    24811 => 44,
    24812 => 44,
    24813 => 44,
    24814 => 44,
    24815 => 44,
    24816 => 44,
    24817 => 44,
    24818 => 44,
    24819 => 43,
    24820 => 43,
    24821 => 43,
    24822 => 43,
    24823 => 43,
    24824 => 43,
    24825 => 43,
    24826 => 43,
    24827 => 43,
    24828 => 43,
    24829 => 43,
    24830 => 43,
    24831 => 43,
    24832 => 43,
    24833 => 43,
    24834 => 43,
    24835 => 43,
    24836 => 43,
    24837 => 43,
    24838 => 43,
    24839 => 43,
    24840 => 43,
    24841 => 43,
    24842 => 43,
    24843 => 43,
    24844 => 43,
    24845 => 43,
    24846 => 43,
    24847 => 43,
    24848 => 43,
    24849 => 43,
    24850 => 43,
    24851 => 43,
    24852 => 43,
    24853 => 43,
    24854 => 43,
    24855 => 43,
    24856 => 43,
    24857 => 43,
    24858 => 43,
    24859 => 43,
    24860 => 43,
    24861 => 43,
    24862 => 43,
    24863 => 43,
    24864 => 43,
    24865 => 43,
    24866 => 43,
    24867 => 43,
    24868 => 43,
    24869 => 43,
    24870 => 43,
    24871 => 43,
    24872 => 43,
    24873 => 43,
    24874 => 43,
    24875 => 43,
    24876 => 43,
    24877 => 43,
    24878 => 43,
    24879 => 43,
    24880 => 43,
    24881 => 43,
    24882 => 43,
    24883 => 43,
    24884 => 43,
    24885 => 43,
    24886 => 43,
    24887 => 43,
    24888 => 43,
    24889 => 43,
    24890 => 43,
    24891 => 43,
    24892 => 43,
    24893 => 43,
    24894 => 43,
    24895 => 43,
    24896 => 43,
    24897 => 43,
    24898 => 43,
    24899 => 43,
    24900 => 43,
    24901 => 43,
    24902 => 43,
    24903 => 43,
    24904 => 43,
    24905 => 43,
    24906 => 43,
    24907 => 43,
    24908 => 43,
    24909 => 43,
    24910 => 43,
    24911 => 43,
    24912 => 43,
    24913 => 43,
    24914 => 43,
    24915 => 43,
    24916 => 43,
    24917 => 43,
    24918 => 43,
    24919 => 43,
    24920 => 43,
    24921 => 43,
    24922 => 43,
    24923 => 43,
    24924 => 43,
    24925 => 43,
    24926 => 43,
    24927 => 43,
    24928 => 43,
    24929 => 43,
    24930 => 43,
    24931 => 43,
    24932 => 43,
    24933 => 43,
    24934 => 43,
    24935 => 43,
    24936 => 43,
    24937 => 43,
    24938 => 43,
    24939 => 43,
    24940 => 43,
    24941 => 43,
    24942 => 43,
    24943 => 43,
    24944 => 43,
    24945 => 43,
    24946 => 43,
    24947 => 43,
    24948 => 43,
    24949 => 43,
    24950 => 43,
    24951 => 43,
    24952 => 43,
    24953 => 43,
    24954 => 43,
    24955 => 43,
    24956 => 43,
    24957 => 43,
    24958 => 43,
    24959 => 43,
    24960 => 43,
    24961 => 43,
    24962 => 43,
    24963 => 43,
    24964 => 43,
    24965 => 43,
    24966 => 43,
    24967 => 43,
    24968 => 43,
    24969 => 43,
    24970 => 43,
    24971 => 43,
    24972 => 43,
    24973 => 43,
    24974 => 43,
    24975 => 43,
    24976 => 43,
    24977 => 43,
    24978 => 43,
    24979 => 43,
    24980 => 43,
    24981 => 43,
    24982 => 43,
    24983 => 43,
    24984 => 43,
    24985 => 43,
    24986 => 43,
    24987 => 43,
    24988 => 43,
    24989 => 43,
    24990 => 43,
    24991 => 43,
    24992 => 43,
    24993 => 43,
    24994 => 43,
    24995 => 43,
    24996 => 43,
    24997 => 43,
    24998 => 43,
    24999 => 43,
    25000 => 43,
    25001 => 43,
    25002 => 43,
    25003 => 43,
    25004 => 43,
    25005 => 43,
    25006 => 43,
    25007 => 43,
    25008 => 43,
    25009 => 43,
    25010 => 43,
    25011 => 43,
    25012 => 43,
    25013 => 43,
    25014 => 43,
    25015 => 43,
    25016 => 43,
    25017 => 43,
    25018 => 43,
    25019 => 43,
    25020 => 43,
    25021 => 43,
    25022 => 43,
    25023 => 43,
    25024 => 43,
    25025 => 43,
    25026 => 43,
    25027 => 43,
    25028 => 43,
    25029 => 43,
    25030 => 43,
    25031 => 43,
    25032 => 43,
    25033 => 43,
    25034 => 43,
    25035 => 43,
    25036 => 43,
    25037 => 43,
    25038 => 43,
    25039 => 43,
    25040 => 43,
    25041 => 43,
    25042 => 43,
    25043 => 43,
    25044 => 43,
    25045 => 43,
    25046 => 42,
    25047 => 42,
    25048 => 42,
    25049 => 42,
    25050 => 42,
    25051 => 42,
    25052 => 42,
    25053 => 42,
    25054 => 42,
    25055 => 42,
    25056 => 42,
    25057 => 42,
    25058 => 42,
    25059 => 42,
    25060 => 42,
    25061 => 42,
    25062 => 42,
    25063 => 42,
    25064 => 42,
    25065 => 42,
    25066 => 42,
    25067 => 42,
    25068 => 42,
    25069 => 42,
    25070 => 42,
    25071 => 42,
    25072 => 42,
    25073 => 42,
    25074 => 42,
    25075 => 42,
    25076 => 42,
    25077 => 42,
    25078 => 42,
    25079 => 42,
    25080 => 42,
    25081 => 42,
    25082 => 42,
    25083 => 42,
    25084 => 42,
    25085 => 42,
    25086 => 42,
    25087 => 42,
    25088 => 42,
    25089 => 42,
    25090 => 42,
    25091 => 42,
    25092 => 42,
    25093 => 42,
    25094 => 42,
    25095 => 42,
    25096 => 42,
    25097 => 42,
    25098 => 42,
    25099 => 42,
    25100 => 42,
    25101 => 42,
    25102 => 42,
    25103 => 42,
    25104 => 42,
    25105 => 42,
    25106 => 42,
    25107 => 42,
    25108 => 42,
    25109 => 42,
    25110 => 42,
    25111 => 42,
    25112 => 42,
    25113 => 42,
    25114 => 42,
    25115 => 42,
    25116 => 42,
    25117 => 42,
    25118 => 42,
    25119 => 42,
    25120 => 42,
    25121 => 42,
    25122 => 42,
    25123 => 42,
    25124 => 42,
    25125 => 42,
    25126 => 42,
    25127 => 42,
    25128 => 42,
    25129 => 42,
    25130 => 42,
    25131 => 42,
    25132 => 42,
    25133 => 42,
    25134 => 42,
    25135 => 42,
    25136 => 42,
    25137 => 42,
    25138 => 42,
    25139 => 42,
    25140 => 42,
    25141 => 42,
    25142 => 42,
    25143 => 42,
    25144 => 42,
    25145 => 42,
    25146 => 42,
    25147 => 42,
    25148 => 42,
    25149 => 42,
    25150 => 42,
    25151 => 42,
    25152 => 42,
    25153 => 42,
    25154 => 42,
    25155 => 42,
    25156 => 42,
    25157 => 42,
    25158 => 42,
    25159 => 42,
    25160 => 42,
    25161 => 42,
    25162 => 42,
    25163 => 42,
    25164 => 42,
    25165 => 42,
    25166 => 42,
    25167 => 42,
    25168 => 42,
    25169 => 42,
    25170 => 42,
    25171 => 42,
    25172 => 42,
    25173 => 42,
    25174 => 42,
    25175 => 42,
    25176 => 42,
    25177 => 42,
    25178 => 42,
    25179 => 42,
    25180 => 42,
    25181 => 42,
    25182 => 42,
    25183 => 42,
    25184 => 42,
    25185 => 42,
    25186 => 42,
    25187 => 42,
    25188 => 42,
    25189 => 42,
    25190 => 42,
    25191 => 42,
    25192 => 42,
    25193 => 42,
    25194 => 42,
    25195 => 42,
    25196 => 42,
    25197 => 42,
    25198 => 42,
    25199 => 42,
    25200 => 42,
    25201 => 42,
    25202 => 42,
    25203 => 42,
    25204 => 42,
    25205 => 42,
    25206 => 42,
    25207 => 42,
    25208 => 42,
    25209 => 42,
    25210 => 42,
    25211 => 42,
    25212 => 42,
    25213 => 42,
    25214 => 42,
    25215 => 42,
    25216 => 42,
    25217 => 42,
    25218 => 42,
    25219 => 42,
    25220 => 42,
    25221 => 42,
    25222 => 42,
    25223 => 42,
    25224 => 42,
    25225 => 42,
    25226 => 42,
    25227 => 42,
    25228 => 42,
    25229 => 42,
    25230 => 42,
    25231 => 42,
    25232 => 42,
    25233 => 42,
    25234 => 42,
    25235 => 42,
    25236 => 42,
    25237 => 42,
    25238 => 42,
    25239 => 42,
    25240 => 42,
    25241 => 42,
    25242 => 42,
    25243 => 42,
    25244 => 42,
    25245 => 42,
    25246 => 42,
    25247 => 42,
    25248 => 42,
    25249 => 42,
    25250 => 42,
    25251 => 42,
    25252 => 42,
    25253 => 42,
    25254 => 42,
    25255 => 42,
    25256 => 42,
    25257 => 42,
    25258 => 42,
    25259 => 42,
    25260 => 42,
    25261 => 42,
    25262 => 42,
    25263 => 42,
    25264 => 42,
    25265 => 42,
    25266 => 42,
    25267 => 42,
    25268 => 41,
    25269 => 41,
    25270 => 41,
    25271 => 41,
    25272 => 41,
    25273 => 41,
    25274 => 41,
    25275 => 41,
    25276 => 41,
    25277 => 41,
    25278 => 41,
    25279 => 41,
    25280 => 41,
    25281 => 41,
    25282 => 41,
    25283 => 41,
    25284 => 41,
    25285 => 41,
    25286 => 41,
    25287 => 41,
    25288 => 41,
    25289 => 41,
    25290 => 41,
    25291 => 41,
    25292 => 41,
    25293 => 41,
    25294 => 41,
    25295 => 41,
    25296 => 41,
    25297 => 41,
    25298 => 41,
    25299 => 41,
    25300 => 41,
    25301 => 41,
    25302 => 41,
    25303 => 41,
    25304 => 41,
    25305 => 41,
    25306 => 41,
    25307 => 41,
    25308 => 41,
    25309 => 41,
    25310 => 41,
    25311 => 41,
    25312 => 41,
    25313 => 41,
    25314 => 41,
    25315 => 41,
    25316 => 41,
    25317 => 41,
    25318 => 41,
    25319 => 41,
    25320 => 41,
    25321 => 41,
    25322 => 41,
    25323 => 41,
    25324 => 41,
    25325 => 41,
    25326 => 41,
    25327 => 41,
    25328 => 41,
    25329 => 41,
    25330 => 41,
    25331 => 41,
    25332 => 41,
    25333 => 41,
    25334 => 41,
    25335 => 41,
    25336 => 41,
    25337 => 41,
    25338 => 41,
    25339 => 41,
    25340 => 41,
    25341 => 41,
    25342 => 41,
    25343 => 41,
    25344 => 41,
    25345 => 41,
    25346 => 41,
    25347 => 41,
    25348 => 41,
    25349 => 41,
    25350 => 41,
    25351 => 41,
    25352 => 41,
    25353 => 41,
    25354 => 41,
    25355 => 41,
    25356 => 41,
    25357 => 41,
    25358 => 41,
    25359 => 41,
    25360 => 41,
    25361 => 41,
    25362 => 41,
    25363 => 41,
    25364 => 41,
    25365 => 41,
    25366 => 41,
    25367 => 41,
    25368 => 41,
    25369 => 41,
    25370 => 41,
    25371 => 41,
    25372 => 41,
    25373 => 41,
    25374 => 41,
    25375 => 41,
    25376 => 41,
    25377 => 41,
    25378 => 41,
    25379 => 41,
    25380 => 41,
    25381 => 41,
    25382 => 41,
    25383 => 41,
    25384 => 41,
    25385 => 41,
    25386 => 41,
    25387 => 41,
    25388 => 41,
    25389 => 41,
    25390 => 41,
    25391 => 41,
    25392 => 41,
    25393 => 41,
    25394 => 41,
    25395 => 41,
    25396 => 41,
    25397 => 41,
    25398 => 41,
    25399 => 41,
    25400 => 41,
    25401 => 41,
    25402 => 41,
    25403 => 41,
    25404 => 41,
    25405 => 41,
    25406 => 41,
    25407 => 41,
    25408 => 41,
    25409 => 41,
    25410 => 41,
    25411 => 41,
    25412 => 41,
    25413 => 41,
    25414 => 41,
    25415 => 41,
    25416 => 41,
    25417 => 41,
    25418 => 41,
    25419 => 41,
    25420 => 41,
    25421 => 41,
    25422 => 41,
    25423 => 41,
    25424 => 41,
    25425 => 41,
    25426 => 41,
    25427 => 41,
    25428 => 41,
    25429 => 41,
    25430 => 41,
    25431 => 41,
    25432 => 41,
    25433 => 41,
    25434 => 41,
    25435 => 41,
    25436 => 41,
    25437 => 41,
    25438 => 41,
    25439 => 41,
    25440 => 41,
    25441 => 41,
    25442 => 41,
    25443 => 41,
    25444 => 41,
    25445 => 41,
    25446 => 41,
    25447 => 41,
    25448 => 41,
    25449 => 41,
    25450 => 41,
    25451 => 41,
    25452 => 41,
    25453 => 41,
    25454 => 41,
    25455 => 41,
    25456 => 41,
    25457 => 41,
    25458 => 41,
    25459 => 41,
    25460 => 41,
    25461 => 41,
    25462 => 41,
    25463 => 41,
    25464 => 41,
    25465 => 41,
    25466 => 41,
    25467 => 41,
    25468 => 41,
    25469 => 41,
    25470 => 41,
    25471 => 41,
    25472 => 41,
    25473 => 41,
    25474 => 41,
    25475 => 41,
    25476 => 41,
    25477 => 41,
    25478 => 41,
    25479 => 41,
    25480 => 41,
    25481 => 41,
    25482 => 41,
    25483 => 41,
    25484 => 41,
    25485 => 41,
    25486 => 40,
    25487 => 40,
    25488 => 40,
    25489 => 40,
    25490 => 40,
    25491 => 40,
    25492 => 40,
    25493 => 40,
    25494 => 40,
    25495 => 40,
    25496 => 40,
    25497 => 40,
    25498 => 40,
    25499 => 40,
    25500 => 40,
    25501 => 40,
    25502 => 40,
    25503 => 40,
    25504 => 40,
    25505 => 40,
    25506 => 40,
    25507 => 40,
    25508 => 40,
    25509 => 40,
    25510 => 40,
    25511 => 40,
    25512 => 40,
    25513 => 40,
    25514 => 40,
    25515 => 40,
    25516 => 40,
    25517 => 40,
    25518 => 40,
    25519 => 40,
    25520 => 40,
    25521 => 40,
    25522 => 40,
    25523 => 40,
    25524 => 40,
    25525 => 40,
    25526 => 40,
    25527 => 40,
    25528 => 40,
    25529 => 40,
    25530 => 40,
    25531 => 40,
    25532 => 40,
    25533 => 40,
    25534 => 40,
    25535 => 40,
    25536 => 40,
    25537 => 40,
    25538 => 40,
    25539 => 40,
    25540 => 40,
    25541 => 40,
    25542 => 40,
    25543 => 40,
    25544 => 40,
    25545 => 40,
    25546 => 40,
    25547 => 40,
    25548 => 40,
    25549 => 40,
    25550 => 40,
    25551 => 40,
    25552 => 40,
    25553 => 40,
    25554 => 40,
    25555 => 40,
    25556 => 40,
    25557 => 40,
    25558 => 40,
    25559 => 40,
    25560 => 40,
    25561 => 40,
    25562 => 40,
    25563 => 40,
    25564 => 40,
    25565 => 40,
    25566 => 40,
    25567 => 40,
    25568 => 40,
    25569 => 40,
    25570 => 40,
    25571 => 40,
    25572 => 40,
    25573 => 40,
    25574 => 40,
    25575 => 40,
    25576 => 40,
    25577 => 40,
    25578 => 40,
    25579 => 40,
    25580 => 40,
    25581 => 40,
    25582 => 40,
    25583 => 40,
    25584 => 40,
    25585 => 40,
    25586 => 40,
    25587 => 40,
    25588 => 40,
    25589 => 40,
    25590 => 40,
    25591 => 40,
    25592 => 40,
    25593 => 40,
    25594 => 40,
    25595 => 40,
    25596 => 40,
    25597 => 40,
    25598 => 40,
    25599 => 40,
    25600 => 40,
    25601 => 40,
    25602 => 40,
    25603 => 40,
    25604 => 40,
    25605 => 40,
    25606 => 40,
    25607 => 40,
    25608 => 40,
    25609 => 40,
    25610 => 40,
    25611 => 40,
    25612 => 40,
    25613 => 40,
    25614 => 40,
    25615 => 40,
    25616 => 40,
    25617 => 40,
    25618 => 40,
    25619 => 40,
    25620 => 40,
    25621 => 40,
    25622 => 40,
    25623 => 40,
    25624 => 40,
    25625 => 40,
    25626 => 40,
    25627 => 40,
    25628 => 40,
    25629 => 40,
    25630 => 40,
    25631 => 40,
    25632 => 40,
    25633 => 40,
    25634 => 40,
    25635 => 40,
    25636 => 40,
    25637 => 40,
    25638 => 40,
    25639 => 40,
    25640 => 40,
    25641 => 40,
    25642 => 40,
    25643 => 40,
    25644 => 40,
    25645 => 40,
    25646 => 40,
    25647 => 40,
    25648 => 40,
    25649 => 40,
    25650 => 40,
    25651 => 40,
    25652 => 40,
    25653 => 40,
    25654 => 40,
    25655 => 40,
    25656 => 40,
    25657 => 40,
    25658 => 40,
    25659 => 40,
    25660 => 40,
    25661 => 40,
    25662 => 40,
    25663 => 40,
    25664 => 40,
    25665 => 40,
    25666 => 40,
    25667 => 40,
    25668 => 40,
    25669 => 40,
    25670 => 40,
    25671 => 40,
    25672 => 40,
    25673 => 40,
    25674 => 40,
    25675 => 40,
    25676 => 40,
    25677 => 40,
    25678 => 40,
    25679 => 40,
    25680 => 40,
    25681 => 40,
    25682 => 40,
    25683 => 40,
    25684 => 40,
    25685 => 40,
    25686 => 40,
    25687 => 40,
    25688 => 40,
    25689 => 40,
    25690 => 40,
    25691 => 40,
    25692 => 40,
    25693 => 40,
    25694 => 40,
    25695 => 40,
    25696 => 40,
    25697 => 40,
    25698 => 40,
    25699 => 40,
    25700 => 39,
    25701 => 39,
    25702 => 39,
    25703 => 39,
    25704 => 39,
    25705 => 39,
    25706 => 39,
    25707 => 39,
    25708 => 39,
    25709 => 39,
    25710 => 39,
    25711 => 39,
    25712 => 39,
    25713 => 39,
    25714 => 39,
    25715 => 39,
    25716 => 39,
    25717 => 39,
    25718 => 39,
    25719 => 39,
    25720 => 39,
    25721 => 39,
    25722 => 39,
    25723 => 39,
    25724 => 39,
    25725 => 39,
    25726 => 39,
    25727 => 39,
    25728 => 39,
    25729 => 39,
    25730 => 39,
    25731 => 39,
    25732 => 39,
    25733 => 39,
    25734 => 39,
    25735 => 39,
    25736 => 39,
    25737 => 39,
    25738 => 39,
    25739 => 39,
    25740 => 39,
    25741 => 39,
    25742 => 39,
    25743 => 39,
    25744 => 39,
    25745 => 39,
    25746 => 39,
    25747 => 39,
    25748 => 39,
    25749 => 39,
    25750 => 39,
    25751 => 39,
    25752 => 39,
    25753 => 39,
    25754 => 39,
    25755 => 39,
    25756 => 39,
    25757 => 39,
    25758 => 39,
    25759 => 39,
    25760 => 39,
    25761 => 39,
    25762 => 39,
    25763 => 39,
    25764 => 39,
    25765 => 39,
    25766 => 39,
    25767 => 39,
    25768 => 39,
    25769 => 39,
    25770 => 39,
    25771 => 39,
    25772 => 39,
    25773 => 39,
    25774 => 39,
    25775 => 39,
    25776 => 39,
    25777 => 39,
    25778 => 39,
    25779 => 39,
    25780 => 39,
    25781 => 39,
    25782 => 39,
    25783 => 39,
    25784 => 39,
    25785 => 39,
    25786 => 39,
    25787 => 39,
    25788 => 39,
    25789 => 39,
    25790 => 39,
    25791 => 39,
    25792 => 39,
    25793 => 39,
    25794 => 39,
    25795 => 39,
    25796 => 39,
    25797 => 39,
    25798 => 39,
    25799 => 39,
    25800 => 39,
    25801 => 39,
    25802 => 39,
    25803 => 39,
    25804 => 39,
    25805 => 39,
    25806 => 39,
    25807 => 39,
    25808 => 39,
    25809 => 39,
    25810 => 39,
    25811 => 39,
    25812 => 39,
    25813 => 39,
    25814 => 39,
    25815 => 39,
    25816 => 39,
    25817 => 39,
    25818 => 39,
    25819 => 39,
    25820 => 39,
    25821 => 39,
    25822 => 39,
    25823 => 39,
    25824 => 39,
    25825 => 39,
    25826 => 39,
    25827 => 39,
    25828 => 39,
    25829 => 39,
    25830 => 39,
    25831 => 39,
    25832 => 39,
    25833 => 39,
    25834 => 39,
    25835 => 39,
    25836 => 39,
    25837 => 39,
    25838 => 39,
    25839 => 39,
    25840 => 39,
    25841 => 39,
    25842 => 39,
    25843 => 39,
    25844 => 39,
    25845 => 39,
    25846 => 39,
    25847 => 39,
    25848 => 39,
    25849 => 39,
    25850 => 39,
    25851 => 39,
    25852 => 39,
    25853 => 39,
    25854 => 39,
    25855 => 39,
    25856 => 39,
    25857 => 39,
    25858 => 39,
    25859 => 39,
    25860 => 39,
    25861 => 39,
    25862 => 39,
    25863 => 39,
    25864 => 39,
    25865 => 39,
    25866 => 39,
    25867 => 39,
    25868 => 39,
    25869 => 39,
    25870 => 39,
    25871 => 39,
    25872 => 39,
    25873 => 39,
    25874 => 39,
    25875 => 39,
    25876 => 39,
    25877 => 39,
    25878 => 39,
    25879 => 39,
    25880 => 39,
    25881 => 39,
    25882 => 39,
    25883 => 39,
    25884 => 39,
    25885 => 39,
    25886 => 39,
    25887 => 39,
    25888 => 39,
    25889 => 39,
    25890 => 39,
    25891 => 39,
    25892 => 39,
    25893 => 39,
    25894 => 39,
    25895 => 39,
    25896 => 39,
    25897 => 39,
    25898 => 39,
    25899 => 39,
    25900 => 39,
    25901 => 39,
    25902 => 39,
    25903 => 39,
    25904 => 39,
    25905 => 39,
    25906 => 39,
    25907 => 39,
    25908 => 39,
    25909 => 39,
    25910 => 39,
    25911 => 38,
    25912 => 38,
    25913 => 38,
    25914 => 38,
    25915 => 38,
    25916 => 38,
    25917 => 38,
    25918 => 38,
    25919 => 38,
    25920 => 38,
    25921 => 38,
    25922 => 38,
    25923 => 38,
    25924 => 38,
    25925 => 38,
    25926 => 38,
    25927 => 38,
    25928 => 38,
    25929 => 38,
    25930 => 38,
    25931 => 38,
    25932 => 38,
    25933 => 38,
    25934 => 38,
    25935 => 38,
    25936 => 38,
    25937 => 38,
    25938 => 38,
    25939 => 38,
    25940 => 38,
    25941 => 38,
    25942 => 38,
    25943 => 38,
    25944 => 38,
    25945 => 38,
    25946 => 38,
    25947 => 38,
    25948 => 38,
    25949 => 38,
    25950 => 38,
    25951 => 38,
    25952 => 38,
    25953 => 38,
    25954 => 38,
    25955 => 38,
    25956 => 38,
    25957 => 38,
    25958 => 38,
    25959 => 38,
    25960 => 38,
    25961 => 38,
    25962 => 38,
    25963 => 38,
    25964 => 38,
    25965 => 38,
    25966 => 38,
    25967 => 38,
    25968 => 38,
    25969 => 38,
    25970 => 38,
    25971 => 38,
    25972 => 38,
    25973 => 38,
    25974 => 38,
    25975 => 38,
    25976 => 38,
    25977 => 38,
    25978 => 38,
    25979 => 38,
    25980 => 38,
    25981 => 38,
    25982 => 38,
    25983 => 38,
    25984 => 38,
    25985 => 38,
    25986 => 38,
    25987 => 38,
    25988 => 38,
    25989 => 38,
    25990 => 38,
    25991 => 38,
    25992 => 38,
    25993 => 38,
    25994 => 38,
    25995 => 38,
    25996 => 38,
    25997 => 38,
    25998 => 38,
    25999 => 38,
    26000 => 38,
    26001 => 38,
    26002 => 38,
    26003 => 38,
    26004 => 38,
    26005 => 38,
    26006 => 38,
    26007 => 38,
    26008 => 38,
    26009 => 38,
    26010 => 38,
    26011 => 38,
    26012 => 38,
    26013 => 38,
    26014 => 38,
    26015 => 38,
    26016 => 38,
    26017 => 38,
    26018 => 38,
    26019 => 38,
    26020 => 38,
    26021 => 38,
    26022 => 38,
    26023 => 38,
    26024 => 38,
    26025 => 38,
    26026 => 38,
    26027 => 38,
    26028 => 38,
    26029 => 38,
    26030 => 38,
    26031 => 38,
    26032 => 38,
    26033 => 38,
    26034 => 38,
    26035 => 38,
    26036 => 38,
    26037 => 38,
    26038 => 38,
    26039 => 38,
    26040 => 38,
    26041 => 38,
    26042 => 38,
    26043 => 38,
    26044 => 38,
    26045 => 38,
    26046 => 38,
    26047 => 38,
    26048 => 38,
    26049 => 38,
    26050 => 38,
    26051 => 38,
    26052 => 38,
    26053 => 38,
    26054 => 38,
    26055 => 38,
    26056 => 38,
    26057 => 38,
    26058 => 38,
    26059 => 38,
    26060 => 38,
    26061 => 38,
    26062 => 38,
    26063 => 38,
    26064 => 38,
    26065 => 38,
    26066 => 38,
    26067 => 38,
    26068 => 38,
    26069 => 38,
    26070 => 38,
    26071 => 38,
    26072 => 38,
    26073 => 38,
    26074 => 38,
    26075 => 38,
    26076 => 38,
    26077 => 38,
    26078 => 38,
    26079 => 38,
    26080 => 38,
    26081 => 38,
    26082 => 38,
    26083 => 38,
    26084 => 38,
    26085 => 38,
    26086 => 38,
    26087 => 38,
    26088 => 38,
    26089 => 38,
    26090 => 38,
    26091 => 38,
    26092 => 38,
    26093 => 38,
    26094 => 38,
    26095 => 38,
    26096 => 38,
    26097 => 38,
    26098 => 38,
    26099 => 38,
    26100 => 38,
    26101 => 38,
    26102 => 38,
    26103 => 38,
    26104 => 38,
    26105 => 38,
    26106 => 38,
    26107 => 38,
    26108 => 38,
    26109 => 38,
    26110 => 38,
    26111 => 38,
    26112 => 38,
    26113 => 38,
    26114 => 38,
    26115 => 38,
    26116 => 38,
    26117 => 38,
    26118 => 37,
    26119 => 37,
    26120 => 37,
    26121 => 37,
    26122 => 37,
    26123 => 37,
    26124 => 37,
    26125 => 37,
    26126 => 37,
    26127 => 37,
    26128 => 37,
    26129 => 37,
    26130 => 37,
    26131 => 37,
    26132 => 37,
    26133 => 37,
    26134 => 37,
    26135 => 37,
    26136 => 37,
    26137 => 37,
    26138 => 37,
    26139 => 37,
    26140 => 37,
    26141 => 37,
    26142 => 37,
    26143 => 37,
    26144 => 37,
    26145 => 37,
    26146 => 37,
    26147 => 37,
    26148 => 37,
    26149 => 37,
    26150 => 37,
    26151 => 37,
    26152 => 37,
    26153 => 37,
    26154 => 37,
    26155 => 37,
    26156 => 37,
    26157 => 37,
    26158 => 37,
    26159 => 37,
    26160 => 37,
    26161 => 37,
    26162 => 37,
    26163 => 37,
    26164 => 37,
    26165 => 37,
    26166 => 37,
    26167 => 37,
    26168 => 37,
    26169 => 37,
    26170 => 37,
    26171 => 37,
    26172 => 37,
    26173 => 37,
    26174 => 37,
    26175 => 37,
    26176 => 37,
    26177 => 37,
    26178 => 37,
    26179 => 37,
    26180 => 37,
    26181 => 37,
    26182 => 37,
    26183 => 37,
    26184 => 37,
    26185 => 37,
    26186 => 37,
    26187 => 37,
    26188 => 37,
    26189 => 37,
    26190 => 37,
    26191 => 37,
    26192 => 37,
    26193 => 37,
    26194 => 37,
    26195 => 37,
    26196 => 37,
    26197 => 37,
    26198 => 37,
    26199 => 37,
    26200 => 37,
    26201 => 37,
    26202 => 37,
    26203 => 37,
    26204 => 37,
    26205 => 37,
    26206 => 37,
    26207 => 37,
    26208 => 37,
    26209 => 37,
    26210 => 37,
    26211 => 37,
    26212 => 37,
    26213 => 37,
    26214 => 37,
    26215 => 37,
    26216 => 37,
    26217 => 37,
    26218 => 37,
    26219 => 37,
    26220 => 37,
    26221 => 37,
    26222 => 37,
    26223 => 37,
    26224 => 37,
    26225 => 37,
    26226 => 37,
    26227 => 37,
    26228 => 37,
    26229 => 37,
    26230 => 37,
    26231 => 37,
    26232 => 37,
    26233 => 37,
    26234 => 37,
    26235 => 37,
    26236 => 37,
    26237 => 37,
    26238 => 37,
    26239 => 37,
    26240 => 37,
    26241 => 37,
    26242 => 37,
    26243 => 37,
    26244 => 37,
    26245 => 37,
    26246 => 37,
    26247 => 37,
    26248 => 37,
    26249 => 37,
    26250 => 37,
    26251 => 37,
    26252 => 37,
    26253 => 37,
    26254 => 37,
    26255 => 37,
    26256 => 37,
    26257 => 37,
    26258 => 37,
    26259 => 37,
    26260 => 37,
    26261 => 37,
    26262 => 37,
    26263 => 37,
    26264 => 37,
    26265 => 37,
    26266 => 37,
    26267 => 37,
    26268 => 37,
    26269 => 37,
    26270 => 37,
    26271 => 37,
    26272 => 37,
    26273 => 37,
    26274 => 37,
    26275 => 37,
    26276 => 37,
    26277 => 37,
    26278 => 37,
    26279 => 37,
    26280 => 37,
    26281 => 37,
    26282 => 37,
    26283 => 37,
    26284 => 37,
    26285 => 37,
    26286 => 37,
    26287 => 37,
    26288 => 37,
    26289 => 37,
    26290 => 37,
    26291 => 37,
    26292 => 37,
    26293 => 37,
    26294 => 37,
    26295 => 37,
    26296 => 37,
    26297 => 37,
    26298 => 37,
    26299 => 37,
    26300 => 37,
    26301 => 37,
    26302 => 37,
    26303 => 37,
    26304 => 37,
    26305 => 37,
    26306 => 37,
    26307 => 37,
    26308 => 37,
    26309 => 37,
    26310 => 37,
    26311 => 37,
    26312 => 37,
    26313 => 37,
    26314 => 37,
    26315 => 37,
    26316 => 37,
    26317 => 37,
    26318 => 37,
    26319 => 37,
    26320 => 37,
    26321 => 37,
    26322 => 37,
    26323 => 36,
    26324 => 36,
    26325 => 36,
    26326 => 36,
    26327 => 36,
    26328 => 36,
    26329 => 36,
    26330 => 36,
    26331 => 36,
    26332 => 36,
    26333 => 36,
    26334 => 36,
    26335 => 36,
    26336 => 36,
    26337 => 36,
    26338 => 36,
    26339 => 36,
    26340 => 36,
    26341 => 36,
    26342 => 36,
    26343 => 36,
    26344 => 36,
    26345 => 36,
    26346 => 36,
    26347 => 36,
    26348 => 36,
    26349 => 36,
    26350 => 36,
    26351 => 36,
    26352 => 36,
    26353 => 36,
    26354 => 36,
    26355 => 36,
    26356 => 36,
    26357 => 36,
    26358 => 36,
    26359 => 36,
    26360 => 36,
    26361 => 36,
    26362 => 36,
    26363 => 36,
    26364 => 36,
    26365 => 36,
    26366 => 36,
    26367 => 36,
    26368 => 36,
    26369 => 36,
    26370 => 36,
    26371 => 36,
    26372 => 36,
    26373 => 36,
    26374 => 36,
    26375 => 36,
    26376 => 36,
    26377 => 36,
    26378 => 36,
    26379 => 36,
    26380 => 36,
    26381 => 36,
    26382 => 36,
    26383 => 36,
    26384 => 36,
    26385 => 36,
    26386 => 36,
    26387 => 36,
    26388 => 36,
    26389 => 36,
    26390 => 36,
    26391 => 36,
    26392 => 36,
    26393 => 36,
    26394 => 36,
    26395 => 36,
    26396 => 36,
    26397 => 36,
    26398 => 36,
    26399 => 36,
    26400 => 36,
    26401 => 36,
    26402 => 36,
    26403 => 36,
    26404 => 36,
    26405 => 36,
    26406 => 36,
    26407 => 36,
    26408 => 36,
    26409 => 36,
    26410 => 36,
    26411 => 36,
    26412 => 36,
    26413 => 36,
    26414 => 36,
    26415 => 36,
    26416 => 36,
    26417 => 36,
    26418 => 36,
    26419 => 36,
    26420 => 36,
    26421 => 36,
    26422 => 36,
    26423 => 36,
    26424 => 36,
    26425 => 36,
    26426 => 36,
    26427 => 36,
    26428 => 36,
    26429 => 36,
    26430 => 36,
    26431 => 36,
    26432 => 36,
    26433 => 36,
    26434 => 36,
    26435 => 36,
    26436 => 36,
    26437 => 36,
    26438 => 36,
    26439 => 36,
    26440 => 36,
    26441 => 36,
    26442 => 36,
    26443 => 36,
    26444 => 36,
    26445 => 36,
    26446 => 36,
    26447 => 36,
    26448 => 36,
    26449 => 36,
    26450 => 36,
    26451 => 36,
    26452 => 36,
    26453 => 36,
    26454 => 36,
    26455 => 36,
    26456 => 36,
    26457 => 36,
    26458 => 36,
    26459 => 36,
    26460 => 36,
    26461 => 36,
    26462 => 36,
    26463 => 36,
    26464 => 36,
    26465 => 36,
    26466 => 36,
    26467 => 36,
    26468 => 36,
    26469 => 36,
    26470 => 36,
    26471 => 36,
    26472 => 36,
    26473 => 36,
    26474 => 36,
    26475 => 36,
    26476 => 36,
    26477 => 36,
    26478 => 36,
    26479 => 36,
    26480 => 36,
    26481 => 36,
    26482 => 36,
    26483 => 36,
    26484 => 36,
    26485 => 36,
    26486 => 36,
    26487 => 36,
    26488 => 36,
    26489 => 36,
    26490 => 36,
    26491 => 36,
    26492 => 36,
    26493 => 36,
    26494 => 36,
    26495 => 36,
    26496 => 36,
    26497 => 36,
    26498 => 36,
    26499 => 36,
    26500 => 36,
    26501 => 36,
    26502 => 36,
    26503 => 36,
    26504 => 36,
    26505 => 36,
    26506 => 36,
    26507 => 36,
    26508 => 36,
    26509 => 36,
    26510 => 36,
    26511 => 36,
    26512 => 36,
    26513 => 36,
    26514 => 36,
    26515 => 36,
    26516 => 36,
    26517 => 36,
    26518 => 36,
    26519 => 36,
    26520 => 36,
    26521 => 36,
    26522 => 36,
    26523 => 36,
    26524 => 36,
    26525 => 35,
    26526 => 35,
    26527 => 35,
    26528 => 35,
    26529 => 35,
    26530 => 35,
    26531 => 35,
    26532 => 35,
    26533 => 35,
    26534 => 35,
    26535 => 35,
    26536 => 35,
    26537 => 35,
    26538 => 35,
    26539 => 35,
    26540 => 35,
    26541 => 35,
    26542 => 35,
    26543 => 35,
    26544 => 35,
    26545 => 35,
    26546 => 35,
    26547 => 35,
    26548 => 35,
    26549 => 35,
    26550 => 35,
    26551 => 35,
    26552 => 35,
    26553 => 35,
    26554 => 35,
    26555 => 35,
    26556 => 35,
    26557 => 35,
    26558 => 35,
    26559 => 35,
    26560 => 35,
    26561 => 35,
    26562 => 35,
    26563 => 35,
    26564 => 35,
    26565 => 35,
    26566 => 35,
    26567 => 35,
    26568 => 35,
    26569 => 35,
    26570 => 35,
    26571 => 35,
    26572 => 35,
    26573 => 35,
    26574 => 35,
    26575 => 35,
    26576 => 35,
    26577 => 35,
    26578 => 35,
    26579 => 35,
    26580 => 35,
    26581 => 35,
    26582 => 35,
    26583 => 35,
    26584 => 35,
    26585 => 35,
    26586 => 35,
    26587 => 35,
    26588 => 35,
    26589 => 35,
    26590 => 35,
    26591 => 35,
    26592 => 35,
    26593 => 35,
    26594 => 35,
    26595 => 35,
    26596 => 35,
    26597 => 35,
    26598 => 35,
    26599 => 35,
    26600 => 35,
    26601 => 35,
    26602 => 35,
    26603 => 35,
    26604 => 35,
    26605 => 35,
    26606 => 35,
    26607 => 35,
    26608 => 35,
    26609 => 35,
    26610 => 35,
    26611 => 35,
    26612 => 35,
    26613 => 35,
    26614 => 35,
    26615 => 35,
    26616 => 35,
    26617 => 35,
    26618 => 35,
    26619 => 35,
    26620 => 35,
    26621 => 35,
    26622 => 35,
    26623 => 35,
    26624 => 35,
    26625 => 35,
    26626 => 35,
    26627 => 35,
    26628 => 35,
    26629 => 35,
    26630 => 35,
    26631 => 35,
    26632 => 35,
    26633 => 35,
    26634 => 35,
    26635 => 35,
    26636 => 35,
    26637 => 35,
    26638 => 35,
    26639 => 35,
    26640 => 35,
    26641 => 35,
    26642 => 35,
    26643 => 35,
    26644 => 35,
    26645 => 35,
    26646 => 35,
    26647 => 35,
    26648 => 35,
    26649 => 35,
    26650 => 35,
    26651 => 35,
    26652 => 35,
    26653 => 35,
    26654 => 35,
    26655 => 35,
    26656 => 35,
    26657 => 35,
    26658 => 35,
    26659 => 35,
    26660 => 35,
    26661 => 35,
    26662 => 35,
    26663 => 35,
    26664 => 35,
    26665 => 35,
    26666 => 35,
    26667 => 35,
    26668 => 35,
    26669 => 35,
    26670 => 35,
    26671 => 35,
    26672 => 35,
    26673 => 35,
    26674 => 35,
    26675 => 35,
    26676 => 35,
    26677 => 35,
    26678 => 35,
    26679 => 35,
    26680 => 35,
    26681 => 35,
    26682 => 35,
    26683 => 35,
    26684 => 35,
    26685 => 35,
    26686 => 35,
    26687 => 35,
    26688 => 35,
    26689 => 35,
    26690 => 35,
    26691 => 35,
    26692 => 35,
    26693 => 35,
    26694 => 35,
    26695 => 35,
    26696 => 35,
    26697 => 35,
    26698 => 35,
    26699 => 35,
    26700 => 35,
    26701 => 35,
    26702 => 35,
    26703 => 35,
    26704 => 35,
    26705 => 35,
    26706 => 35,
    26707 => 35,
    26708 => 35,
    26709 => 35,
    26710 => 35,
    26711 => 35,
    26712 => 35,
    26713 => 35,
    26714 => 35,
    26715 => 35,
    26716 => 35,
    26717 => 35,
    26718 => 35,
    26719 => 35,
    26720 => 35,
    26721 => 35,
    26722 => 35,
    26723 => 35,
    26724 => 34,
    26725 => 34,
    26726 => 34,
    26727 => 34,
    26728 => 34,
    26729 => 34,
    26730 => 34,
    26731 => 34,
    26732 => 34,
    26733 => 34,
    26734 => 34,
    26735 => 34,
    26736 => 34,
    26737 => 34,
    26738 => 34,
    26739 => 34,
    26740 => 34,
    26741 => 34,
    26742 => 34,
    26743 => 34,
    26744 => 34,
    26745 => 34,
    26746 => 34,
    26747 => 34,
    26748 => 34,
    26749 => 34,
    26750 => 34,
    26751 => 34,
    26752 => 34,
    26753 => 34,
    26754 => 34,
    26755 => 34,
    26756 => 34,
    26757 => 34,
    26758 => 34,
    26759 => 34,
    26760 => 34,
    26761 => 34,
    26762 => 34,
    26763 => 34,
    26764 => 34,
    26765 => 34,
    26766 => 34,
    26767 => 34,
    26768 => 34,
    26769 => 34,
    26770 => 34,
    26771 => 34,
    26772 => 34,
    26773 => 34,
    26774 => 34,
    26775 => 34,
    26776 => 34,
    26777 => 34,
    26778 => 34,
    26779 => 34,
    26780 => 34,
    26781 => 34,
    26782 => 34,
    26783 => 34,
    26784 => 34,
    26785 => 34,
    26786 => 34,
    26787 => 34,
    26788 => 34,
    26789 => 34,
    26790 => 34,
    26791 => 34,
    26792 => 34,
    26793 => 34,
    26794 => 34,
    26795 => 34,
    26796 => 34,
    26797 => 34,
    26798 => 34,
    26799 => 34,
    26800 => 34,
    26801 => 34,
    26802 => 34,
    26803 => 34,
    26804 => 34,
    26805 => 34,
    26806 => 34,
    26807 => 34,
    26808 => 34,
    26809 => 34,
    26810 => 34,
    26811 => 34,
    26812 => 34,
    26813 => 34,
    26814 => 34,
    26815 => 34,
    26816 => 34,
    26817 => 34,
    26818 => 34,
    26819 => 34,
    26820 => 34,
    26821 => 34,
    26822 => 34,
    26823 => 34,
    26824 => 34,
    26825 => 34,
    26826 => 34,
    26827 => 34,
    26828 => 34,
    26829 => 34,
    26830 => 34,
    26831 => 34,
    26832 => 34,
    26833 => 34,
    26834 => 34,
    26835 => 34,
    26836 => 34,
    26837 => 34,
    26838 => 34,
    26839 => 34,
    26840 => 34,
    26841 => 34,
    26842 => 34,
    26843 => 34,
    26844 => 34,
    26845 => 34,
    26846 => 34,
    26847 => 34,
    26848 => 34,
    26849 => 34,
    26850 => 34,
    26851 => 34,
    26852 => 34,
    26853 => 34,
    26854 => 34,
    26855 => 34,
    26856 => 34,
    26857 => 34,
    26858 => 34,
    26859 => 34,
    26860 => 34,
    26861 => 34,
    26862 => 34,
    26863 => 34,
    26864 => 34,
    26865 => 34,
    26866 => 34,
    26867 => 34,
    26868 => 34,
    26869 => 34,
    26870 => 34,
    26871 => 34,
    26872 => 34,
    26873 => 34,
    26874 => 34,
    26875 => 34,
    26876 => 34,
    26877 => 34,
    26878 => 34,
    26879 => 34,
    26880 => 34,
    26881 => 34,
    26882 => 34,
    26883 => 34,
    26884 => 34,
    26885 => 34,
    26886 => 34,
    26887 => 34,
    26888 => 34,
    26889 => 34,
    26890 => 34,
    26891 => 34,
    26892 => 34,
    26893 => 34,
    26894 => 34,
    26895 => 34,
    26896 => 34,
    26897 => 34,
    26898 => 34,
    26899 => 34,
    26900 => 34,
    26901 => 34,
    26902 => 34,
    26903 => 34,
    26904 => 34,
    26905 => 34,
    26906 => 34,
    26907 => 34,
    26908 => 34,
    26909 => 34,
    26910 => 34,
    26911 => 34,
    26912 => 34,
    26913 => 34,
    26914 => 34,
    26915 => 34,
    26916 => 34,
    26917 => 34,
    26918 => 34,
    26919 => 34,
    26920 => 34,
    26921 => 33,
    26922 => 33,
    26923 => 33,
    26924 => 33,
    26925 => 33,
    26926 => 33,
    26927 => 33,
    26928 => 33,
    26929 => 33,
    26930 => 33,
    26931 => 33,
    26932 => 33,
    26933 => 33,
    26934 => 33,
    26935 => 33,
    26936 => 33,
    26937 => 33,
    26938 => 33,
    26939 => 33,
    26940 => 33,
    26941 => 33,
    26942 => 33,
    26943 => 33,
    26944 => 33,
    26945 => 33,
    26946 => 33,
    26947 => 33,
    26948 => 33,
    26949 => 33,
    26950 => 33,
    26951 => 33,
    26952 => 33,
    26953 => 33,
    26954 => 33,
    26955 => 33,
    26956 => 33,
    26957 => 33,
    26958 => 33,
    26959 => 33,
    26960 => 33,
    26961 => 33,
    26962 => 33,
    26963 => 33,
    26964 => 33,
    26965 => 33,
    26966 => 33,
    26967 => 33,
    26968 => 33,
    26969 => 33,
    26970 => 33,
    26971 => 33,
    26972 => 33,
    26973 => 33,
    26974 => 33,
    26975 => 33,
    26976 => 33,
    26977 => 33,
    26978 => 33,
    26979 => 33,
    26980 => 33,
    26981 => 33,
    26982 => 33,
    26983 => 33,
    26984 => 33,
    26985 => 33,
    26986 => 33,
    26987 => 33,
    26988 => 33,
    26989 => 33,
    26990 => 33,
    26991 => 33,
    26992 => 33,
    26993 => 33,
    26994 => 33,
    26995 => 33,
    26996 => 33,
    26997 => 33,
    26998 => 33,
    26999 => 33,
    27000 => 33,
    27001 => 33,
    27002 => 33,
    27003 => 33,
    27004 => 33,
    27005 => 33,
    27006 => 33,
    27007 => 33,
    27008 => 33,
    27009 => 33,
    27010 => 33,
    27011 => 33,
    27012 => 33,
    27013 => 33,
    27014 => 33,
    27015 => 33,
    27016 => 33,
    27017 => 33,
    27018 => 33,
    27019 => 33,
    27020 => 33,
    27021 => 33,
    27022 => 33,
    27023 => 33,
    27024 => 33,
    27025 => 33,
    27026 => 33,
    27027 => 33,
    27028 => 33,
    27029 => 33,
    27030 => 33,
    27031 => 33,
    27032 => 33,
    27033 => 33,
    27034 => 33,
    27035 => 33,
    27036 => 33,
    27037 => 33,
    27038 => 33,
    27039 => 33,
    27040 => 33,
    27041 => 33,
    27042 => 33,
    27043 => 33,
    27044 => 33,
    27045 => 33,
    27046 => 33,
    27047 => 33,
    27048 => 33,
    27049 => 33,
    27050 => 33,
    27051 => 33,
    27052 => 33,
    27053 => 33,
    27054 => 33,
    27055 => 33,
    27056 => 33,
    27057 => 33,
    27058 => 33,
    27059 => 33,
    27060 => 33,
    27061 => 33,
    27062 => 33,
    27063 => 33,
    27064 => 33,
    27065 => 33,
    27066 => 33,
    27067 => 33,
    27068 => 33,
    27069 => 33,
    27070 => 33,
    27071 => 33,
    27072 => 33,
    27073 => 33,
    27074 => 33,
    27075 => 33,
    27076 => 33,
    27077 => 33,
    27078 => 33,
    27079 => 33,
    27080 => 33,
    27081 => 33,
    27082 => 33,
    27083 => 33,
    27084 => 33,
    27085 => 33,
    27086 => 33,
    27087 => 33,
    27088 => 33,
    27089 => 33,
    27090 => 33,
    27091 => 33,
    27092 => 33,
    27093 => 33,
    27094 => 33,
    27095 => 33,
    27096 => 33,
    27097 => 33,
    27098 => 33,
    27099 => 33,
    27100 => 33,
    27101 => 33,
    27102 => 33,
    27103 => 33,
    27104 => 33,
    27105 => 33,
    27106 => 33,
    27107 => 33,
    27108 => 33,
    27109 => 33,
    27110 => 33,
    27111 => 33,
    27112 => 33,
    27113 => 33,
    27114 => 33,
    27115 => 32,
    27116 => 32,
    27117 => 32,
    27118 => 32,
    27119 => 32,
    27120 => 32,
    27121 => 32,
    27122 => 32,
    27123 => 32,
    27124 => 32,
    27125 => 32,
    27126 => 32,
    27127 => 32,
    27128 => 32,
    27129 => 32,
    27130 => 32,
    27131 => 32,
    27132 => 32,
    27133 => 32,
    27134 => 32,
    27135 => 32,
    27136 => 32,
    27137 => 32,
    27138 => 32,
    27139 => 32,
    27140 => 32,
    27141 => 32,
    27142 => 32,
    27143 => 32,
    27144 => 32,
    27145 => 32,
    27146 => 32,
    27147 => 32,
    27148 => 32,
    27149 => 32,
    27150 => 32,
    27151 => 32,
    27152 => 32,
    27153 => 32,
    27154 => 32,
    27155 => 32,
    27156 => 32,
    27157 => 32,
    27158 => 32,
    27159 => 32,
    27160 => 32,
    27161 => 32,
    27162 => 32,
    27163 => 32,
    27164 => 32,
    27165 => 32,
    27166 => 32,
    27167 => 32,
    27168 => 32,
    27169 => 32,
    27170 => 32,
    27171 => 32,
    27172 => 32,
    27173 => 32,
    27174 => 32,
    27175 => 32,
    27176 => 32,
    27177 => 32,
    27178 => 32,
    27179 => 32,
    27180 => 32,
    27181 => 32,
    27182 => 32,
    27183 => 32,
    27184 => 32,
    27185 => 32,
    27186 => 32,
    27187 => 32,
    27188 => 32,
    27189 => 32,
    27190 => 32,
    27191 => 32,
    27192 => 32,
    27193 => 32,
    27194 => 32,
    27195 => 32,
    27196 => 32,
    27197 => 32,
    27198 => 32,
    27199 => 32,
    27200 => 32,
    27201 => 32,
    27202 => 32,
    27203 => 32,
    27204 => 32,
    27205 => 32,
    27206 => 32,
    27207 => 32,
    27208 => 32,
    27209 => 32,
    27210 => 32,
    27211 => 32,
    27212 => 32,
    27213 => 32,
    27214 => 32,
    27215 => 32,
    27216 => 32,
    27217 => 32,
    27218 => 32,
    27219 => 32,
    27220 => 32,
    27221 => 32,
    27222 => 32,
    27223 => 32,
    27224 => 32,
    27225 => 32,
    27226 => 32,
    27227 => 32,
    27228 => 32,
    27229 => 32,
    27230 => 32,
    27231 => 32,
    27232 => 32,
    27233 => 32,
    27234 => 32,
    27235 => 32,
    27236 => 32,
    27237 => 32,
    27238 => 32,
    27239 => 32,
    27240 => 32,
    27241 => 32,
    27242 => 32,
    27243 => 32,
    27244 => 32,
    27245 => 32,
    27246 => 32,
    27247 => 32,
    27248 => 32,
    27249 => 32,
    27250 => 32,
    27251 => 32,
    27252 => 32,
    27253 => 32,
    27254 => 32,
    27255 => 32,
    27256 => 32,
    27257 => 32,
    27258 => 32,
    27259 => 32,
    27260 => 32,
    27261 => 32,
    27262 => 32,
    27263 => 32,
    27264 => 32,
    27265 => 32,
    27266 => 32,
    27267 => 32,
    27268 => 32,
    27269 => 32,
    27270 => 32,
    27271 => 32,
    27272 => 32,
    27273 => 32,
    27274 => 32,
    27275 => 32,
    27276 => 32,
    27277 => 32,
    27278 => 32,
    27279 => 32,
    27280 => 32,
    27281 => 32,
    27282 => 32,
    27283 => 32,
    27284 => 32,
    27285 => 32,
    27286 => 32,
    27287 => 32,
    27288 => 32,
    27289 => 32,
    27290 => 32,
    27291 => 32,
    27292 => 32,
    27293 => 32,
    27294 => 32,
    27295 => 32,
    27296 => 32,
    27297 => 32,
    27298 => 32,
    27299 => 32,
    27300 => 32,
    27301 => 32,
    27302 => 32,
    27303 => 32,
    27304 => 32,
    27305 => 32,
    27306 => 32,
    27307 => 31,
    27308 => 31,
    27309 => 31,
    27310 => 31,
    27311 => 31,
    27312 => 31,
    27313 => 31,
    27314 => 31,
    27315 => 31,
    27316 => 31,
    27317 => 31,
    27318 => 31,
    27319 => 31,
    27320 => 31,
    27321 => 31,
    27322 => 31,
    27323 => 31,
    27324 => 31,
    27325 => 31,
    27326 => 31,
    27327 => 31,
    27328 => 31,
    27329 => 31,
    27330 => 31,
    27331 => 31,
    27332 => 31,
    27333 => 31,
    27334 => 31,
    27335 => 31,
    27336 => 31,
    27337 => 31,
    27338 => 31,
    27339 => 31,
    27340 => 31,
    27341 => 31,
    27342 => 31,
    27343 => 31,
    27344 => 31,
    27345 => 31,
    27346 => 31,
    27347 => 31,
    27348 => 31,
    27349 => 31,
    27350 => 31,
    27351 => 31,
    27352 => 31,
    27353 => 31,
    27354 => 31,
    27355 => 31,
    27356 => 31,
    27357 => 31,
    27358 => 31,
    27359 => 31,
    27360 => 31,
    27361 => 31,
    27362 => 31,
    27363 => 31,
    27364 => 31,
    27365 => 31,
    27366 => 31,
    27367 => 31,
    27368 => 31,
    27369 => 31,
    27370 => 31,
    27371 => 31,
    27372 => 31,
    27373 => 31,
    27374 => 31,
    27375 => 31,
    27376 => 31,
    27377 => 31,
    27378 => 31,
    27379 => 31,
    27380 => 31,
    27381 => 31,
    27382 => 31,
    27383 => 31,
    27384 => 31,
    27385 => 31,
    27386 => 31,
    27387 => 31,
    27388 => 31,
    27389 => 31,
    27390 => 31,
    27391 => 31,
    27392 => 31,
    27393 => 31,
    27394 => 31,
    27395 => 31,
    27396 => 31,
    27397 => 31,
    27398 => 31,
    27399 => 31,
    27400 => 31,
    27401 => 31,
    27402 => 31,
    27403 => 31,
    27404 => 31,
    27405 => 31,
    27406 => 31,
    27407 => 31,
    27408 => 31,
    27409 => 31,
    27410 => 31,
    27411 => 31,
    27412 => 31,
    27413 => 31,
    27414 => 31,
    27415 => 31,
    27416 => 31,
    27417 => 31,
    27418 => 31,
    27419 => 31,
    27420 => 31,
    27421 => 31,
    27422 => 31,
    27423 => 31,
    27424 => 31,
    27425 => 31,
    27426 => 31,
    27427 => 31,
    27428 => 31,
    27429 => 31,
    27430 => 31,
    27431 => 31,
    27432 => 31,
    27433 => 31,
    27434 => 31,
    27435 => 31,
    27436 => 31,
    27437 => 31,
    27438 => 31,
    27439 => 31,
    27440 => 31,
    27441 => 31,
    27442 => 31,
    27443 => 31,
    27444 => 31,
    27445 => 31,
    27446 => 31,
    27447 => 31,
    27448 => 31,
    27449 => 31,
    27450 => 31,
    27451 => 31,
    27452 => 31,
    27453 => 31,
    27454 => 31,
    27455 => 31,
    27456 => 31,
    27457 => 31,
    27458 => 31,
    27459 => 31,
    27460 => 31,
    27461 => 31,
    27462 => 31,
    27463 => 31,
    27464 => 31,
    27465 => 31,
    27466 => 31,
    27467 => 31,
    27468 => 31,
    27469 => 31,
    27470 => 31,
    27471 => 31,
    27472 => 31,
    27473 => 31,
    27474 => 31,
    27475 => 31,
    27476 => 31,
    27477 => 31,
    27478 => 31,
    27479 => 31,
    27480 => 31,
    27481 => 31,
    27482 => 31,
    27483 => 31,
    27484 => 31,
    27485 => 31,
    27486 => 31,
    27487 => 31,
    27488 => 31,
    27489 => 31,
    27490 => 31,
    27491 => 31,
    27492 => 31,
    27493 => 31,
    27494 => 31,
    27495 => 31,
    27496 => 31,
    27497 => 30,
    27498 => 30,
    27499 => 30,
    27500 => 30,
    27501 => 30,
    27502 => 30,
    27503 => 30,
    27504 => 30,
    27505 => 30,
    27506 => 30,
    27507 => 30,
    27508 => 30,
    27509 => 30,
    27510 => 30,
    27511 => 30,
    27512 => 30,
    27513 => 30,
    27514 => 30,
    27515 => 30,
    27516 => 30,
    27517 => 30,
    27518 => 30,
    27519 => 30,
    27520 => 30,
    27521 => 30,
    27522 => 30,
    27523 => 30,
    27524 => 30,
    27525 => 30,
    27526 => 30,
    27527 => 30,
    27528 => 30,
    27529 => 30,
    27530 => 30,
    27531 => 30,
    27532 => 30,
    27533 => 30,
    27534 => 30,
    27535 => 30,
    27536 => 30,
    27537 => 30,
    27538 => 30,
    27539 => 30,
    27540 => 30,
    27541 => 30,
    27542 => 30,
    27543 => 30,
    27544 => 30,
    27545 => 30,
    27546 => 30,
    27547 => 30,
    27548 => 30,
    27549 => 30,
    27550 => 30,
    27551 => 30,
    27552 => 30,
    27553 => 30,
    27554 => 30,
    27555 => 30,
    27556 => 30,
    27557 => 30,
    27558 => 30,
    27559 => 30,
    27560 => 30,
    27561 => 30,
    27562 => 30,
    27563 => 30,
    27564 => 30,
    27565 => 30,
    27566 => 30,
    27567 => 30,
    27568 => 30,
    27569 => 30,
    27570 => 30,
    27571 => 30,
    27572 => 30,
    27573 => 30,
    27574 => 30,
    27575 => 30,
    27576 => 30,
    27577 => 30,
    27578 => 30,
    27579 => 30,
    27580 => 30,
    27581 => 30,
    27582 => 30,
    27583 => 30,
    27584 => 30,
    27585 => 30,
    27586 => 30,
    27587 => 30,
    27588 => 30,
    27589 => 30,
    27590 => 30,
    27591 => 30,
    27592 => 30,
    27593 => 30,
    27594 => 30,
    27595 => 30,
    27596 => 30,
    27597 => 30,
    27598 => 30,
    27599 => 30,
    27600 => 30,
    27601 => 30,
    27602 => 30,
    27603 => 30,
    27604 => 30,
    27605 => 30,
    27606 => 30,
    27607 => 30,
    27608 => 30,
    27609 => 30,
    27610 => 30,
    27611 => 30,
    27612 => 30,
    27613 => 30,
    27614 => 30,
    27615 => 30,
    27616 => 30,
    27617 => 30,
    27618 => 30,
    27619 => 30,
    27620 => 30,
    27621 => 30,
    27622 => 30,
    27623 => 30,
    27624 => 30,
    27625 => 30,
    27626 => 30,
    27627 => 30,
    27628 => 30,
    27629 => 30,
    27630 => 30,
    27631 => 30,
    27632 => 30,
    27633 => 30,
    27634 => 30,
    27635 => 30,
    27636 => 30,
    27637 => 30,
    27638 => 30,
    27639 => 30,
    27640 => 30,
    27641 => 30,
    27642 => 30,
    27643 => 30,
    27644 => 30,
    27645 => 30,
    27646 => 30,
    27647 => 30,
    27648 => 30,
    27649 => 30,
    27650 => 30,
    27651 => 30,
    27652 => 30,
    27653 => 30,
    27654 => 30,
    27655 => 30,
    27656 => 30,
    27657 => 30,
    27658 => 30,
    27659 => 30,
    27660 => 30,
    27661 => 30,
    27662 => 30,
    27663 => 30,
    27664 => 30,
    27665 => 30,
    27666 => 30,
    27667 => 30,
    27668 => 30,
    27669 => 30,
    27670 => 30,
    27671 => 30,
    27672 => 30,
    27673 => 30,
    27674 => 30,
    27675 => 30,
    27676 => 30,
    27677 => 30,
    27678 => 30,
    27679 => 30,
    27680 => 30,
    27681 => 30,
    27682 => 30,
    27683 => 30,
    27684 => 30,
    27685 => 30,
    27686 => 29,
    27687 => 29,
    27688 => 29,
    27689 => 29,
    27690 => 29,
    27691 => 29,
    27692 => 29,
    27693 => 29,
    27694 => 29,
    27695 => 29,
    27696 => 29,
    27697 => 29,
    27698 => 29,
    27699 => 29,
    27700 => 29,
    27701 => 29,
    27702 => 29,
    27703 => 29,
    27704 => 29,
    27705 => 29,
    27706 => 29,
    27707 => 29,
    27708 => 29,
    27709 => 29,
    27710 => 29,
    27711 => 29,
    27712 => 29,
    27713 => 29,
    27714 => 29,
    27715 => 29,
    27716 => 29,
    27717 => 29,
    27718 => 29,
    27719 => 29,
    27720 => 29,
    27721 => 29,
    27722 => 29,
    27723 => 29,
    27724 => 29,
    27725 => 29,
    27726 => 29,
    27727 => 29,
    27728 => 29,
    27729 => 29,
    27730 => 29,
    27731 => 29,
    27732 => 29,
    27733 => 29,
    27734 => 29,
    27735 => 29,
    27736 => 29,
    27737 => 29,
    27738 => 29,
    27739 => 29,
    27740 => 29,
    27741 => 29,
    27742 => 29,
    27743 => 29,
    27744 => 29,
    27745 => 29,
    27746 => 29,
    27747 => 29,
    27748 => 29,
    27749 => 29,
    27750 => 29,
    27751 => 29,
    27752 => 29,
    27753 => 29,
    27754 => 29,
    27755 => 29,
    27756 => 29,
    27757 => 29,
    27758 => 29,
    27759 => 29,
    27760 => 29,
    27761 => 29,
    27762 => 29,
    27763 => 29,
    27764 => 29,
    27765 => 29,
    27766 => 29,
    27767 => 29,
    27768 => 29,
    27769 => 29,
    27770 => 29,
    27771 => 29,
    27772 => 29,
    27773 => 29,
    27774 => 29,
    27775 => 29,
    27776 => 29,
    27777 => 29,
    27778 => 29,
    27779 => 29,
    27780 => 29,
    27781 => 29,
    27782 => 29,
    27783 => 29,
    27784 => 29,
    27785 => 29,
    27786 => 29,
    27787 => 29,
    27788 => 29,
    27789 => 29,
    27790 => 29,
    27791 => 29,
    27792 => 29,
    27793 => 29,
    27794 => 29,
    27795 => 29,
    27796 => 29,
    27797 => 29,
    27798 => 29,
    27799 => 29,
    27800 => 29,
    27801 => 29,
    27802 => 29,
    27803 => 29,
    27804 => 29,
    27805 => 29,
    27806 => 29,
    27807 => 29,
    27808 => 29,
    27809 => 29,
    27810 => 29,
    27811 => 29,
    27812 => 29,
    27813 => 29,
    27814 => 29,
    27815 => 29,
    27816 => 29,
    27817 => 29,
    27818 => 29,
    27819 => 29,
    27820 => 29,
    27821 => 29,
    27822 => 29,
    27823 => 29,
    27824 => 29,
    27825 => 29,
    27826 => 29,
    27827 => 29,
    27828 => 29,
    27829 => 29,
    27830 => 29,
    27831 => 29,
    27832 => 29,
    27833 => 29,
    27834 => 29,
    27835 => 29,
    27836 => 29,
    27837 => 29,
    27838 => 29,
    27839 => 29,
    27840 => 29,
    27841 => 29,
    27842 => 29,
    27843 => 29,
    27844 => 29,
    27845 => 29,
    27846 => 29,
    27847 => 29,
    27848 => 29,
    27849 => 29,
    27850 => 29,
    27851 => 29,
    27852 => 29,
    27853 => 29,
    27854 => 29,
    27855 => 29,
    27856 => 29,
    27857 => 29,
    27858 => 29,
    27859 => 29,
    27860 => 29,
    27861 => 29,
    27862 => 29,
    27863 => 29,
    27864 => 29,
    27865 => 29,
    27866 => 29,
    27867 => 29,
    27868 => 29,
    27869 => 29,
    27870 => 29,
    27871 => 29,
    27872 => 28,
    27873 => 28,
    27874 => 28,
    27875 => 28,
    27876 => 28,
    27877 => 28,
    27878 => 28,
    27879 => 28,
    27880 => 28,
    27881 => 28,
    27882 => 28,
    27883 => 28,
    27884 => 28,
    27885 => 28,
    27886 => 28,
    27887 => 28,
    27888 => 28,
    27889 => 28,
    27890 => 28,
    27891 => 28,
    27892 => 28,
    27893 => 28,
    27894 => 28,
    27895 => 28,
    27896 => 28,
    27897 => 28,
    27898 => 28,
    27899 => 28,
    27900 => 28,
    27901 => 28,
    27902 => 28,
    27903 => 28,
    27904 => 28,
    27905 => 28,
    27906 => 28,
    27907 => 28,
    27908 => 28,
    27909 => 28,
    27910 => 28,
    27911 => 28,
    27912 => 28,
    27913 => 28,
    27914 => 28,
    27915 => 28,
    27916 => 28,
    27917 => 28,
    27918 => 28,
    27919 => 28,
    27920 => 28,
    27921 => 28,
    27922 => 28,
    27923 => 28,
    27924 => 28,
    27925 => 28,
    27926 => 28,
    27927 => 28,
    27928 => 28,
    27929 => 28,
    27930 => 28,
    27931 => 28,
    27932 => 28,
    27933 => 28,
    27934 => 28,
    27935 => 28,
    27936 => 28,
    27937 => 28,
    27938 => 28,
    27939 => 28,
    27940 => 28,
    27941 => 28,
    27942 => 28,
    27943 => 28,
    27944 => 28,
    27945 => 28,
    27946 => 28,
    27947 => 28,
    27948 => 28,
    27949 => 28,
    27950 => 28,
    27951 => 28,
    27952 => 28,
    27953 => 28,
    27954 => 28,
    27955 => 28,
    27956 => 28,
    27957 => 28,
    27958 => 28,
    27959 => 28,
    27960 => 28,
    27961 => 28,
    27962 => 28,
    27963 => 28,
    27964 => 28,
    27965 => 28,
    27966 => 28,
    27967 => 28,
    27968 => 28,
    27969 => 28,
    27970 => 28,
    27971 => 28,
    27972 => 28,
    27973 => 28,
    27974 => 28,
    27975 => 28,
    27976 => 28,
    27977 => 28,
    27978 => 28,
    27979 => 28,
    27980 => 28,
    27981 => 28,
    27982 => 28,
    27983 => 28,
    27984 => 28,
    27985 => 28,
    27986 => 28,
    27987 => 28,
    27988 => 28,
    27989 => 28,
    27990 => 28,
    27991 => 28,
    27992 => 28,
    27993 => 28,
    27994 => 28,
    27995 => 28,
    27996 => 28,
    27997 => 28,
    27998 => 28,
    27999 => 28,
    28000 => 28,
    28001 => 28,
    28002 => 28,
    28003 => 28,
    28004 => 28,
    28005 => 28,
    28006 => 28,
    28007 => 28,
    28008 => 28,
    28009 => 28,
    28010 => 28,
    28011 => 28,
    28012 => 28,
    28013 => 28,
    28014 => 28,
    28015 => 28,
    28016 => 28,
    28017 => 28,
    28018 => 28,
    28019 => 28,
    28020 => 28,
    28021 => 28,
    28022 => 28,
    28023 => 28,
    28024 => 28,
    28025 => 28,
    28026 => 28,
    28027 => 28,
    28028 => 28,
    28029 => 28,
    28030 => 28,
    28031 => 28,
    28032 => 28,
    28033 => 28,
    28034 => 28,
    28035 => 28,
    28036 => 28,
    28037 => 28,
    28038 => 28,
    28039 => 28,
    28040 => 28,
    28041 => 28,
    28042 => 28,
    28043 => 28,
    28044 => 28,
    28045 => 28,
    28046 => 28,
    28047 => 28,
    28048 => 28,
    28049 => 28,
    28050 => 28,
    28051 => 28,
    28052 => 28,
    28053 => 28,
    28054 => 28,
    28055 => 28,
    28056 => 28,
    28057 => 27,
    28058 => 27,
    28059 => 27,
    28060 => 27,
    28061 => 27,
    28062 => 27,
    28063 => 27,
    28064 => 27,
    28065 => 27,
    28066 => 27,
    28067 => 27,
    28068 => 27,
    28069 => 27,
    28070 => 27,
    28071 => 27,
    28072 => 27,
    28073 => 27,
    28074 => 27,
    28075 => 27,
    28076 => 27,
    28077 => 27,
    28078 => 27,
    28079 => 27,
    28080 => 27,
    28081 => 27,
    28082 => 27,
    28083 => 27,
    28084 => 27,
    28085 => 27,
    28086 => 27,
    28087 => 27,
    28088 => 27,
    28089 => 27,
    28090 => 27,
    28091 => 27,
    28092 => 27,
    28093 => 27,
    28094 => 27,
    28095 => 27,
    28096 => 27,
    28097 => 27,
    28098 => 27,
    28099 => 27,
    28100 => 27,
    28101 => 27,
    28102 => 27,
    28103 => 27,
    28104 => 27,
    28105 => 27,
    28106 => 27,
    28107 => 27,
    28108 => 27,
    28109 => 27,
    28110 => 27,
    28111 => 27,
    28112 => 27,
    28113 => 27,
    28114 => 27,
    28115 => 27,
    28116 => 27,
    28117 => 27,
    28118 => 27,
    28119 => 27,
    28120 => 27,
    28121 => 27,
    28122 => 27,
    28123 => 27,
    28124 => 27,
    28125 => 27,
    28126 => 27,
    28127 => 27,
    28128 => 27,
    28129 => 27,
    28130 => 27,
    28131 => 27,
    28132 => 27,
    28133 => 27,
    28134 => 27,
    28135 => 27,
    28136 => 27,
    28137 => 27,
    28138 => 27,
    28139 => 27,
    28140 => 27,
    28141 => 27,
    28142 => 27,
    28143 => 27,
    28144 => 27,
    28145 => 27,
    28146 => 27,
    28147 => 27,
    28148 => 27,
    28149 => 27,
    28150 => 27,
    28151 => 27,
    28152 => 27,
    28153 => 27,
    28154 => 27,
    28155 => 27,
    28156 => 27,
    28157 => 27,
    28158 => 27,
    28159 => 27,
    28160 => 27,
    28161 => 27,
    28162 => 27,
    28163 => 27,
    28164 => 27,
    28165 => 27,
    28166 => 27,
    28167 => 27,
    28168 => 27,
    28169 => 27,
    28170 => 27,
    28171 => 27,
    28172 => 27,
    28173 => 27,
    28174 => 27,
    28175 => 27,
    28176 => 27,
    28177 => 27,
    28178 => 27,
    28179 => 27,
    28180 => 27,
    28181 => 27,
    28182 => 27,
    28183 => 27,
    28184 => 27,
    28185 => 27,
    28186 => 27,
    28187 => 27,
    28188 => 27,
    28189 => 27,
    28190 => 27,
    28191 => 27,
    28192 => 27,
    28193 => 27,
    28194 => 27,
    28195 => 27,
    28196 => 27,
    28197 => 27,
    28198 => 27,
    28199 => 27,
    28200 => 27,
    28201 => 27,
    28202 => 27,
    28203 => 27,
    28204 => 27,
    28205 => 27,
    28206 => 27,
    28207 => 27,
    28208 => 27,
    28209 => 27,
    28210 => 27,
    28211 => 27,
    28212 => 27,
    28213 => 27,
    28214 => 27,
    28215 => 27,
    28216 => 27,
    28217 => 27,
    28218 => 27,
    28219 => 27,
    28220 => 27,
    28221 => 27,
    28222 => 27,
    28223 => 27,
    28224 => 27,
    28225 => 27,
    28226 => 27,
    28227 => 27,
    28228 => 27,
    28229 => 27,
    28230 => 27,
    28231 => 27,
    28232 => 27,
    28233 => 27,
    28234 => 27,
    28235 => 27,
    28236 => 27,
    28237 => 27,
    28238 => 27,
    28239 => 27,
    28240 => 26,
    28241 => 26,
    28242 => 26,
    28243 => 26,
    28244 => 26,
    28245 => 26,
    28246 => 26,
    28247 => 26,
    28248 => 26,
    28249 => 26,
    28250 => 26,
    28251 => 26,
    28252 => 26,
    28253 => 26,
    28254 => 26,
    28255 => 26,
    28256 => 26,
    28257 => 26,
    28258 => 26,
    28259 => 26,
    28260 => 26,
    28261 => 26,
    28262 => 26,
    28263 => 26,
    28264 => 26,
    28265 => 26,
    28266 => 26,
    28267 => 26,
    28268 => 26,
    28269 => 26,
    28270 => 26,
    28271 => 26,
    28272 => 26,
    28273 => 26,
    28274 => 26,
    28275 => 26,
    28276 => 26,
    28277 => 26,
    28278 => 26,
    28279 => 26,
    28280 => 26,
    28281 => 26,
    28282 => 26,
    28283 => 26,
    28284 => 26,
    28285 => 26,
    28286 => 26,
    28287 => 26,
    28288 => 26,
    28289 => 26,
    28290 => 26,
    28291 => 26,
    28292 => 26,
    28293 => 26,
    28294 => 26,
    28295 => 26,
    28296 => 26,
    28297 => 26,
    28298 => 26,
    28299 => 26,
    28300 => 26,
    28301 => 26,
    28302 => 26,
    28303 => 26,
    28304 => 26,
    28305 => 26,
    28306 => 26,
    28307 => 26,
    28308 => 26,
    28309 => 26,
    28310 => 26,
    28311 => 26,
    28312 => 26,
    28313 => 26,
    28314 => 26,
    28315 => 26,
    28316 => 26,
    28317 => 26,
    28318 => 26,
    28319 => 26,
    28320 => 26,
    28321 => 26,
    28322 => 26,
    28323 => 26,
    28324 => 26,
    28325 => 26,
    28326 => 26,
    28327 => 26,
    28328 => 26,
    28329 => 26,
    28330 => 26,
    28331 => 26,
    28332 => 26,
    28333 => 26,
    28334 => 26,
    28335 => 26,
    28336 => 26,
    28337 => 26,
    28338 => 26,
    28339 => 26,
    28340 => 26,
    28341 => 26,
    28342 => 26,
    28343 => 26,
    28344 => 26,
    28345 => 26,
    28346 => 26,
    28347 => 26,
    28348 => 26,
    28349 => 26,
    28350 => 26,
    28351 => 26,
    28352 => 26,
    28353 => 26,
    28354 => 26,
    28355 => 26,
    28356 => 26,
    28357 => 26,
    28358 => 26,
    28359 => 26,
    28360 => 26,
    28361 => 26,
    28362 => 26,
    28363 => 26,
    28364 => 26,
    28365 => 26,
    28366 => 26,
    28367 => 26,
    28368 => 26,
    28369 => 26,
    28370 => 26,
    28371 => 26,
    28372 => 26,
    28373 => 26,
    28374 => 26,
    28375 => 26,
    28376 => 26,
    28377 => 26,
    28378 => 26,
    28379 => 26,
    28380 => 26,
    28381 => 26,
    28382 => 26,
    28383 => 26,
    28384 => 26,
    28385 => 26,
    28386 => 26,
    28387 => 26,
    28388 => 26,
    28389 => 26,
    28390 => 26,
    28391 => 26,
    28392 => 26,
    28393 => 26,
    28394 => 26,
    28395 => 26,
    28396 => 26,
    28397 => 26,
    28398 => 26,
    28399 => 26,
    28400 => 26,
    28401 => 26,
    28402 => 26,
    28403 => 26,
    28404 => 26,
    28405 => 26,
    28406 => 26,
    28407 => 26,
    28408 => 26,
    28409 => 26,
    28410 => 26,
    28411 => 26,
    28412 => 26,
    28413 => 26,
    28414 => 26,
    28415 => 26,
    28416 => 26,
    28417 => 26,
    28418 => 26,
    28419 => 26,
    28420 => 26,
    28421 => 26,
    28422 => 25,
    28423 => 25,
    28424 => 25,
    28425 => 25,
    28426 => 25,
    28427 => 25,
    28428 => 25,
    28429 => 25,
    28430 => 25,
    28431 => 25,
    28432 => 25,
    28433 => 25,
    28434 => 25,
    28435 => 25,
    28436 => 25,
    28437 => 25,
    28438 => 25,
    28439 => 25,
    28440 => 25,
    28441 => 25,
    28442 => 25,
    28443 => 25,
    28444 => 25,
    28445 => 25,
    28446 => 25,
    28447 => 25,
    28448 => 25,
    28449 => 25,
    28450 => 25,
    28451 => 25,
    28452 => 25,
    28453 => 25,
    28454 => 25,
    28455 => 25,
    28456 => 25,
    28457 => 25,
    28458 => 25,
    28459 => 25,
    28460 => 25,
    28461 => 25,
    28462 => 25,
    28463 => 25,
    28464 => 25,
    28465 => 25,
    28466 => 25,
    28467 => 25,
    28468 => 25,
    28469 => 25,
    28470 => 25,
    28471 => 25,
    28472 => 25,
    28473 => 25,
    28474 => 25,
    28475 => 25,
    28476 => 25,
    28477 => 25,
    28478 => 25,
    28479 => 25,
    28480 => 25,
    28481 => 25,
    28482 => 25,
    28483 => 25,
    28484 => 25,
    28485 => 25,
    28486 => 25,
    28487 => 25,
    28488 => 25,
    28489 => 25,
    28490 => 25,
    28491 => 25,
    28492 => 25,
    28493 => 25,
    28494 => 25,
    28495 => 25,
    28496 => 25,
    28497 => 25,
    28498 => 25,
    28499 => 25,
    28500 => 25,
    28501 => 25,
    28502 => 25,
    28503 => 25,
    28504 => 25,
    28505 => 25,
    28506 => 25,
    28507 => 25,
    28508 => 25,
    28509 => 25,
    28510 => 25,
    28511 => 25,
    28512 => 25,
    28513 => 25,
    28514 => 25,
    28515 => 25,
    28516 => 25,
    28517 => 25,
    28518 => 25,
    28519 => 25,
    28520 => 25,
    28521 => 25,
    28522 => 25,
    28523 => 25,
    28524 => 25,
    28525 => 25,
    28526 => 25,
    28527 => 25,
    28528 => 25,
    28529 => 25,
    28530 => 25,
    28531 => 25,
    28532 => 25,
    28533 => 25,
    28534 => 25,
    28535 => 25,
    28536 => 25,
    28537 => 25,
    28538 => 25,
    28539 => 25,
    28540 => 25,
    28541 => 25,
    28542 => 25,
    28543 => 25,
    28544 => 25,
    28545 => 25,
    28546 => 25,
    28547 => 25,
    28548 => 25,
    28549 => 25,
    28550 => 25,
    28551 => 25,
    28552 => 25,
    28553 => 25,
    28554 => 25,
    28555 => 25,
    28556 => 25,
    28557 => 25,
    28558 => 25,
    28559 => 25,
    28560 => 25,
    28561 => 25,
    28562 => 25,
    28563 => 25,
    28564 => 25,
    28565 => 25,
    28566 => 25,
    28567 => 25,
    28568 => 25,
    28569 => 25,
    28570 => 25,
    28571 => 25,
    28572 => 25,
    28573 => 25,
    28574 => 25,
    28575 => 25,
    28576 => 25,
    28577 => 25,
    28578 => 25,
    28579 => 25,
    28580 => 25,
    28581 => 25,
    28582 => 25,
    28583 => 25,
    28584 => 25,
    28585 => 25,
    28586 => 25,
    28587 => 25,
    28588 => 25,
    28589 => 25,
    28590 => 25,
    28591 => 25,
    28592 => 25,
    28593 => 25,
    28594 => 25,
    28595 => 25,
    28596 => 25,
    28597 => 25,
    28598 => 25,
    28599 => 25,
    28600 => 25,
    28601 => 25,
    28602 => 24,
    28603 => 24,
    28604 => 24,
    28605 => 24,
    28606 => 24,
    28607 => 24,
    28608 => 24,
    28609 => 24,
    28610 => 24,
    28611 => 24,
    28612 => 24,
    28613 => 24,
    28614 => 24,
    28615 => 24,
    28616 => 24,
    28617 => 24,
    28618 => 24,
    28619 => 24,
    28620 => 24,
    28621 => 24,
    28622 => 24,
    28623 => 24,
    28624 => 24,
    28625 => 24,
    28626 => 24,
    28627 => 24,
    28628 => 24,
    28629 => 24,
    28630 => 24,
    28631 => 24,
    28632 => 24,
    28633 => 24,
    28634 => 24,
    28635 => 24,
    28636 => 24,
    28637 => 24,
    28638 => 24,
    28639 => 24,
    28640 => 24,
    28641 => 24,
    28642 => 24,
    28643 => 24,
    28644 => 24,
    28645 => 24,
    28646 => 24,
    28647 => 24,
    28648 => 24,
    28649 => 24,
    28650 => 24,
    28651 => 24,
    28652 => 24,
    28653 => 24,
    28654 => 24,
    28655 => 24,
    28656 => 24,
    28657 => 24,
    28658 => 24,
    28659 => 24,
    28660 => 24,
    28661 => 24,
    28662 => 24,
    28663 => 24,
    28664 => 24,
    28665 => 24,
    28666 => 24,
    28667 => 24,
    28668 => 24,
    28669 => 24,
    28670 => 24,
    28671 => 24,
    28672 => 24,
    28673 => 24,
    28674 => 24,
    28675 => 24,
    28676 => 24,
    28677 => 24,
    28678 => 24,
    28679 => 24,
    28680 => 24,
    28681 => 24,
    28682 => 24,
    28683 => 24,
    28684 => 24,
    28685 => 24,
    28686 => 24,
    28687 => 24,
    28688 => 24,
    28689 => 24,
    28690 => 24,
    28691 => 24,
    28692 => 24,
    28693 => 24,
    28694 => 24,
    28695 => 24,
    28696 => 24,
    28697 => 24,
    28698 => 24,
    28699 => 24,
    28700 => 24,
    28701 => 24,
    28702 => 24,
    28703 => 24,
    28704 => 24,
    28705 => 24,
    28706 => 24,
    28707 => 24,
    28708 => 24,
    28709 => 24,
    28710 => 24,
    28711 => 24,
    28712 => 24,
    28713 => 24,
    28714 => 24,
    28715 => 24,
    28716 => 24,
    28717 => 24,
    28718 => 24,
    28719 => 24,
    28720 => 24,
    28721 => 24,
    28722 => 24,
    28723 => 24,
    28724 => 24,
    28725 => 24,
    28726 => 24,
    28727 => 24,
    28728 => 24,
    28729 => 24,
    28730 => 24,
    28731 => 24,
    28732 => 24,
    28733 => 24,
    28734 => 24,
    28735 => 24,
    28736 => 24,
    28737 => 24,
    28738 => 24,
    28739 => 24,
    28740 => 24,
    28741 => 24,
    28742 => 24,
    28743 => 24,
    28744 => 24,
    28745 => 24,
    28746 => 24,
    28747 => 24,
    28748 => 24,
    28749 => 24,
    28750 => 24,
    28751 => 24,
    28752 => 24,
    28753 => 24,
    28754 => 24,
    28755 => 24,
    28756 => 24,
    28757 => 24,
    28758 => 24,
    28759 => 24,
    28760 => 24,
    28761 => 24,
    28762 => 24,
    28763 => 24,
    28764 => 24,
    28765 => 24,
    28766 => 24,
    28767 => 24,
    28768 => 24,
    28769 => 24,
    28770 => 24,
    28771 => 24,
    28772 => 24,
    28773 => 24,
    28774 => 24,
    28775 => 24,
    28776 => 24,
    28777 => 24,
    28778 => 24,
    28779 => 24,
    28780 => 24,
    28781 => 23,
    28782 => 23,
    28783 => 23,
    28784 => 23,
    28785 => 23,
    28786 => 23,
    28787 => 23,
    28788 => 23,
    28789 => 23,
    28790 => 23,
    28791 => 23,
    28792 => 23,
    28793 => 23,
    28794 => 23,
    28795 => 23,
    28796 => 23,
    28797 => 23,
    28798 => 23,
    28799 => 23,
    28800 => 23,
    28801 => 23,
    28802 => 23,
    28803 => 23,
    28804 => 23,
    28805 => 23,
    28806 => 23,
    28807 => 23,
    28808 => 23,
    28809 => 23,
    28810 => 23,
    28811 => 23,
    28812 => 23,
    28813 => 23,
    28814 => 23,
    28815 => 23,
    28816 => 23,
    28817 => 23,
    28818 => 23,
    28819 => 23,
    28820 => 23,
    28821 => 23,
    28822 => 23,
    28823 => 23,
    28824 => 23,
    28825 => 23,
    28826 => 23,
    28827 => 23,
    28828 => 23,
    28829 => 23,
    28830 => 23,
    28831 => 23,
    28832 => 23,
    28833 => 23,
    28834 => 23,
    28835 => 23,
    28836 => 23,
    28837 => 23,
    28838 => 23,
    28839 => 23,
    28840 => 23,
    28841 => 23,
    28842 => 23,
    28843 => 23,
    28844 => 23,
    28845 => 23,
    28846 => 23,
    28847 => 23,
    28848 => 23,
    28849 => 23,
    28850 => 23,
    28851 => 23,
    28852 => 23,
    28853 => 23,
    28854 => 23,
    28855 => 23,
    28856 => 23,
    28857 => 23,
    28858 => 23,
    28859 => 23,
    28860 => 23,
    28861 => 23,
    28862 => 23,
    28863 => 23,
    28864 => 23,
    28865 => 23,
    28866 => 23,
    28867 => 23,
    28868 => 23,
    28869 => 23,
    28870 => 23,
    28871 => 23,
    28872 => 23,
    28873 => 23,
    28874 => 23,
    28875 => 23,
    28876 => 23,
    28877 => 23,
    28878 => 23,
    28879 => 23,
    28880 => 23,
    28881 => 23,
    28882 => 23,
    28883 => 23,
    28884 => 23,
    28885 => 23,
    28886 => 23,
    28887 => 23,
    28888 => 23,
    28889 => 23,
    28890 => 23,
    28891 => 23,
    28892 => 23,
    28893 => 23,
    28894 => 23,
    28895 => 23,
    28896 => 23,
    28897 => 23,
    28898 => 23,
    28899 => 23,
    28900 => 23,
    28901 => 23,
    28902 => 23,
    28903 => 23,
    28904 => 23,
    28905 => 23,
    28906 => 23,
    28907 => 23,
    28908 => 23,
    28909 => 23,
    28910 => 23,
    28911 => 23,
    28912 => 23,
    28913 => 23,
    28914 => 23,
    28915 => 23,
    28916 => 23,
    28917 => 23,
    28918 => 23,
    28919 => 23,
    28920 => 23,
    28921 => 23,
    28922 => 23,
    28923 => 23,
    28924 => 23,
    28925 => 23,
    28926 => 23,
    28927 => 23,
    28928 => 23,
    28929 => 23,
    28930 => 23,
    28931 => 23,
    28932 => 23,
    28933 => 23,
    28934 => 23,
    28935 => 23,
    28936 => 23,
    28937 => 23,
    28938 => 23,
    28939 => 23,
    28940 => 23,
    28941 => 23,
    28942 => 23,
    28943 => 23,
    28944 => 23,
    28945 => 23,
    28946 => 23,
    28947 => 23,
    28948 => 23,
    28949 => 23,
    28950 => 23,
    28951 => 23,
    28952 => 23,
    28953 => 23,
    28954 => 23,
    28955 => 23,
    28956 => 23,
    28957 => 23,
    28958 => 23,
    28959 => 22,
    28960 => 22,
    28961 => 22,
    28962 => 22,
    28963 => 22,
    28964 => 22,
    28965 => 22,
    28966 => 22,
    28967 => 22,
    28968 => 22,
    28969 => 22,
    28970 => 22,
    28971 => 22,
    28972 => 22,
    28973 => 22,
    28974 => 22,
    28975 => 22,
    28976 => 22,
    28977 => 22,
    28978 => 22,
    28979 => 22,
    28980 => 22,
    28981 => 22,
    28982 => 22,
    28983 => 22,
    28984 => 22,
    28985 => 22,
    28986 => 22,
    28987 => 22,
    28988 => 22,
    28989 => 22,
    28990 => 22,
    28991 => 22,
    28992 => 22,
    28993 => 22,
    28994 => 22,
    28995 => 22,
    28996 => 22,
    28997 => 22,
    28998 => 22,
    28999 => 22,
    29000 => 22,
    29001 => 22,
    29002 => 22,
    29003 => 22,
    29004 => 22,
    29005 => 22,
    29006 => 22,
    29007 => 22,
    29008 => 22,
    29009 => 22,
    29010 => 22,
    29011 => 22,
    29012 => 22,
    29013 => 22,
    29014 => 22,
    29015 => 22,
    29016 => 22,
    29017 => 22,
    29018 => 22,
    29019 => 22,
    29020 => 22,
    29021 => 22,
    29022 => 22,
    29023 => 22,
    29024 => 22,
    29025 => 22,
    29026 => 22,
    29027 => 22,
    29028 => 22,
    29029 => 22,
    29030 => 22,
    29031 => 22,
    29032 => 22,
    29033 => 22,
    29034 => 22,
    29035 => 22,
    29036 => 22,
    29037 => 22,
    29038 => 22,
    29039 => 22,
    29040 => 22,
    29041 => 22,
    29042 => 22,
    29043 => 22,
    29044 => 22,
    29045 => 22,
    29046 => 22,
    29047 => 22,
    29048 => 22,
    29049 => 22,
    29050 => 22,
    29051 => 22,
    29052 => 22,
    29053 => 22,
    29054 => 22,
    29055 => 22,
    29056 => 22,
    29057 => 22,
    29058 => 22,
    29059 => 22,
    29060 => 22,
    29061 => 22,
    29062 => 22,
    29063 => 22,
    29064 => 22,
    29065 => 22,
    29066 => 22,
    29067 => 22,
    29068 => 22,
    29069 => 22,
    29070 => 22,
    29071 => 22,
    29072 => 22,
    29073 => 22,
    29074 => 22,
    29075 => 22,
    29076 => 22,
    29077 => 22,
    29078 => 22,
    29079 => 22,
    29080 => 22,
    29081 => 22,
    29082 => 22,
    29083 => 22,
    29084 => 22,
    29085 => 22,
    29086 => 22,
    29087 => 22,
    29088 => 22,
    29089 => 22,
    29090 => 22,
    29091 => 22,
    29092 => 22,
    29093 => 22,
    29094 => 22,
    29095 => 22,
    29096 => 22,
    29097 => 22,
    29098 => 22,
    29099 => 22,
    29100 => 22,
    29101 => 22,
    29102 => 22,
    29103 => 22,
    29104 => 22,
    29105 => 22,
    29106 => 22,
    29107 => 22,
    29108 => 22,
    29109 => 22,
    29110 => 22,
    29111 => 22,
    29112 => 22,
    29113 => 22,
    29114 => 22,
    29115 => 22,
    29116 => 22,
    29117 => 22,
    29118 => 22,
    29119 => 22,
    29120 => 22,
    29121 => 22,
    29122 => 22,
    29123 => 22,
    29124 => 22,
    29125 => 22,
    29126 => 22,
    29127 => 22,
    29128 => 22,
    29129 => 22,
    29130 => 22,
    29131 => 22,
    29132 => 22,
    29133 => 22,
    29134 => 22,
    29135 => 22,
    29136 => 21,
    29137 => 21,
    29138 => 21,
    29139 => 21,
    29140 => 21,
    29141 => 21,
    29142 => 21,
    29143 => 21,
    29144 => 21,
    29145 => 21,
    29146 => 21,
    29147 => 21,
    29148 => 21,
    29149 => 21,
    29150 => 21,
    29151 => 21,
    29152 => 21,
    29153 => 21,
    29154 => 21,
    29155 => 21,
    29156 => 21,
    29157 => 21,
    29158 => 21,
    29159 => 21,
    29160 => 21,
    29161 => 21,
    29162 => 21,
    29163 => 21,
    29164 => 21,
    29165 => 21,
    29166 => 21,
    29167 => 21,
    29168 => 21,
    29169 => 21,
    29170 => 21,
    29171 => 21,
    29172 => 21,
    29173 => 21,
    29174 => 21,
    29175 => 21,
    29176 => 21,
    29177 => 21,
    29178 => 21,
    29179 => 21,
    29180 => 21,
    29181 => 21,
    29182 => 21,
    29183 => 21,
    29184 => 21,
    29185 => 21,
    29186 => 21,
    29187 => 21,
    29188 => 21,
    29189 => 21,
    29190 => 21,
    29191 => 21,
    29192 => 21,
    29193 => 21,
    29194 => 21,
    29195 => 21,
    29196 => 21,
    29197 => 21,
    29198 => 21,
    29199 => 21,
    29200 => 21,
    29201 => 21,
    29202 => 21,
    29203 => 21,
    29204 => 21,
    29205 => 21,
    29206 => 21,
    29207 => 21,
    29208 => 21,
    29209 => 21,
    29210 => 21,
    29211 => 21,
    29212 => 21,
    29213 => 21,
    29214 => 21,
    29215 => 21,
    29216 => 21,
    29217 => 21,
    29218 => 21,
    29219 => 21,
    29220 => 21,
    29221 => 21,
    29222 => 21,
    29223 => 21,
    29224 => 21,
    29225 => 21,
    29226 => 21,
    29227 => 21,
    29228 => 21,
    29229 => 21,
    29230 => 21,
    29231 => 21,
    29232 => 21,
    29233 => 21,
    29234 => 21,
    29235 => 21,
    29236 => 21,
    29237 => 21,
    29238 => 21,
    29239 => 21,
    29240 => 21,
    29241 => 21,
    29242 => 21,
    29243 => 21,
    29244 => 21,
    29245 => 21,
    29246 => 21,
    29247 => 21,
    29248 => 21,
    29249 => 21,
    29250 => 21,
    29251 => 21,
    29252 => 21,
    29253 => 21,
    29254 => 21,
    29255 => 21,
    29256 => 21,
    29257 => 21,
    29258 => 21,
    29259 => 21,
    29260 => 21,
    29261 => 21,
    29262 => 21,
    29263 => 21,
    29264 => 21,
    29265 => 21,
    29266 => 21,
    29267 => 21,
    29268 => 21,
    29269 => 21,
    29270 => 21,
    29271 => 21,
    29272 => 21,
    29273 => 21,
    29274 => 21,
    29275 => 21,
    29276 => 21,
    29277 => 21,
    29278 => 21,
    29279 => 21,
    29280 => 21,
    29281 => 21,
    29282 => 21,
    29283 => 21,
    29284 => 21,
    29285 => 21,
    29286 => 21,
    29287 => 21,
    29288 => 21,
    29289 => 21,
    29290 => 21,
    29291 => 21,
    29292 => 21,
    29293 => 21,
    29294 => 21,
    29295 => 21,
    29296 => 21,
    29297 => 21,
    29298 => 21,
    29299 => 21,
    29300 => 21,
    29301 => 21,
    29302 => 21,
    29303 => 21,
    29304 => 21,
    29305 => 21,
    29306 => 21,
    29307 => 21,
    29308 => 21,
    29309 => 21,
    29310 => 21,
    29311 => 21,
    29312 => 20,
    29313 => 20,
    29314 => 20,
    29315 => 20,
    29316 => 20,
    29317 => 20,
    29318 => 20,
    29319 => 20,
    29320 => 20,
    29321 => 20,
    29322 => 20,
    29323 => 20,
    29324 => 20,
    29325 => 20,
    29326 => 20,
    29327 => 20,
    29328 => 20,
    29329 => 20,
    29330 => 20,
    29331 => 20,
    29332 => 20,
    29333 => 20,
    29334 => 20,
    29335 => 20,
    29336 => 20,
    29337 => 20,
    29338 => 20,
    29339 => 20,
    29340 => 20,
    29341 => 20,
    29342 => 20,
    29343 => 20,
    29344 => 20,
    29345 => 20,
    29346 => 20,
    29347 => 20,
    29348 => 20,
    29349 => 20,
    29350 => 20,
    29351 => 20,
    29352 => 20,
    29353 => 20,
    29354 => 20,
    29355 => 20,
    29356 => 20,
    29357 => 20,
    29358 => 20,
    29359 => 20,
    29360 => 20,
    29361 => 20,
    29362 => 20,
    29363 => 20,
    29364 => 20,
    29365 => 20,
    29366 => 20,
    29367 => 20,
    29368 => 20,
    29369 => 20,
    29370 => 20,
    29371 => 20,
    29372 => 20,
    29373 => 20,
    29374 => 20,
    29375 => 20,
    29376 => 20,
    29377 => 20,
    29378 => 20,
    29379 => 20,
    29380 => 20,
    29381 => 20,
    29382 => 20,
    29383 => 20,
    29384 => 20,
    29385 => 20,
    29386 => 20,
    29387 => 20,
    29388 => 20,
    29389 => 20,
    29390 => 20,
    29391 => 20,
    29392 => 20,
    29393 => 20,
    29394 => 20,
    29395 => 20,
    29396 => 20,
    29397 => 20,
    29398 => 20,
    29399 => 20,
    29400 => 20,
    29401 => 20,
    29402 => 20,
    29403 => 20,
    29404 => 20,
    29405 => 20,
    29406 => 20,
    29407 => 20,
    29408 => 20,
    29409 => 20,
    29410 => 20,
    29411 => 20,
    29412 => 20,
    29413 => 20,
    29414 => 20,
    29415 => 20,
    29416 => 20,
    29417 => 20,
    29418 => 20,
    29419 => 20,
    29420 => 20,
    29421 => 20,
    29422 => 20,
    29423 => 20,
    29424 => 20,
    29425 => 20,
    29426 => 20,
    29427 => 20,
    29428 => 20,
    29429 => 20,
    29430 => 20,
    29431 => 20,
    29432 => 20,
    29433 => 20,
    29434 => 20,
    29435 => 20,
    29436 => 20,
    29437 => 20,
    29438 => 20,
    29439 => 20,
    29440 => 20,
    29441 => 20,
    29442 => 20,
    29443 => 20,
    29444 => 20,
    29445 => 20,
    29446 => 20,
    29447 => 20,
    29448 => 20,
    29449 => 20,
    29450 => 20,
    29451 => 20,
    29452 => 20,
    29453 => 20,
    29454 => 20,
    29455 => 20,
    29456 => 20,
    29457 => 20,
    29458 => 20,
    29459 => 20,
    29460 => 20,
    29461 => 20,
    29462 => 20,
    29463 => 20,
    29464 => 20,
    29465 => 20,
    29466 => 20,
    29467 => 20,
    29468 => 20,
    29469 => 20,
    29470 => 20,
    29471 => 20,
    29472 => 20,
    29473 => 20,
    29474 => 20,
    29475 => 20,
    29476 => 20,
    29477 => 20,
    29478 => 20,
    29479 => 20,
    29480 => 20,
    29481 => 20,
    29482 => 20,
    29483 => 20,
    29484 => 20,
    29485 => 20,
    29486 => 19,
    29487 => 19,
    29488 => 19,
    29489 => 19,
    29490 => 19,
    29491 => 19,
    29492 => 19,
    29493 => 19,
    29494 => 19,
    29495 => 19,
    29496 => 19,
    29497 => 19,
    29498 => 19,
    29499 => 19,
    29500 => 19,
    29501 => 19,
    29502 => 19,
    29503 => 19,
    29504 => 19,
    29505 => 19,
    29506 => 19,
    29507 => 19,
    29508 => 19,
    29509 => 19,
    29510 => 19,
    29511 => 19,
    29512 => 19,
    29513 => 19,
    29514 => 19,
    29515 => 19,
    29516 => 19,
    29517 => 19,
    29518 => 19,
    29519 => 19,
    29520 => 19,
    29521 => 19,
    29522 => 19,
    29523 => 19,
    29524 => 19,
    29525 => 19,
    29526 => 19,
    29527 => 19,
    29528 => 19,
    29529 => 19,
    29530 => 19,
    29531 => 19,
    29532 => 19,
    29533 => 19,
    29534 => 19,
    29535 => 19,
    29536 => 19,
    29537 => 19,
    29538 => 19,
    29539 => 19,
    29540 => 19,
    29541 => 19,
    29542 => 19,
    29543 => 19,
    29544 => 19,
    29545 => 19,
    29546 => 19,
    29547 => 19,
    29548 => 19,
    29549 => 19,
    29550 => 19,
    29551 => 19,
    29552 => 19,
    29553 => 19,
    29554 => 19,
    29555 => 19,
    29556 => 19,
    29557 => 19,
    29558 => 19,
    29559 => 19,
    29560 => 19,
    29561 => 19,
    29562 => 19,
    29563 => 19,
    29564 => 19,
    29565 => 19,
    29566 => 19,
    29567 => 19,
    29568 => 19,
    29569 => 19,
    29570 => 19,
    29571 => 19,
    29572 => 19,
    29573 => 19,
    29574 => 19,
    29575 => 19,
    29576 => 19,
    29577 => 19,
    29578 => 19,
    29579 => 19,
    29580 => 19,
    29581 => 19,
    29582 => 19,
    29583 => 19,
    29584 => 19,
    29585 => 19,
    29586 => 19,
    29587 => 19,
    29588 => 19,
    29589 => 19,
    29590 => 19,
    29591 => 19,
    29592 => 19,
    29593 => 19,
    29594 => 19,
    29595 => 19,
    29596 => 19,
    29597 => 19,
    29598 => 19,
    29599 => 19,
    29600 => 19,
    29601 => 19,
    29602 => 19,
    29603 => 19,
    29604 => 19,
    29605 => 19,
    29606 => 19,
    29607 => 19,
    29608 => 19,
    29609 => 19,
    29610 => 19,
    29611 => 19,
    29612 => 19,
    29613 => 19,
    29614 => 19,
    29615 => 19,
    29616 => 19,
    29617 => 19,
    29618 => 19,
    29619 => 19,
    29620 => 19,
    29621 => 19,
    29622 => 19,
    29623 => 19,
    29624 => 19,
    29625 => 19,
    29626 => 19,
    29627 => 19,
    29628 => 19,
    29629 => 19,
    29630 => 19,
    29631 => 19,
    29632 => 19,
    29633 => 19,
    29634 => 19,
    29635 => 19,
    29636 => 19,
    29637 => 19,
    29638 => 19,
    29639 => 19,
    29640 => 19,
    29641 => 19,
    29642 => 19,
    29643 => 19,
    29644 => 19,
    29645 => 19,
    29646 => 19,
    29647 => 19,
    29648 => 19,
    29649 => 19,
    29650 => 19,
    29651 => 19,
    29652 => 19,
    29653 => 19,
    29654 => 19,
    29655 => 19,
    29656 => 19,
    29657 => 19,
    29658 => 19,
    29659 => 19,
    29660 => 18,
    29661 => 18,
    29662 => 18,
    29663 => 18,
    29664 => 18,
    29665 => 18,
    29666 => 18,
    29667 => 18,
    29668 => 18,
    29669 => 18,
    29670 => 18,
    29671 => 18,
    29672 => 18,
    29673 => 18,
    29674 => 18,
    29675 => 18,
    29676 => 18,
    29677 => 18,
    29678 => 18,
    29679 => 18,
    29680 => 18,
    29681 => 18,
    29682 => 18,
    29683 => 18,
    29684 => 18,
    29685 => 18,
    29686 => 18,
    29687 => 18,
    29688 => 18,
    29689 => 18,
    29690 => 18,
    29691 => 18,
    29692 => 18,
    29693 => 18,
    29694 => 18,
    29695 => 18,
    29696 => 18,
    29697 => 18,
    29698 => 18,
    29699 => 18,
    29700 => 18,
    29701 => 18,
    29702 => 18,
    29703 => 18,
    29704 => 18,
    29705 => 18,
    29706 => 18,
    29707 => 18,
    29708 => 18,
    29709 => 18,
    29710 => 18,
    29711 => 18,
    29712 => 18,
    29713 => 18,
    29714 => 18,
    29715 => 18,
    29716 => 18,
    29717 => 18,
    29718 => 18,
    29719 => 18,
    29720 => 18,
    29721 => 18,
    29722 => 18,
    29723 => 18,
    29724 => 18,
    29725 => 18,
    29726 => 18,
    29727 => 18,
    29728 => 18,
    29729 => 18,
    29730 => 18,
    29731 => 18,
    29732 => 18,
    29733 => 18,
    29734 => 18,
    29735 => 18,
    29736 => 18,
    29737 => 18,
    29738 => 18,
    29739 => 18,
    29740 => 18,
    29741 => 18,
    29742 => 18,
    29743 => 18,
    29744 => 18,
    29745 => 18,
    29746 => 18,
    29747 => 18,
    29748 => 18,
    29749 => 18,
    29750 => 18,
    29751 => 18,
    29752 => 18,
    29753 => 18,
    29754 => 18,
    29755 => 18,
    29756 => 18,
    29757 => 18,
    29758 => 18,
    29759 => 18,
    29760 => 18,
    29761 => 18,
    29762 => 18,
    29763 => 18,
    29764 => 18,
    29765 => 18,
    29766 => 18,
    29767 => 18,
    29768 => 18,
    29769 => 18,
    29770 => 18,
    29771 => 18,
    29772 => 18,
    29773 => 18,
    29774 => 18,
    29775 => 18,
    29776 => 18,
    29777 => 18,
    29778 => 18,
    29779 => 18,
    29780 => 18,
    29781 => 18,
    29782 => 18,
    29783 => 18,
    29784 => 18,
    29785 => 18,
    29786 => 18,
    29787 => 18,
    29788 => 18,
    29789 => 18,
    29790 => 18,
    29791 => 18,
    29792 => 18,
    29793 => 18,
    29794 => 18,
    29795 => 18,
    29796 => 18,
    29797 => 18,
    29798 => 18,
    29799 => 18,
    29800 => 18,
    29801 => 18,
    29802 => 18,
    29803 => 18,
    29804 => 18,
    29805 => 18,
    29806 => 18,
    29807 => 18,
    29808 => 18,
    29809 => 18,
    29810 => 18,
    29811 => 18,
    29812 => 18,
    29813 => 18,
    29814 => 18,
    29815 => 18,
    29816 => 18,
    29817 => 18,
    29818 => 18,
    29819 => 18,
    29820 => 18,
    29821 => 18,
    29822 => 18,
    29823 => 18,
    29824 => 18,
    29825 => 18,
    29826 => 18,
    29827 => 18,
    29828 => 18,
    29829 => 18,
    29830 => 18,
    29831 => 18,
    29832 => 18,
    29833 => 17,
    29834 => 17,
    29835 => 17,
    29836 => 17,
    29837 => 17,
    29838 => 17,
    29839 => 17,
    29840 => 17,
    29841 => 17,
    29842 => 17,
    29843 => 17,
    29844 => 17,
    29845 => 17,
    29846 => 17,
    29847 => 17,
    29848 => 17,
    29849 => 17,
    29850 => 17,
    29851 => 17,
    29852 => 17,
    29853 => 17,
    29854 => 17,
    29855 => 17,
    29856 => 17,
    29857 => 17,
    29858 => 17,
    29859 => 17,
    29860 => 17,
    29861 => 17,
    29862 => 17,
    29863 => 17,
    29864 => 17,
    29865 => 17,
    29866 => 17,
    29867 => 17,
    29868 => 17,
    29869 => 17,
    29870 => 17,
    29871 => 17,
    29872 => 17,
    29873 => 17,
    29874 => 17,
    29875 => 17,
    29876 => 17,
    29877 => 17,
    29878 => 17,
    29879 => 17,
    29880 => 17,
    29881 => 17,
    29882 => 17,
    29883 => 17,
    29884 => 17,
    29885 => 17,
    29886 => 17,
    29887 => 17,
    29888 => 17,
    29889 => 17,
    29890 => 17,
    29891 => 17,
    29892 => 17,
    29893 => 17,
    29894 => 17,
    29895 => 17,
    29896 => 17,
    29897 => 17,
    29898 => 17,
    29899 => 17,
    29900 => 17,
    29901 => 17,
    29902 => 17,
    29903 => 17,
    29904 => 17,
    29905 => 17,
    29906 => 17,
    29907 => 17,
    29908 => 17,
    29909 => 17,
    29910 => 17,
    29911 => 17,
    29912 => 17,
    29913 => 17,
    29914 => 17,
    29915 => 17,
    29916 => 17,
    29917 => 17,
    29918 => 17,
    29919 => 17,
    29920 => 17,
    29921 => 17,
    29922 => 17,
    29923 => 17,
    29924 => 17,
    29925 => 17,
    29926 => 17,
    29927 => 17,
    29928 => 17,
    29929 => 17,
    29930 => 17,
    29931 => 17,
    29932 => 17,
    29933 => 17,
    29934 => 17,
    29935 => 17,
    29936 => 17,
    29937 => 17,
    29938 => 17,
    29939 => 17,
    29940 => 17,
    29941 => 17,
    29942 => 17,
    29943 => 17,
    29944 => 17,
    29945 => 17,
    29946 => 17,
    29947 => 17,
    29948 => 17,
    29949 => 17,
    29950 => 17,
    29951 => 17,
    29952 => 17,
    29953 => 17,
    29954 => 17,
    29955 => 17,
    29956 => 17,
    29957 => 17,
    29958 => 17,
    29959 => 17,
    29960 => 17,
    29961 => 17,
    29962 => 17,
    29963 => 17,
    29964 => 17,
    29965 => 17,
    29966 => 17,
    29967 => 17,
    29968 => 17,
    29969 => 17,
    29970 => 17,
    29971 => 17,
    29972 => 17,
    29973 => 17,
    29974 => 17,
    29975 => 17,
    29976 => 17,
    29977 => 17,
    29978 => 17,
    29979 => 17,
    29980 => 17,
    29981 => 17,
    29982 => 17,
    29983 => 17,
    29984 => 17,
    29985 => 17,
    29986 => 17,
    29987 => 17,
    29988 => 17,
    29989 => 17,
    29990 => 17,
    29991 => 17,
    29992 => 17,
    29993 => 17,
    29994 => 17,
    29995 => 17,
    29996 => 17,
    29997 => 17,
    29998 => 17,
    29999 => 17,
    30000 => 17,
    30001 => 17,
    30002 => 17,
    30003 => 17,
    30004 => 16,
    30005 => 16,
    30006 => 16,
    30007 => 16,
    30008 => 16,
    30009 => 16,
    30010 => 16,
    30011 => 16,
    30012 => 16,
    30013 => 16,
    30014 => 16,
    30015 => 16,
    30016 => 16,
    30017 => 16,
    30018 => 16,
    30019 => 16,
    30020 => 16,
    30021 => 16,
    30022 => 16,
    30023 => 16,
    30024 => 16,
    30025 => 16,
    30026 => 16,
    30027 => 16,
    30028 => 16,
    30029 => 16,
    30030 => 16,
    30031 => 16,
    30032 => 16,
    30033 => 16,
    30034 => 16,
    30035 => 16,
    30036 => 16,
    30037 => 16,
    30038 => 16,
    30039 => 16,
    30040 => 16,
    30041 => 16,
    30042 => 16,
    30043 => 16,
    30044 => 16,
    30045 => 16,
    30046 => 16,
    30047 => 16,
    30048 => 16,
    30049 => 16,
    30050 => 16,
    30051 => 16,
    30052 => 16,
    30053 => 16,
    30054 => 16,
    30055 => 16,
    30056 => 16,
    30057 => 16,
    30058 => 16,
    30059 => 16,
    30060 => 16,
    30061 => 16,
    30062 => 16,
    30063 => 16,
    30064 => 16,
    30065 => 16,
    30066 => 16,
    30067 => 16,
    30068 => 16,
    30069 => 16,
    30070 => 16,
    30071 => 16,
    30072 => 16,
    30073 => 16,
    30074 => 16,
    30075 => 16,
    30076 => 16,
    30077 => 16,
    30078 => 16,
    30079 => 16,
    30080 => 16,
    30081 => 16,
    30082 => 16,
    30083 => 16,
    30084 => 16,
    30085 => 16,
    30086 => 16,
    30087 => 16,
    30088 => 16,
    30089 => 16,
    30090 => 16,
    30091 => 16,
    30092 => 16,
    30093 => 16,
    30094 => 16,
    30095 => 16,
    30096 => 16,
    30097 => 16,
    30098 => 16,
    30099 => 16,
    30100 => 16,
    30101 => 16,
    30102 => 16,
    30103 => 16,
    30104 => 16,
    30105 => 16,
    30106 => 16,
    30107 => 16,
    30108 => 16,
    30109 => 16,
    30110 => 16,
    30111 => 16,
    30112 => 16,
    30113 => 16,
    30114 => 16,
    30115 => 16,
    30116 => 16,
    30117 => 16,
    30118 => 16,
    30119 => 16,
    30120 => 16,
    30121 => 16,
    30122 => 16,
    30123 => 16,
    30124 => 16,
    30125 => 16,
    30126 => 16,
    30127 => 16,
    30128 => 16,
    30129 => 16,
    30130 => 16,
    30131 => 16,
    30132 => 16,
    30133 => 16,
    30134 => 16,
    30135 => 16,
    30136 => 16,
    30137 => 16,
    30138 => 16,
    30139 => 16,
    30140 => 16,
    30141 => 16,
    30142 => 16,
    30143 => 16,
    30144 => 16,
    30145 => 16,
    30146 => 16,
    30147 => 16,
    30148 => 16,
    30149 => 16,
    30150 => 16,
    30151 => 16,
    30152 => 16,
    30153 => 16,
    30154 => 16,
    30155 => 16,
    30156 => 16,
    30157 => 16,
    30158 => 16,
    30159 => 16,
    30160 => 16,
    30161 => 16,
    30162 => 16,
    30163 => 16,
    30164 => 16,
    30165 => 16,
    30166 => 16,
    30167 => 16,
    30168 => 16,
    30169 => 16,
    30170 => 16,
    30171 => 16,
    30172 => 16,
    30173 => 16,
    30174 => 16,
    30175 => 16,
    30176 => 15,
    30177 => 15,
    30178 => 15,
    30179 => 15,
    30180 => 15,
    30181 => 15,
    30182 => 15,
    30183 => 15,
    30184 => 15,
    30185 => 15,
    30186 => 15,
    30187 => 15,
    30188 => 15,
    30189 => 15,
    30190 => 15,
    30191 => 15,
    30192 => 15,
    30193 => 15,
    30194 => 15,
    30195 => 15,
    30196 => 15,
    30197 => 15,
    30198 => 15,
    30199 => 15,
    30200 => 15,
    30201 => 15,
    30202 => 15,
    30203 => 15,
    30204 => 15,
    30205 => 15,
    30206 => 15,
    30207 => 15,
    30208 => 15,
    30209 => 15,
    30210 => 15,
    30211 => 15,
    30212 => 15,
    30213 => 15,
    30214 => 15,
    30215 => 15,
    30216 => 15,
    30217 => 15,
    30218 => 15,
    30219 => 15,
    30220 => 15,
    30221 => 15,
    30222 => 15,
    30223 => 15,
    30224 => 15,
    30225 => 15,
    30226 => 15,
    30227 => 15,
    30228 => 15,
    30229 => 15,
    30230 => 15,
    30231 => 15,
    30232 => 15,
    30233 => 15,
    30234 => 15,
    30235 => 15,
    30236 => 15,
    30237 => 15,
    30238 => 15,
    30239 => 15,
    30240 => 15,
    30241 => 15,
    30242 => 15,
    30243 => 15,
    30244 => 15,
    30245 => 15,
    30246 => 15,
    30247 => 15,
    30248 => 15,
    30249 => 15,
    30250 => 15,
    30251 => 15,
    30252 => 15,
    30253 => 15,
    30254 => 15,
    30255 => 15,
    30256 => 15,
    30257 => 15,
    30258 => 15,
    30259 => 15,
    30260 => 15,
    30261 => 15,
    30262 => 15,
    30263 => 15,
    30264 => 15,
    30265 => 15,
    30266 => 15,
    30267 => 15,
    30268 => 15,
    30269 => 15,
    30270 => 15,
    30271 => 15,
    30272 => 15,
    30273 => 15,
    30274 => 15,
    30275 => 15,
    30276 => 15,
    30277 => 15,
    30278 => 15,
    30279 => 15,
    30280 => 15,
    30281 => 15,
    30282 => 15,
    30283 => 15,
    30284 => 15,
    30285 => 15,
    30286 => 15,
    30287 => 15,
    30288 => 15,
    30289 => 15,
    30290 => 15,
    30291 => 15,
    30292 => 15,
    30293 => 15,
    30294 => 15,
    30295 => 15,
    30296 => 15,
    30297 => 15,
    30298 => 15,
    30299 => 15,
    30300 => 15,
    30301 => 15,
    30302 => 15,
    30303 => 15,
    30304 => 15,
    30305 => 15,
    30306 => 15,
    30307 => 15,
    30308 => 15,
    30309 => 15,
    30310 => 15,
    30311 => 15,
    30312 => 15,
    30313 => 15,
    30314 => 15,
    30315 => 15,
    30316 => 15,
    30317 => 15,
    30318 => 15,
    30319 => 15,
    30320 => 15,
    30321 => 15,
    30322 => 15,
    30323 => 15,
    30324 => 15,
    30325 => 15,
    30326 => 15,
    30327 => 15,
    30328 => 15,
    30329 => 15,
    30330 => 15,
    30331 => 15,
    30332 => 15,
    30333 => 15,
    30334 => 15,
    30335 => 15,
    30336 => 15,
    30337 => 15,
    30338 => 15,
    30339 => 15,
    30340 => 15,
    30341 => 15,
    30342 => 15,
    30343 => 15,
    30344 => 15,
    30345 => 15,
    30346 => 14,
    30347 => 14,
    30348 => 14,
    30349 => 14,
    30350 => 14,
    30351 => 14,
    30352 => 14,
    30353 => 14,
    30354 => 14,
    30355 => 14,
    30356 => 14,
    30357 => 14,
    30358 => 14,
    30359 => 14,
    30360 => 14,
    30361 => 14,
    30362 => 14,
    30363 => 14,
    30364 => 14,
    30365 => 14,
    30366 => 14,
    30367 => 14,
    30368 => 14,
    30369 => 14,
    30370 => 14,
    30371 => 14,
    30372 => 14,
    30373 => 14,
    30374 => 14,
    30375 => 14,
    30376 => 14,
    30377 => 14,
    30378 => 14,
    30379 => 14,
    30380 => 14,
    30381 => 14,
    30382 => 14,
    30383 => 14,
    30384 => 14,
    30385 => 14,
    30386 => 14,
    30387 => 14,
    30388 => 14,
    30389 => 14,
    30390 => 14,
    30391 => 14,
    30392 => 14,
    30393 => 14,
    30394 => 14,
    30395 => 14,
    30396 => 14,
    30397 => 14,
    30398 => 14,
    30399 => 14,
    30400 => 14,
    30401 => 14,
    30402 => 14,
    30403 => 14,
    30404 => 14,
    30405 => 14,
    30406 => 14,
    30407 => 14,
    30408 => 14,
    30409 => 14,
    30410 => 14,
    30411 => 14,
    30412 => 14,
    30413 => 14,
    30414 => 14,
    30415 => 14,
    30416 => 14,
    30417 => 14,
    30418 => 14,
    30419 => 14,
    30420 => 14,
    30421 => 14,
    30422 => 14,
    30423 => 14,
    30424 => 14,
    30425 => 14,
    30426 => 14,
    30427 => 14,
    30428 => 14,
    30429 => 14,
    30430 => 14,
    30431 => 14,
    30432 => 14,
    30433 => 14,
    30434 => 14,
    30435 => 14,
    30436 => 14,
    30437 => 14,
    30438 => 14,
    30439 => 14,
    30440 => 14,
    30441 => 14,
    30442 => 14,
    30443 => 14,
    30444 => 14,
    30445 => 14,
    30446 => 14,
    30447 => 14,
    30448 => 14,
    30449 => 14,
    30450 => 14,
    30451 => 14,
    30452 => 14,
    30453 => 14,
    30454 => 14,
    30455 => 14,
    30456 => 14,
    30457 => 14,
    30458 => 14,
    30459 => 14,
    30460 => 14,
    30461 => 14,
    30462 => 14,
    30463 => 14,
    30464 => 14,
    30465 => 14,
    30466 => 14,
    30467 => 14,
    30468 => 14,
    30469 => 14,
    30470 => 14,
    30471 => 14,
    30472 => 14,
    30473 => 14,
    30474 => 14,
    30475 => 14,
    30476 => 14,
    30477 => 14,
    30478 => 14,
    30479 => 14,
    30480 => 14,
    30481 => 14,
    30482 => 14,
    30483 => 14,
    30484 => 14,
    30485 => 14,
    30486 => 14,
    30487 => 14,
    30488 => 14,
    30489 => 14,
    30490 => 14,
    30491 => 14,
    30492 => 14,
    30493 => 14,
    30494 => 14,
    30495 => 14,
    30496 => 14,
    30497 => 14,
    30498 => 14,
    30499 => 14,
    30500 => 14,
    30501 => 14,
    30502 => 14,
    30503 => 14,
    30504 => 14,
    30505 => 14,
    30506 => 14,
    30507 => 14,
    30508 => 14,
    30509 => 14,
    30510 => 14,
    30511 => 14,
    30512 => 14,
    30513 => 14,
    30514 => 14,
    30515 => 14,
    30516 => 13,
    30517 => 13,
    30518 => 13,
    30519 => 13,
    30520 => 13,
    30521 => 13,
    30522 => 13,
    30523 => 13,
    30524 => 13,
    30525 => 13,
    30526 => 13,
    30527 => 13,
    30528 => 13,
    30529 => 13,
    30530 => 13,
    30531 => 13,
    30532 => 13,
    30533 => 13,
    30534 => 13,
    30535 => 13,
    30536 => 13,
    30537 => 13,
    30538 => 13,
    30539 => 13,
    30540 => 13,
    30541 => 13,
    30542 => 13,
    30543 => 13,
    30544 => 13,
    30545 => 13,
    30546 => 13,
    30547 => 13,
    30548 => 13,
    30549 => 13,
    30550 => 13,
    30551 => 13,
    30552 => 13,
    30553 => 13,
    30554 => 13,
    30555 => 13,
    30556 => 13,
    30557 => 13,
    30558 => 13,
    30559 => 13,
    30560 => 13,
    30561 => 13,
    30562 => 13,
    30563 => 13,
    30564 => 13,
    30565 => 13,
    30566 => 13,
    30567 => 13,
    30568 => 13,
    30569 => 13,
    30570 => 13,
    30571 => 13,
    30572 => 13,
    30573 => 13,
    30574 => 13,
    30575 => 13,
    30576 => 13,
    30577 => 13,
    30578 => 13,
    30579 => 13,
    30580 => 13,
    30581 => 13,
    30582 => 13,
    30583 => 13,
    30584 => 13,
    30585 => 13,
    30586 => 13,
    30587 => 13,
    30588 => 13,
    30589 => 13,
    30590 => 13,
    30591 => 13,
    30592 => 13,
    30593 => 13,
    30594 => 13,
    30595 => 13,
    30596 => 13,
    30597 => 13,
    30598 => 13,
    30599 => 13,
    30600 => 13,
    30601 => 13,
    30602 => 13,
    30603 => 13,
    30604 => 13,
    30605 => 13,
    30606 => 13,
    30607 => 13,
    30608 => 13,
    30609 => 13,
    30610 => 13,
    30611 => 13,
    30612 => 13,
    30613 => 13,
    30614 => 13,
    30615 => 13,
    30616 => 13,
    30617 => 13,
    30618 => 13,
    30619 => 13,
    30620 => 13,
    30621 => 13,
    30622 => 13,
    30623 => 13,
    30624 => 13,
    30625 => 13,
    30626 => 13,
    30627 => 13,
    30628 => 13,
    30629 => 13,
    30630 => 13,
    30631 => 13,
    30632 => 13,
    30633 => 13,
    30634 => 13,
    30635 => 13,
    30636 => 13,
    30637 => 13,
    30638 => 13,
    30639 => 13,
    30640 => 13,
    30641 => 13,
    30642 => 13,
    30643 => 13,
    30644 => 13,
    30645 => 13,
    30646 => 13,
    30647 => 13,
    30648 => 13,
    30649 => 13,
    30650 => 13,
    30651 => 13,
    30652 => 13,
    30653 => 13,
    30654 => 13,
    30655 => 13,
    30656 => 13,
    30657 => 13,
    30658 => 13,
    30659 => 13,
    30660 => 13,
    30661 => 13,
    30662 => 13,
    30663 => 13,
    30664 => 13,
    30665 => 13,
    30666 => 13,
    30667 => 13,
    30668 => 13,
    30669 => 13,
    30670 => 13,
    30671 => 13,
    30672 => 13,
    30673 => 13,
    30674 => 13,
    30675 => 13,
    30676 => 13,
    30677 => 13,
    30678 => 13,
    30679 => 13,
    30680 => 13,
    30681 => 13,
    30682 => 13,
    30683 => 13,
    30684 => 13,
    30685 => 12,
    30686 => 12,
    30687 => 12,
    30688 => 12,
    30689 => 12,
    30690 => 12,
    30691 => 12,
    30692 => 12,
    30693 => 12,
    30694 => 12,
    30695 => 12,
    30696 => 12,
    30697 => 12,
    30698 => 12,
    30699 => 12,
    30700 => 12,
    30701 => 12,
    30702 => 12,
    30703 => 12,
    30704 => 12,
    30705 => 12,
    30706 => 12,
    30707 => 12,
    30708 => 12,
    30709 => 12,
    30710 => 12,
    30711 => 12,
    30712 => 12,
    30713 => 12,
    30714 => 12,
    30715 => 12,
    30716 => 12,
    30717 => 12,
    30718 => 12,
    30719 => 12,
    30720 => 12,
    30721 => 12,
    30722 => 12,
    30723 => 12,
    30724 => 12,
    30725 => 12,
    30726 => 12,
    30727 => 12,
    30728 => 12,
    30729 => 12,
    30730 => 12,
    30731 => 12,
    30732 => 12,
    30733 => 12,
    30734 => 12,
    30735 => 12,
    30736 => 12,
    30737 => 12,
    30738 => 12,
    30739 => 12,
    30740 => 12,
    30741 => 12,
    30742 => 12,
    30743 => 12,
    30744 => 12,
    30745 => 12,
    30746 => 12,
    30747 => 12,
    30748 => 12,
    30749 => 12,
    30750 => 12,
    30751 => 12,
    30752 => 12,
    30753 => 12,
    30754 => 12,
    30755 => 12,
    30756 => 12,
    30757 => 12,
    30758 => 12,
    30759 => 12,
    30760 => 12,
    30761 => 12,
    30762 => 12,
    30763 => 12,
    30764 => 12,
    30765 => 12,
    30766 => 12,
    30767 => 12,
    30768 => 12,
    30769 => 12,
    30770 => 12,
    30771 => 12,
    30772 => 12,
    30773 => 12,
    30774 => 12,
    30775 => 12,
    30776 => 12,
    30777 => 12,
    30778 => 12,
    30779 => 12,
    30780 => 12,
    30781 => 12,
    30782 => 12,
    30783 => 12,
    30784 => 12,
    30785 => 12,
    30786 => 12,
    30787 => 12,
    30788 => 12,
    30789 => 12,
    30790 => 12,
    30791 => 12,
    30792 => 12,
    30793 => 12,
    30794 => 12,
    30795 => 12,
    30796 => 12,
    30797 => 12,
    30798 => 12,
    30799 => 12,
    30800 => 12,
    30801 => 12,
    30802 => 12,
    30803 => 12,
    30804 => 12,
    30805 => 12,
    30806 => 12,
    30807 => 12,
    30808 => 12,
    30809 => 12,
    30810 => 12,
    30811 => 12,
    30812 => 12,
    30813 => 12,
    30814 => 12,
    30815 => 12,
    30816 => 12,
    30817 => 12,
    30818 => 12,
    30819 => 12,
    30820 => 12,
    30821 => 12,
    30822 => 12,
    30823 => 12,
    30824 => 12,
    30825 => 12,
    30826 => 12,
    30827 => 12,
    30828 => 12,
    30829 => 12,
    30830 => 12,
    30831 => 12,
    30832 => 12,
    30833 => 12,
    30834 => 12,
    30835 => 12,
    30836 => 12,
    30837 => 12,
    30838 => 12,
    30839 => 12,
    30840 => 12,
    30841 => 12,
    30842 => 12,
    30843 => 12,
    30844 => 12,
    30845 => 12,
    30846 => 12,
    30847 => 12,
    30848 => 12,
    30849 => 12,
    30850 => 12,
    30851 => 12,
    30852 => 12,
    30853 => 12,
    30854 => 11,
    30855 => 11,
    30856 => 11,
    30857 => 11,
    30858 => 11,
    30859 => 11,
    30860 => 11,
    30861 => 11,
    30862 => 11,
    30863 => 11,
    30864 => 11,
    30865 => 11,
    30866 => 11,
    30867 => 11,
    30868 => 11,
    30869 => 11,
    30870 => 11,
    30871 => 11,
    30872 => 11,
    30873 => 11,
    30874 => 11,
    30875 => 11,
    30876 => 11,
    30877 => 11,
    30878 => 11,
    30879 => 11,
    30880 => 11,
    30881 => 11,
    30882 => 11,
    30883 => 11,
    30884 => 11,
    30885 => 11,
    30886 => 11,
    30887 => 11,
    30888 => 11,
    30889 => 11,
    30890 => 11,
    30891 => 11,
    30892 => 11,
    30893 => 11,
    30894 => 11,
    30895 => 11,
    30896 => 11,
    30897 => 11,
    30898 => 11,
    30899 => 11,
    30900 => 11,
    30901 => 11,
    30902 => 11,
    30903 => 11,
    30904 => 11,
    30905 => 11,
    30906 => 11,
    30907 => 11,
    30908 => 11,
    30909 => 11,
    30910 => 11,
    30911 => 11,
    30912 => 11,
    30913 => 11,
    30914 => 11,
    30915 => 11,
    30916 => 11,
    30917 => 11,
    30918 => 11,
    30919 => 11,
    30920 => 11,
    30921 => 11,
    30922 => 11,
    30923 => 11,
    30924 => 11,
    30925 => 11,
    30926 => 11,
    30927 => 11,
    30928 => 11,
    30929 => 11,
    30930 => 11,
    30931 => 11,
    30932 => 11,
    30933 => 11,
    30934 => 11,
    30935 => 11,
    30936 => 11,
    30937 => 11,
    30938 => 11,
    30939 => 11,
    30940 => 11,
    30941 => 11,
    30942 => 11,
    30943 => 11,
    30944 => 11,
    30945 => 11,
    30946 => 11,
    30947 => 11,
    30948 => 11,
    30949 => 11,
    30950 => 11,
    30951 => 11,
    30952 => 11,
    30953 => 11,
    30954 => 11,
    30955 => 11,
    30956 => 11,
    30957 => 11,
    30958 => 11,
    30959 => 11,
    30960 => 11,
    30961 => 11,
    30962 => 11,
    30963 => 11,
    30964 => 11,
    30965 => 11,
    30966 => 11,
    30967 => 11,
    30968 => 11,
    30969 => 11,
    30970 => 11,
    30971 => 11,
    30972 => 11,
    30973 => 11,
    30974 => 11,
    30975 => 11,
    30976 => 11,
    30977 => 11,
    30978 => 11,
    30979 => 11,
    30980 => 11,
    30981 => 11,
    30982 => 11,
    30983 => 11,
    30984 => 11,
    30985 => 11,
    30986 => 11,
    30987 => 11,
    30988 => 11,
    30989 => 11,
    30990 => 11,
    30991 => 11,
    30992 => 11,
    30993 => 11,
    30994 => 11,
    30995 => 11,
    30996 => 11,
    30997 => 11,
    30998 => 11,
    30999 => 11,
    31000 => 11,
    31001 => 11,
    31002 => 11,
    31003 => 11,
    31004 => 11,
    31005 => 11,
    31006 => 11,
    31007 => 11,
    31008 => 11,
    31009 => 11,
    31010 => 11,
    31011 => 11,
    31012 => 11,
    31013 => 11,
    31014 => 11,
    31015 => 11,
    31016 => 11,
    31017 => 11,
    31018 => 11,
    31019 => 11,
    31020 => 11,
    31021 => 11,
    31022 => 10,
    31023 => 10,
    31024 => 10,
    31025 => 10,
    31026 => 10,
    31027 => 10,
    31028 => 10,
    31029 => 10,
    31030 => 10,
    31031 => 10,
    31032 => 10,
    31033 => 10,
    31034 => 10,
    31035 => 10,
    31036 => 10,
    31037 => 10,
    31038 => 10,
    31039 => 10,
    31040 => 10,
    31041 => 10,
    31042 => 10,
    31043 => 10,
    31044 => 10,
    31045 => 10,
    31046 => 10,
    31047 => 10,
    31048 => 10,
    31049 => 10,
    31050 => 10,
    31051 => 10,
    31052 => 10,
    31053 => 10,
    31054 => 10,
    31055 => 10,
    31056 => 10,
    31057 => 10,
    31058 => 10,
    31059 => 10,
    31060 => 10,
    31061 => 10,
    31062 => 10,
    31063 => 10,
    31064 => 10,
    31065 => 10,
    31066 => 10,
    31067 => 10,
    31068 => 10,
    31069 => 10,
    31070 => 10,
    31071 => 10,
    31072 => 10,
    31073 => 10,
    31074 => 10,
    31075 => 10,
    31076 => 10,
    31077 => 10,
    31078 => 10,
    31079 => 10,
    31080 => 10,
    31081 => 10,
    31082 => 10,
    31083 => 10,
    31084 => 10,
    31085 => 10,
    31086 => 10,
    31087 => 10,
    31088 => 10,
    31089 => 10,
    31090 => 10,
    31091 => 10,
    31092 => 10,
    31093 => 10,
    31094 => 10,
    31095 => 10,
    31096 => 10,
    31097 => 10,
    31098 => 10,
    31099 => 10,
    31100 => 10,
    31101 => 10,
    31102 => 10,
    31103 => 10,
    31104 => 10,
    31105 => 10,
    31106 => 10,
    31107 => 10,
    31108 => 10,
    31109 => 10,
    31110 => 10,
    31111 => 10,
    31112 => 10,
    31113 => 10,
    31114 => 10,
    31115 => 10,
    31116 => 10,
    31117 => 10,
    31118 => 10,
    31119 => 10,
    31120 => 10,
    31121 => 10,
    31122 => 10,
    31123 => 10,
    31124 => 10,
    31125 => 10,
    31126 => 10,
    31127 => 10,
    31128 => 10,
    31129 => 10,
    31130 => 10,
    31131 => 10,
    31132 => 10,
    31133 => 10,
    31134 => 10,
    31135 => 10,
    31136 => 10,
    31137 => 10,
    31138 => 10,
    31139 => 10,
    31140 => 10,
    31141 => 10,
    31142 => 10,
    31143 => 10,
    31144 => 10,
    31145 => 10,
    31146 => 10,
    31147 => 10,
    31148 => 10,
    31149 => 10,
    31150 => 10,
    31151 => 10,
    31152 => 10,
    31153 => 10,
    31154 => 10,
    31155 => 10,
    31156 => 10,
    31157 => 10,
    31158 => 10,
    31159 => 10,
    31160 => 10,
    31161 => 10,
    31162 => 10,
    31163 => 10,
    31164 => 10,
    31165 => 10,
    31166 => 10,
    31167 => 10,
    31168 => 10,
    31169 => 10,
    31170 => 10,
    31171 => 10,
    31172 => 10,
    31173 => 10,
    31174 => 10,
    31175 => 10,
    31176 => 10,
    31177 => 10,
    31178 => 10,
    31179 => 10,
    31180 => 10,
    31181 => 10,
    31182 => 10,
    31183 => 10,
    31184 => 10,
    31185 => 10,
    31186 => 10,
    31187 => 10,
    31188 => 10,
    31189 => 10,
    31190 => 9,
    31191 => 9,
    31192 => 9,
    31193 => 9,
    31194 => 9,
    31195 => 9,
    31196 => 9,
    31197 => 9,
    31198 => 9,
    31199 => 9,
    31200 => 9,
    31201 => 9,
    31202 => 9,
    31203 => 9,
    31204 => 9,
    31205 => 9,
    31206 => 9,
    31207 => 9,
    31208 => 9,
    31209 => 9,
    31210 => 9,
    31211 => 9,
    31212 => 9,
    31213 => 9,
    31214 => 9,
    31215 => 9,
    31216 => 9,
    31217 => 9,
    31218 => 9,
    31219 => 9,
    31220 => 9,
    31221 => 9,
    31222 => 9,
    31223 => 9,
    31224 => 9,
    31225 => 9,
    31226 => 9,
    31227 => 9,
    31228 => 9,
    31229 => 9,
    31230 => 9,
    31231 => 9,
    31232 => 9,
    31233 => 9,
    31234 => 9,
    31235 => 9,
    31236 => 9,
    31237 => 9,
    31238 => 9,
    31239 => 9,
    31240 => 9,
    31241 => 9,
    31242 => 9,
    31243 => 9,
    31244 => 9,
    31245 => 9,
    31246 => 9,
    31247 => 9,
    31248 => 9,
    31249 => 9,
    31250 => 9,
    31251 => 9,
    31252 => 9,
    31253 => 9,
    31254 => 9,
    31255 => 9,
    31256 => 9,
    31257 => 9,
    31258 => 9,
    31259 => 9,
    31260 => 9,
    31261 => 9,
    31262 => 9,
    31263 => 9,
    31264 => 9,
    31265 => 9,
    31266 => 9,
    31267 => 9,
    31268 => 9,
    31269 => 9,
    31270 => 9,
    31271 => 9,
    31272 => 9,
    31273 => 9,
    31274 => 9,
    31275 => 9,
    31276 => 9,
    31277 => 9,
    31278 => 9,
    31279 => 9,
    31280 => 9,
    31281 => 9,
    31282 => 9,
    31283 => 9,
    31284 => 9,
    31285 => 9,
    31286 => 9,
    31287 => 9,
    31288 => 9,
    31289 => 9,
    31290 => 9,
    31291 => 9,
    31292 => 9,
    31293 => 9,
    31294 => 9,
    31295 => 9,
    31296 => 9,
    31297 => 9,
    31298 => 9,
    31299 => 9,
    31300 => 9,
    31301 => 9,
    31302 => 9,
    31303 => 9,
    31304 => 9,
    31305 => 9,
    31306 => 9,
    31307 => 9,
    31308 => 9,
    31309 => 9,
    31310 => 9,
    31311 => 9,
    31312 => 9,
    31313 => 9,
    31314 => 9,
    31315 => 9,
    31316 => 9,
    31317 => 9,
    31318 => 9,
    31319 => 9,
    31320 => 9,
    31321 => 9,
    31322 => 9,
    31323 => 9,
    31324 => 9,
    31325 => 9,
    31326 => 9,
    31327 => 9,
    31328 => 9,
    31329 => 9,
    31330 => 9,
    31331 => 9,
    31332 => 9,
    31333 => 9,
    31334 => 9,
    31335 => 9,
    31336 => 9,
    31337 => 9,
    31338 => 9,
    31339 => 9,
    31340 => 9,
    31341 => 9,
    31342 => 9,
    31343 => 9,
    31344 => 9,
    31345 => 9,
    31346 => 9,
    31347 => 9,
    31348 => 9,
    31349 => 9,
    31350 => 9,
    31351 => 9,
    31352 => 9,
    31353 => 9,
    31354 => 9,
    31355 => 9,
    31356 => 9,
    31357 => 8,
    31358 => 8,
    31359 => 8,
    31360 => 8,
    31361 => 8,
    31362 => 8,
    31363 => 8,
    31364 => 8,
    31365 => 8,
    31366 => 8,
    31367 => 8,
    31368 => 8,
    31369 => 8,
    31370 => 8,
    31371 => 8,
    31372 => 8,
    31373 => 8,
    31374 => 8,
    31375 => 8,
    31376 => 8,
    31377 => 8,
    31378 => 8,
    31379 => 8,
    31380 => 8,
    31381 => 8,
    31382 => 8,
    31383 => 8,
    31384 => 8,
    31385 => 8,
    31386 => 8,
    31387 => 8,
    31388 => 8,
    31389 => 8,
    31390 => 8,
    31391 => 8,
    31392 => 8,
    31393 => 8,
    31394 => 8,
    31395 => 8,
    31396 => 8,
    31397 => 8,
    31398 => 8,
    31399 => 8,
    31400 => 8,
    31401 => 8,
    31402 => 8,
    31403 => 8,
    31404 => 8,
    31405 => 8,
    31406 => 8,
    31407 => 8,
    31408 => 8,
    31409 => 8,
    31410 => 8,
    31411 => 8,
    31412 => 8,
    31413 => 8,
    31414 => 8,
    31415 => 8,
    31416 => 8,
    31417 => 8,
    31418 => 8,
    31419 => 8,
    31420 => 8,
    31421 => 8,
    31422 => 8,
    31423 => 8,
    31424 => 8,
    31425 => 8,
    31426 => 8,
    31427 => 8,
    31428 => 8,
    31429 => 8,
    31430 => 8,
    31431 => 8,
    31432 => 8,
    31433 => 8,
    31434 => 8,
    31435 => 8,
    31436 => 8,
    31437 => 8,
    31438 => 8,
    31439 => 8,
    31440 => 8,
    31441 => 8,
    31442 => 8,
    31443 => 8,
    31444 => 8,
    31445 => 8,
    31446 => 8,
    31447 => 8,
    31448 => 8,
    31449 => 8,
    31450 => 8,
    31451 => 8,
    31452 => 8,
    31453 => 8,
    31454 => 8,
    31455 => 8,
    31456 => 8,
    31457 => 8,
    31458 => 8,
    31459 => 8,
    31460 => 8,
    31461 => 8,
    31462 => 8,
    31463 => 8,
    31464 => 8,
    31465 => 8,
    31466 => 8,
    31467 => 8,
    31468 => 8,
    31469 => 8,
    31470 => 8,
    31471 => 8,
    31472 => 8,
    31473 => 8,
    31474 => 8,
    31475 => 8,
    31476 => 8,
    31477 => 8,
    31478 => 8,
    31479 => 8,
    31480 => 8,
    31481 => 8,
    31482 => 8,
    31483 => 8,
    31484 => 8,
    31485 => 8,
    31486 => 8,
    31487 => 8,
    31488 => 8,
    31489 => 8,
    31490 => 8,
    31491 => 8,
    31492 => 8,
    31493 => 8,
    31494 => 8,
    31495 => 8,
    31496 => 8,
    31497 => 8,
    31498 => 8,
    31499 => 8,
    31500 => 8,
    31501 => 8,
    31502 => 8,
    31503 => 8,
    31504 => 8,
    31505 => 8,
    31506 => 8,
    31507 => 8,
    31508 => 8,
    31509 => 8,
    31510 => 8,
    31511 => 8,
    31512 => 8,
    31513 => 8,
    31514 => 8,
    31515 => 8,
    31516 => 8,
    31517 => 8,
    31518 => 8,
    31519 => 8,
    31520 => 8,
    31521 => 8,
    31522 => 8,
    31523 => 8,
    31524 => 7,
    31525 => 7,
    31526 => 7,
    31527 => 7,
    31528 => 7,
    31529 => 7,
    31530 => 7,
    31531 => 7,
    31532 => 7,
    31533 => 7,
    31534 => 7,
    31535 => 7,
    31536 => 7,
    31537 => 7,
    31538 => 7,
    31539 => 7,
    31540 => 7,
    31541 => 7,
    31542 => 7,
    31543 => 7,
    31544 => 7,
    31545 => 7,
    31546 => 7,
    31547 => 7,
    31548 => 7,
    31549 => 7,
    31550 => 7,
    31551 => 7,
    31552 => 7,
    31553 => 7,
    31554 => 7,
    31555 => 7,
    31556 => 7,
    31557 => 7,
    31558 => 7,
    31559 => 7,
    31560 => 7,
    31561 => 7,
    31562 => 7,
    31563 => 7,
    31564 => 7,
    31565 => 7,
    31566 => 7,
    31567 => 7,
    31568 => 7,
    31569 => 7,
    31570 => 7,
    31571 => 7,
    31572 => 7,
    31573 => 7,
    31574 => 7,
    31575 => 7,
    31576 => 7,
    31577 => 7,
    31578 => 7,
    31579 => 7,
    31580 => 7,
    31581 => 7,
    31582 => 7,
    31583 => 7,
    31584 => 7,
    31585 => 7,
    31586 => 7,
    31587 => 7,
    31588 => 7,
    31589 => 7,
    31590 => 7,
    31591 => 7,
    31592 => 7,
    31593 => 7,
    31594 => 7,
    31595 => 7,
    31596 => 7,
    31597 => 7,
    31598 => 7,
    31599 => 7,
    31600 => 7,
    31601 => 7,
    31602 => 7,
    31603 => 7,
    31604 => 7,
    31605 => 7,
    31606 => 7,
    31607 => 7,
    31608 => 7,
    31609 => 7,
    31610 => 7,
    31611 => 7,
    31612 => 7,
    31613 => 7,
    31614 => 7,
    31615 => 7,
    31616 => 7,
    31617 => 7,
    31618 => 7,
    31619 => 7,
    31620 => 7,
    31621 => 7,
    31622 => 7,
    31623 => 7,
    31624 => 7,
    31625 => 7,
    31626 => 7,
    31627 => 7,
    31628 => 7,
    31629 => 7,
    31630 => 7,
    31631 => 7,
    31632 => 7,
    31633 => 7,
    31634 => 7,
    31635 => 7,
    31636 => 7,
    31637 => 7,
    31638 => 7,
    31639 => 7,
    31640 => 7,
    31641 => 7,
    31642 => 7,
    31643 => 7,
    31644 => 7,
    31645 => 7,
    31646 => 7,
    31647 => 7,
    31648 => 7,
    31649 => 7,
    31650 => 7,
    31651 => 7,
    31652 => 7,
    31653 => 7,
    31654 => 7,
    31655 => 7,
    31656 => 7,
    31657 => 7,
    31658 => 7,
    31659 => 7,
    31660 => 7,
    31661 => 7,
    31662 => 7,
    31663 => 7,
    31664 => 7,
    31665 => 7,
    31666 => 7,
    31667 => 7,
    31668 => 7,
    31669 => 7,
    31670 => 7,
    31671 => 7,
    31672 => 7,
    31673 => 7,
    31674 => 7,
    31675 => 7,
    31676 => 7,
    31677 => 7,
    31678 => 7,
    31679 => 7,
    31680 => 7,
    31681 => 7,
    31682 => 7,
    31683 => 7,
    31684 => 7,
    31685 => 7,
    31686 => 7,
    31687 => 7,
    31688 => 7,
    31689 => 7,
    31690 => 6,
    31691 => 6,
    31692 => 6,
    31693 => 6,
    31694 => 6,
    31695 => 6,
    31696 => 6,
    31697 => 6,
    31698 => 6,
    31699 => 6,
    31700 => 6,
    31701 => 6,
    31702 => 6,
    31703 => 6,
    31704 => 6,
    31705 => 6,
    31706 => 6,
    31707 => 6,
    31708 => 6,
    31709 => 6,
    31710 => 6,
    31711 => 6,
    31712 => 6,
    31713 => 6,
    31714 => 6,
    31715 => 6,
    31716 => 6,
    31717 => 6,
    31718 => 6,
    31719 => 6,
    31720 => 6,
    31721 => 6,
    31722 => 6,
    31723 => 6,
    31724 => 6,
    31725 => 6,
    31726 => 6,
    31727 => 6,
    31728 => 6,
    31729 => 6,
    31730 => 6,
    31731 => 6,
    31732 => 6,
    31733 => 6,
    31734 => 6,
    31735 => 6,
    31736 => 6,
    31737 => 6,
    31738 => 6,
    31739 => 6,
    31740 => 6,
    31741 => 6,
    31742 => 6,
    31743 => 6,
    31744 => 6,
    31745 => 6,
    31746 => 6,
    31747 => 6,
    31748 => 6,
    31749 => 6,
    31750 => 6,
    31751 => 6,
    31752 => 6,
    31753 => 6,
    31754 => 6,
    31755 => 6,
    31756 => 6,
    31757 => 6,
    31758 => 6,
    31759 => 6,
    31760 => 6,
    31761 => 6,
    31762 => 6,
    31763 => 6,
    31764 => 6,
    31765 => 6,
    31766 => 6,
    31767 => 6,
    31768 => 6,
    31769 => 6,
    31770 => 6,
    31771 => 6,
    31772 => 6,
    31773 => 6,
    31774 => 6,
    31775 => 6,
    31776 => 6,
    31777 => 6,
    31778 => 6,
    31779 => 6,
    31780 => 6,
    31781 => 6,
    31782 => 6,
    31783 => 6,
    31784 => 6,
    31785 => 6,
    31786 => 6,
    31787 => 6,
    31788 => 6,
    31789 => 6,
    31790 => 6,
    31791 => 6,
    31792 => 6,
    31793 => 6,
    31794 => 6,
    31795 => 6,
    31796 => 6,
    31797 => 6,
    31798 => 6,
    31799 => 6,
    31800 => 6,
    31801 => 6,
    31802 => 6,
    31803 => 6,
    31804 => 6,
    31805 => 6,
    31806 => 6,
    31807 => 6,
    31808 => 6,
    31809 => 6,
    31810 => 6,
    31811 => 6,
    31812 => 6,
    31813 => 6,
    31814 => 6,
    31815 => 6,
    31816 => 6,
    31817 => 6,
    31818 => 6,
    31819 => 6,
    31820 => 6,
    31821 => 6,
    31822 => 6,
    31823 => 6,
    31824 => 6,
    31825 => 6,
    31826 => 6,
    31827 => 6,
    31828 => 6,
    31829 => 6,
    31830 => 6,
    31831 => 6,
    31832 => 6,
    31833 => 6,
    31834 => 6,
    31835 => 6,
    31836 => 6,
    31837 => 6,
    31838 => 6,
    31839 => 6,
    31840 => 6,
    31841 => 6,
    31842 => 6,
    31843 => 6,
    31844 => 6,
    31845 => 6,
    31846 => 6,
    31847 => 6,
    31848 => 6,
    31849 => 6,
    31850 => 6,
    31851 => 6,
    31852 => 6,
    31853 => 6,
    31854 => 6,
    31855 => 6,
    31856 => 6,
    31857 => 5,
    31858 => 5,
    31859 => 5,
    31860 => 5,
    31861 => 5,
    31862 => 5,
    31863 => 5,
    31864 => 5,
    31865 => 5,
    31866 => 5,
    31867 => 5,
    31868 => 5,
    31869 => 5,
    31870 => 5,
    31871 => 5,
    31872 => 5,
    31873 => 5,
    31874 => 5,
    31875 => 5,
    31876 => 5,
    31877 => 5,
    31878 => 5,
    31879 => 5,
    31880 => 5,
    31881 => 5,
    31882 => 5,
    31883 => 5,
    31884 => 5,
    31885 => 5,
    31886 => 5,
    31887 => 5,
    31888 => 5,
    31889 => 5,
    31890 => 5,
    31891 => 5,
    31892 => 5,
    31893 => 5,
    31894 => 5,
    31895 => 5,
    31896 => 5,
    31897 => 5,
    31898 => 5,
    31899 => 5,
    31900 => 5,
    31901 => 5,
    31902 => 5,
    31903 => 5,
    31904 => 5,
    31905 => 5,
    31906 => 5,
    31907 => 5,
    31908 => 5,
    31909 => 5,
    31910 => 5,
    31911 => 5,
    31912 => 5,
    31913 => 5,
    31914 => 5,
    31915 => 5,
    31916 => 5,
    31917 => 5,
    31918 => 5,
    31919 => 5,
    31920 => 5,
    31921 => 5,
    31922 => 5,
    31923 => 5,
    31924 => 5,
    31925 => 5,
    31926 => 5,
    31927 => 5,
    31928 => 5,
    31929 => 5,
    31930 => 5,
    31931 => 5,
    31932 => 5,
    31933 => 5,
    31934 => 5,
    31935 => 5,
    31936 => 5,
    31937 => 5,
    31938 => 5,
    31939 => 5,
    31940 => 5,
    31941 => 5,
    31942 => 5,
    31943 => 5,
    31944 => 5,
    31945 => 5,
    31946 => 5,
    31947 => 5,
    31948 => 5,
    31949 => 5,
    31950 => 5,
    31951 => 5,
    31952 => 5,
    31953 => 5,
    31954 => 5,
    31955 => 5,
    31956 => 5,
    31957 => 5,
    31958 => 5,
    31959 => 5,
    31960 => 5,
    31961 => 5,
    31962 => 5,
    31963 => 5,
    31964 => 5,
    31965 => 5,
    31966 => 5,
    31967 => 5,
    31968 => 5,
    31969 => 5,
    31970 => 5,
    31971 => 5,
    31972 => 5,
    31973 => 5,
    31974 => 5,
    31975 => 5,
    31976 => 5,
    31977 => 5,
    31978 => 5,
    31979 => 5,
    31980 => 5,
    31981 => 5,
    31982 => 5,
    31983 => 5,
    31984 => 5,
    31985 => 5,
    31986 => 5,
    31987 => 5,
    31988 => 5,
    31989 => 5,
    31990 => 5,
    31991 => 5,
    31992 => 5,
    31993 => 5,
    31994 => 5,
    31995 => 5,
    31996 => 5,
    31997 => 5,
    31998 => 5,
    31999 => 5,
    32000 => 5,
    32001 => 5,
    32002 => 5,
    32003 => 5,
    32004 => 5,
    32005 => 5,
    32006 => 5,
    32007 => 5,
    32008 => 5,
    32009 => 5,
    32010 => 5,
    32011 => 5,
    32012 => 5,
    32013 => 5,
    32014 => 5,
    32015 => 5,
    32016 => 5,
    32017 => 5,
    32018 => 5,
    32019 => 5,
    32020 => 5,
    32021 => 5,
    32022 => 5,
    32023 => 4,
    32024 => 4,
    32025 => 4,
    32026 => 4,
    32027 => 4,
    32028 => 4,
    32029 => 4,
    32030 => 4,
    32031 => 4,
    32032 => 4,
    32033 => 4,
    32034 => 4,
    32035 => 4,
    32036 => 4,
    32037 => 4,
    32038 => 4,
    32039 => 4,
    32040 => 4,
    32041 => 4,
    32042 => 4,
    32043 => 4,
    32044 => 4,
    32045 => 4,
    32046 => 4,
    32047 => 4,
    32048 => 4,
    32049 => 4,
    32050 => 4,
    32051 => 4,
    32052 => 4,
    32053 => 4,
    32054 => 4,
    32055 => 4,
    32056 => 4,
    32057 => 4,
    32058 => 4,
    32059 => 4,
    32060 => 4,
    32061 => 4,
    32062 => 4,
    32063 => 4,
    32064 => 4,
    32065 => 4,
    32066 => 4,
    32067 => 4,
    32068 => 4,
    32069 => 4,
    32070 => 4,
    32071 => 4,
    32072 => 4,
    32073 => 4,
    32074 => 4,
    32075 => 4,
    32076 => 4,
    32077 => 4,
    32078 => 4,
    32079 => 4,
    32080 => 4,
    32081 => 4,
    32082 => 4,
    32083 => 4,
    32084 => 4,
    32085 => 4,
    32086 => 4,
    32087 => 4,
    32088 => 4,
    32089 => 4,
    32090 => 4,
    32091 => 4,
    32092 => 4,
    32093 => 4,
    32094 => 4,
    32095 => 4,
    32096 => 4,
    32097 => 4,
    32098 => 4,
    32099 => 4,
    32100 => 4,
    32101 => 4,
    32102 => 4,
    32103 => 4,
    32104 => 4,
    32105 => 4,
    32106 => 4,
    32107 => 4,
    32108 => 4,
    32109 => 4,
    32110 => 4,
    32111 => 4,
    32112 => 4,
    32113 => 4,
    32114 => 4,
    32115 => 4,
    32116 => 4,
    32117 => 4,
    32118 => 4,
    32119 => 4,
    32120 => 4,
    32121 => 4,
    32122 => 4,
    32123 => 4,
    32124 => 4,
    32125 => 4,
    32126 => 4,
    32127 => 4,
    32128 => 4,
    32129 => 4,
    32130 => 4,
    32131 => 4,
    32132 => 4,
    32133 => 4,
    32134 => 4,
    32135 => 4,
    32136 => 4,
    32137 => 4,
    32138 => 4,
    32139 => 4,
    32140 => 4,
    32141 => 4,
    32142 => 4,
    32143 => 4,
    32144 => 4,
    32145 => 4,
    32146 => 4,
    32147 => 4,
    32148 => 4,
    32149 => 4,
    32150 => 4,
    32151 => 4,
    32152 => 4,
    32153 => 4,
    32154 => 4,
    32155 => 4,
    32156 => 4,
    32157 => 4,
    32158 => 4,
    32159 => 4,
    32160 => 4,
    32161 => 4,
    32162 => 4,
    32163 => 4,
    32164 => 4,
    32165 => 4,
    32166 => 4,
    32167 => 4,
    32168 => 4,
    32169 => 4,
    32170 => 4,
    32171 => 4,
    32172 => 4,
    32173 => 4,
    32174 => 4,
    32175 => 4,
    32176 => 4,
    32177 => 4,
    32178 => 4,
    32179 => 4,
    32180 => 4,
    32181 => 4,
    32182 => 4,
    32183 => 4,
    32184 => 4,
    32185 => 4,
    32186 => 4,
    32187 => 4,
    32188 => 4,
    32189 => 3,
    32190 => 3,
    32191 => 3,
    32192 => 3,
    32193 => 3,
    32194 => 3,
    32195 => 3,
    32196 => 3,
    32197 => 3,
    32198 => 3,
    32199 => 3,
    32200 => 3,
    32201 => 3,
    32202 => 3,
    32203 => 3,
    32204 => 3,
    32205 => 3,
    32206 => 3,
    32207 => 3,
    32208 => 3,
    32209 => 3,
    32210 => 3,
    32211 => 3,
    32212 => 3,
    32213 => 3,
    32214 => 3,
    32215 => 3,
    32216 => 3,
    32217 => 3,
    32218 => 3,
    32219 => 3,
    32220 => 3,
    32221 => 3,
    32222 => 3,
    32223 => 3,
    32224 => 3,
    32225 => 3,
    32226 => 3,
    32227 => 3,
    32228 => 3,
    32229 => 3,
    32230 => 3,
    32231 => 3,
    32232 => 3,
    32233 => 3,
    32234 => 3,
    32235 => 3,
    32236 => 3,
    32237 => 3,
    32238 => 3,
    32239 => 3,
    32240 => 3,
    32241 => 3,
    32242 => 3,
    32243 => 3,
    32244 => 3,
    32245 => 3,
    32246 => 3,
    32247 => 3,
    32248 => 3,
    32249 => 3,
    32250 => 3,
    32251 => 3,
    32252 => 3,
    32253 => 3,
    32254 => 3,
    32255 => 3,
    32256 => 3,
    32257 => 3,
    32258 => 3,
    32259 => 3,
    32260 => 3,
    32261 => 3,
    32262 => 3,
    32263 => 3,
    32264 => 3,
    32265 => 3,
    32266 => 3,
    32267 => 3,
    32268 => 3,
    32269 => 3,
    32270 => 3,
    32271 => 3,
    32272 => 3,
    32273 => 3,
    32274 => 3,
    32275 => 3,
    32276 => 3,
    32277 => 3,
    32278 => 3,
    32279 => 3,
    32280 => 3,
    32281 => 3,
    32282 => 3,
    32283 => 3,
    32284 => 3,
    32285 => 3,
    32286 => 3,
    32287 => 3,
    32288 => 3,
    32289 => 3,
    32290 => 3,
    32291 => 3,
    32292 => 3,
    32293 => 3,
    32294 => 3,
    32295 => 3,
    32296 => 3,
    32297 => 3,
    32298 => 3,
    32299 => 3,
    32300 => 3,
    32301 => 3,
    32302 => 3,
    32303 => 3,
    32304 => 3,
    32305 => 3,
    32306 => 3,
    32307 => 3,
    32308 => 3,
    32309 => 3,
    32310 => 3,
    32311 => 3,
    32312 => 3,
    32313 => 3,
    32314 => 3,
    32315 => 3,
    32316 => 3,
    32317 => 3,
    32318 => 3,
    32319 => 3,
    32320 => 3,
    32321 => 3,
    32322 => 3,
    32323 => 3,
    32324 => 3,
    32325 => 3,
    32326 => 3,
    32327 => 3,
    32328 => 3,
    32329 => 3,
    32330 => 3,
    32331 => 3,
    32332 => 3,
    32333 => 3,
    32334 => 3,
    32335 => 3,
    32336 => 3,
    32337 => 3,
    32338 => 3,
    32339 => 3,
    32340 => 3,
    32341 => 3,
    32342 => 3,
    32343 => 3,
    32344 => 3,
    32345 => 3,
    32346 => 3,
    32347 => 3,
    32348 => 3,
    32349 => 3,
    32350 => 3,
    32351 => 3,
    32352 => 3,
    32353 => 3,
    32354 => 2,
    32355 => 2,
    32356 => 2,
    32357 => 2,
    32358 => 2,
    32359 => 2,
    32360 => 2,
    32361 => 2,
    32362 => 2,
    32363 => 2,
    32364 => 2,
    32365 => 2,
    32366 => 2,
    32367 => 2,
    32368 => 2,
    32369 => 2,
    32370 => 2,
    32371 => 2,
    32372 => 2,
    32373 => 2,
    32374 => 2,
    32375 => 2,
    32376 => 2,
    32377 => 2,
    32378 => 2,
    32379 => 2,
    32380 => 2,
    32381 => 2,
    32382 => 2,
    32383 => 2,
    32384 => 2,
    32385 => 2,
    32386 => 2,
    32387 => 2,
    32388 => 2,
    32389 => 2,
    32390 => 2,
    32391 => 2,
    32392 => 2,
    32393 => 2,
    32394 => 2,
    32395 => 2,
    32396 => 2,
    32397 => 2,
    32398 => 2,
    32399 => 2,
    32400 => 2,
    32401 => 2,
    32402 => 2,
    32403 => 2,
    32404 => 2,
    32405 => 2,
    32406 => 2,
    32407 => 2,
    32408 => 2,
    32409 => 2,
    32410 => 2,
    32411 => 2,
    32412 => 2,
    32413 => 2,
    32414 => 2,
    32415 => 2,
    32416 => 2,
    32417 => 2,
    32418 => 2,
    32419 => 2,
    32420 => 2,
    32421 => 2,
    32422 => 2,
    32423 => 2,
    32424 => 2,
    32425 => 2,
    32426 => 2,
    32427 => 2,
    32428 => 2,
    32429 => 2,
    32430 => 2,
    32431 => 2,
    32432 => 2,
    32433 => 2,
    32434 => 2,
    32435 => 2,
    32436 => 2,
    32437 => 2,
    32438 => 2,
    32439 => 2,
    32440 => 2,
    32441 => 2,
    32442 => 2,
    32443 => 2,
    32444 => 2,
    32445 => 2,
    32446 => 2,
    32447 => 2,
    32448 => 2,
    32449 => 2,
    32450 => 2,
    32451 => 2,
    32452 => 2,
    32453 => 2,
    32454 => 2,
    32455 => 2,
    32456 => 2,
    32457 => 2,
    32458 => 2,
    32459 => 2,
    32460 => 2,
    32461 => 2,
    32462 => 2,
    32463 => 2,
    32464 => 2,
    32465 => 2,
    32466 => 2,
    32467 => 2,
    32468 => 2,
    32469 => 2,
    32470 => 2,
    32471 => 2,
    32472 => 2,
    32473 => 2,
    32474 => 2,
    32475 => 2,
    32476 => 2,
    32477 => 2,
    32478 => 2,
    32479 => 2,
    32480 => 2,
    32481 => 2,
    32482 => 2,
    32483 => 2,
    32484 => 2,
    32485 => 2,
    32486 => 2,
    32487 => 2,
    32488 => 2,
    32489 => 2,
    32490 => 2,
    32491 => 2,
    32492 => 2,
    32493 => 2,
    32494 => 2,
    32495 => 2,
    32496 => 2,
    32497 => 2,
    32498 => 2,
    32499 => 2,
    32500 => 2,
    32501 => 2,
    32502 => 2,
    32503 => 2,
    32504 => 2,
    32505 => 2,
    32506 => 2,
    32507 => 2,
    32508 => 2,
    32509 => 2,
    32510 => 2,
    32511 => 2,
    32512 => 2,
    32513 => 2,
    32514 => 2,
    32515 => 2,
    32516 => 2,
    32517 => 2,
    32518 => 2,
    32519 => 2,
    32520 => 1,
    32521 => 1,
    32522 => 1,
    32523 => 1,
    32524 => 1,
    32525 => 1,
    32526 => 1,
    32527 => 1,
    32528 => 1,
    32529 => 1,
    32530 => 1,
    32531 => 1,
    32532 => 1,
    32533 => 1,
    32534 => 1,
    32535 => 1,
    32536 => 1,
    32537 => 1,
    32538 => 1,
    32539 => 1,
    32540 => 1,
    32541 => 1,
    32542 => 1,
    32543 => 1,
    32544 => 1,
    32545 => 1,
    32546 => 1,
    32547 => 1,
    32548 => 1,
    32549 => 1,
    32550 => 1,
    32551 => 1,
    32552 => 1,
    32553 => 1,
    32554 => 1,
    32555 => 1,
    32556 => 1,
    32557 => 1,
    32558 => 1,
    32559 => 1,
    32560 => 1,
    32561 => 1,
    32562 => 1,
    32563 => 1,
    32564 => 1,
    32565 => 1,
    32566 => 1,
    32567 => 1,
    32568 => 1,
    32569 => 1,
    32570 => 1,
    32571 => 1,
    32572 => 1,
    32573 => 1,
    32574 => 1,
    32575 => 1,
    32576 => 1,
    32577 => 1,
    32578 => 1,
    32579 => 1,
    32580 => 1,
    32581 => 1,
    32582 => 1,
    32583 => 1,
    32584 => 1,
    32585 => 1,
    32586 => 1,
    32587 => 1,
    32588 => 1,
    32589 => 1,
    32590 => 1,
    32591 => 1,
    32592 => 1,
    32593 => 1,
    32594 => 1,
    32595 => 1,
    32596 => 1,
    32597 => 1,
    32598 => 1,
    32599 => 1,
    32600 => 1,
    32601 => 1,
    32602 => 1,
    32603 => 1,
    32604 => 1,
    32605 => 1,
    32606 => 1,
    32607 => 1,
    32608 => 1,
    32609 => 1,
    32610 => 1,
    32611 => 1,
    32612 => 1,
    32613 => 1,
    32614 => 1,
    32615 => 1,
    32616 => 1,
    32617 => 1,
    32618 => 1,
    32619 => 1,
    32620 => 1,
    32621 => 1,
    32622 => 1,
    32623 => 1,
    32624 => 1,
    32625 => 1,
    32626 => 1,
    32627 => 1,
    32628 => 1,
    32629 => 1,
    32630 => 1,
    32631 => 1,
    32632 => 1,
    32633 => 1,
    32634 => 1,
    32635 => 1,
    32636 => 1,
    32637 => 1,
    32638 => 1,
    32639 => 1,
    32640 => 1,
    32641 => 1,
    32642 => 1,
    32643 => 1,
    32644 => 1,
    32645 => 1,
    32646 => 1,
    32647 => 1,
    32648 => 1,
    32649 => 1,
    32650 => 1,
    32651 => 1,
    32652 => 1,
    32653 => 1,
    32654 => 1,
    32655 => 1,
    32656 => 1,
    32657 => 1,
    32658 => 1,
    32659 => 1,
    32660 => 1,
    32661 => 1,
    32662 => 1,
    32663 => 1,
    32664 => 1,
    32665 => 1,
    32666 => 1,
    32667 => 1,
    32668 => 1,
    32669 => 1,
    32670 => 1,
    32671 => 1,
    32672 => 1,
    32673 => 1,
    32674 => 1,
    32675 => 1,
    32676 => 1,
    32677 => 1,
    32678 => 1,
    32679 => 1,
    32680 => 1,
    32681 => 1,
    32682 => 1,
    32683 => 1,
    32684 => 1,
    32685 => 1,
    32686 => 0,
    32687 => 0,
    32688 => 0,
    32689 => 0,
    32690 => 0,
    32691 => 0,
    32692 => 0,
    32693 => 0,
    32694 => 0,
    32695 => 0,
    32696 => 0,
    32697 => 0,
    32698 => 0,
    32699 => 0,
    32700 => 0,
    32701 => 0,
    32702 => 0,
    32703 => 0,
    32704 => 0,
    32705 => 0,
    32706 => 0,
    32707 => 0,
    32708 => 0,
    32709 => 0,
    32710 => 0,
    32711 => 0,
    32712 => 0,
    32713 => 0,
    32714 => 0,
    32715 => 0,
    32716 => 0,
    32717 => 0,
    32718 => 0,
    32719 => 0,
    32720 => 0,
    32721 => 0,
    32722 => 0,
    32723 => 0,
    32724 => 0,
    32725 => 0,
    32726 => 0,
    32727 => 0,
    32728 => 0,
    32729 => 0,
    32730 => 0,
    32731 => 0,
    32732 => 0,
    32733 => 0,
    32734 => 0,
    32735 => 0,
    32736 => 0,
    32737 => 0,
    32738 => 0,
    32739 => 0,
    32740 => 0,
    32741 => 0,
    32742 => 0,
    32743 => 0,
    32744 => 0,
    32745 => 0,
    32746 => 0,
    32747 => 0,
    32748 => 0,
    32749 => 0,
    32750 => 0,
    32751 => 0,
    32752 => 0,
    32753 => 0,
    32754 => 0,
    32755 => 0,
    32756 => 0,
    32757 => 0,
    32758 => 0,
    32759 => 0,
    32760 => 0,
    32761 => 0,
    32762 => 0,
    32763 => 0,
    32764 => 0,
    32765 => 0,
    32766 => 0,
    32767 => 0,
    32768 => 0,
    32769 => 0,
    32770 => 0,
    32771 => 0,
    32772 => 0,
    32773 => 0,
    32774 => 0,
    32775 => 0,
    32776 => 0,
    32777 => 0,
    32778 => 0,
    32779 => 0,
    32780 => 0,
    32781 => 0,
    32782 => 0,
    32783 => 0,
    32784 => 0,
    32785 => 0,
    32786 => 0,
    32787 => 0,
    32788 => 0,
    32789 => 0,
    32790 => 0,
    32791 => 0,
    32792 => 0,
    32793 => 0,
    32794 => 0,
    32795 => 0,
    32796 => 0,
    32797 => 0,
    32798 => 0,
    32799 => 0,
    32800 => 0,
    32801 => 0,
    32802 => 0,
    32803 => 0,
    32804 => 0,
    32805 => 0,
    32806 => 0,
    32807 => 0,
    32808 => 0,
    32809 => 0,
    32810 => 0,
    32811 => 0,
    32812 => 0,
    32813 => 0,
    32814 => 0,
    32815 => 0,
    32816 => 0,
    32817 => 0,
    32818 => 0,
    32819 => 0,
    32820 => 0,
    32821 => 0,
    32822 => 0,
    32823 => 0,
    32824 => 0,
    32825 => 0,
    32826 => 0,
    32827 => 0,
    32828 => 0,
    32829 => 0,
    32830 => 0,
    32831 => 0,
    32832 => 0,
    32833 => 0,
    32834 => 0,
    32835 => 0,
    32836 => 0,
    32837 => 0,
    32838 => 0,
    32839 => 0,
    32840 => 0,
    32841 => 0,
    32842 => 0,
    32843 => 0,
    32844 => 0,
    32845 => 0,
    32846 => 0,
    32847 => 0,
    32848 => 0,
    32849 => 0,
    32850 => 0,
    32851 => -1,
    32852 => -1,
    32853 => -1,
    32854 => -1,
    32855 => -1,
    32856 => -1,
    32857 => -1,
    32858 => -1,
    32859 => -1,
    32860 => -1,
    32861 => -1,
    32862 => -1,
    32863 => -1,
    32864 => -1,
    32865 => -1,
    32866 => -1,
    32867 => -1,
    32868 => -1,
    32869 => -1,
    32870 => -1,
    32871 => -1,
    32872 => -1,
    32873 => -1,
    32874 => -1,
    32875 => -1,
    32876 => -1,
    32877 => -1,
    32878 => -1,
    32879 => -1,
    32880 => -1,
    32881 => -1,
    32882 => -1,
    32883 => -1,
    32884 => -1,
    32885 => -1,
    32886 => -1,
    32887 => -1,
    32888 => -1,
    32889 => -1,
    32890 => -1,
    32891 => -1,
    32892 => -1,
    32893 => -1,
    32894 => -1,
    32895 => -1,
    32896 => -1,
    32897 => -1,
    32898 => -1,
    32899 => -1,
    32900 => -1,
    32901 => -1,
    32902 => -1,
    32903 => -1,
    32904 => -1,
    32905 => -1,
    32906 => -1,
    32907 => -1,
    32908 => -1,
    32909 => -1,
    32910 => -1,
    32911 => -1,
    32912 => -1,
    32913 => -1,
    32914 => -1,
    32915 => -1,
    32916 => -1,
    32917 => -1,
    32918 => -1,
    32919 => -1,
    32920 => -1,
    32921 => -1,
    32922 => -1,
    32923 => -1,
    32924 => -1,
    32925 => -1,
    32926 => -1,
    32927 => -1,
    32928 => -1,
    32929 => -1,
    32930 => -1,
    32931 => -1,
    32932 => -1,
    32933 => -1,
    32934 => -1,
    32935 => -1,
    32936 => -1,
    32937 => -1,
    32938 => -1,
    32939 => -1,
    32940 => -1,
    32941 => -1,
    32942 => -1,
    32943 => -1,
    32944 => -1,
    32945 => -1,
    32946 => -1,
    32947 => -1,
    32948 => -1,
    32949 => -1,
    32950 => -1,
    32951 => -1,
    32952 => -1,
    32953 => -1,
    32954 => -1,
    32955 => -1,
    32956 => -1,
    32957 => -1,
    32958 => -1,
    32959 => -1,
    32960 => -1,
    32961 => -1,
    32962 => -1,
    32963 => -1,
    32964 => -1,
    32965 => -1,
    32966 => -1,
    32967 => -1,
    32968 => -1,
    32969 => -1,
    32970 => -1,
    32971 => -1,
    32972 => -1,
    32973 => -1,
    32974 => -1,
    32975 => -1,
    32976 => -1,
    32977 => -1,
    32978 => -1,
    32979 => -1,
    32980 => -1,
    32981 => -1,
    32982 => -1,
    32983 => -1,
    32984 => -1,
    32985 => -1,
    32986 => -1,
    32987 => -1,
    32988 => -1,
    32989 => -1,
    32990 => -1,
    32991 => -1,
    32992 => -1,
    32993 => -1,
    32994 => -1,
    32995 => -1,
    32996 => -1,
    32997 => -1,
    32998 => -1,
    32999 => -1,
    33000 => -1,
    33001 => -1,
    33002 => -1,
    33003 => -1,
    33004 => -1,
    33005 => -1,
    33006 => -1,
    33007 => -1,
    33008 => -1,
    33009 => -1,
    33010 => -1,
    33011 => -1,
    33012 => -1,
    33013 => -1,
    33014 => -1,
    33015 => -1,
    33016 => -1,
    33017 => -2,
    33018 => -2,
    33019 => -2,
    33020 => -2,
    33021 => -2,
    33022 => -2,
    33023 => -2,
    33024 => -2,
    33025 => -2,
    33026 => -2,
    33027 => -2,
    33028 => -2,
    33029 => -2,
    33030 => -2,
    33031 => -2,
    33032 => -2,
    33033 => -2,
    33034 => -2,
    33035 => -2,
    33036 => -2,
    33037 => -2,
    33038 => -2,
    33039 => -2,
    33040 => -2,
    33041 => -2,
    33042 => -2,
    33043 => -2,
    33044 => -2,
    33045 => -2,
    33046 => -2,
    33047 => -2,
    33048 => -2,
    33049 => -2,
    33050 => -2,
    33051 => -2,
    33052 => -2,
    33053 => -2,
    33054 => -2,
    33055 => -2,
    33056 => -2,
    33057 => -2,
    33058 => -2,
    33059 => -2,
    33060 => -2,
    33061 => -2,
    33062 => -2,
    33063 => -2,
    33064 => -2,
    33065 => -2,
    33066 => -2,
    33067 => -2,
    33068 => -2,
    33069 => -2,
    33070 => -2,
    33071 => -2,
    33072 => -2,
    33073 => -2,
    33074 => -2,
    33075 => -2,
    33076 => -2,
    33077 => -2,
    33078 => -2,
    33079 => -2,
    33080 => -2,
    33081 => -2,
    33082 => -2,
    33083 => -2,
    33084 => -2,
    33085 => -2,
    33086 => -2,
    33087 => -2,
    33088 => -2,
    33089 => -2,
    33090 => -2,
    33091 => -2,
    33092 => -2,
    33093 => -2,
    33094 => -2,
    33095 => -2,
    33096 => -2,
    33097 => -2,
    33098 => -2,
    33099 => -2,
    33100 => -2,
    33101 => -2,
    33102 => -2,
    33103 => -2,
    33104 => -2,
    33105 => -2,
    33106 => -2,
    33107 => -2,
    33108 => -2,
    33109 => -2,
    33110 => -2,
    33111 => -2,
    33112 => -2,
    33113 => -2,
    33114 => -2,
    33115 => -2,
    33116 => -2,
    33117 => -2,
    33118 => -2,
    33119 => -2,
    33120 => -2,
    33121 => -2,
    33122 => -2,
    33123 => -2,
    33124 => -2,
    33125 => -2,
    33126 => -2,
    33127 => -2,
    33128 => -2,
    33129 => -2,
    33130 => -2,
    33131 => -2,
    33132 => -2,
    33133 => -2,
    33134 => -2,
    33135 => -2,
    33136 => -2,
    33137 => -2,
    33138 => -2,
    33139 => -2,
    33140 => -2,
    33141 => -2,
    33142 => -2,
    33143 => -2,
    33144 => -2,
    33145 => -2,
    33146 => -2,
    33147 => -2,
    33148 => -2,
    33149 => -2,
    33150 => -2,
    33151 => -2,
    33152 => -2,
    33153 => -2,
    33154 => -2,
    33155 => -2,
    33156 => -2,
    33157 => -2,
    33158 => -2,
    33159 => -2,
    33160 => -2,
    33161 => -2,
    33162 => -2,
    33163 => -2,
    33164 => -2,
    33165 => -2,
    33166 => -2,
    33167 => -2,
    33168 => -2,
    33169 => -2,
    33170 => -2,
    33171 => -2,
    33172 => -2,
    33173 => -2,
    33174 => -2,
    33175 => -2,
    33176 => -2,
    33177 => -2,
    33178 => -2,
    33179 => -2,
    33180 => -2,
    33181 => -2,
    33182 => -2,
    33183 => -3,
    33184 => -3,
    33185 => -3,
    33186 => -3,
    33187 => -3,
    33188 => -3,
    33189 => -3,
    33190 => -3,
    33191 => -3,
    33192 => -3,
    33193 => -3,
    33194 => -3,
    33195 => -3,
    33196 => -3,
    33197 => -3,
    33198 => -3,
    33199 => -3,
    33200 => -3,
    33201 => -3,
    33202 => -3,
    33203 => -3,
    33204 => -3,
    33205 => -3,
    33206 => -3,
    33207 => -3,
    33208 => -3,
    33209 => -3,
    33210 => -3,
    33211 => -3,
    33212 => -3,
    33213 => -3,
    33214 => -3,
    33215 => -3,
    33216 => -3,
    33217 => -3,
    33218 => -3,
    33219 => -3,
    33220 => -3,
    33221 => -3,
    33222 => -3,
    33223 => -3,
    33224 => -3,
    33225 => -3,
    33226 => -3,
    33227 => -3,
    33228 => -3,
    33229 => -3,
    33230 => -3,
    33231 => -3,
    33232 => -3,
    33233 => -3,
    33234 => -3,
    33235 => -3,
    33236 => -3,
    33237 => -3,
    33238 => -3,
    33239 => -3,
    33240 => -3,
    33241 => -3,
    33242 => -3,
    33243 => -3,
    33244 => -3,
    33245 => -3,
    33246 => -3,
    33247 => -3,
    33248 => -3,
    33249 => -3,
    33250 => -3,
    33251 => -3,
    33252 => -3,
    33253 => -3,
    33254 => -3,
    33255 => -3,
    33256 => -3,
    33257 => -3,
    33258 => -3,
    33259 => -3,
    33260 => -3,
    33261 => -3,
    33262 => -3,
    33263 => -3,
    33264 => -3,
    33265 => -3,
    33266 => -3,
    33267 => -3,
    33268 => -3,
    33269 => -3,
    33270 => -3,
    33271 => -3,
    33272 => -3,
    33273 => -3,
    33274 => -3,
    33275 => -3,
    33276 => -3,
    33277 => -3,
    33278 => -3,
    33279 => -3,
    33280 => -3,
    33281 => -3,
    33282 => -3,
    33283 => -3,
    33284 => -3,
    33285 => -3,
    33286 => -3,
    33287 => -3,
    33288 => -3,
    33289 => -3,
    33290 => -3,
    33291 => -3,
    33292 => -3,
    33293 => -3,
    33294 => -3,
    33295 => -3,
    33296 => -3,
    33297 => -3,
    33298 => -3,
    33299 => -3,
    33300 => -3,
    33301 => -3,
    33302 => -3,
    33303 => -3,
    33304 => -3,
    33305 => -3,
    33306 => -3,
    33307 => -3,
    33308 => -3,
    33309 => -3,
    33310 => -3,
    33311 => -3,
    33312 => -3,
    33313 => -3,
    33314 => -3,
    33315 => -3,
    33316 => -3,
    33317 => -3,
    33318 => -3,
    33319 => -3,
    33320 => -3,
    33321 => -3,
    33322 => -3,
    33323 => -3,
    33324 => -3,
    33325 => -3,
    33326 => -3,
    33327 => -3,
    33328 => -3,
    33329 => -3,
    33330 => -3,
    33331 => -3,
    33332 => -3,
    33333 => -3,
    33334 => -3,
    33335 => -3,
    33336 => -3,
    33337 => -3,
    33338 => -3,
    33339 => -3,
    33340 => -3,
    33341 => -3,
    33342 => -3,
    33343 => -3,
    33344 => -3,
    33345 => -3,
    33346 => -3,
    33347 => -3,
    33348 => -4,
    33349 => -4,
    33350 => -4,
    33351 => -4,
    33352 => -4,
    33353 => -4,
    33354 => -4,
    33355 => -4,
    33356 => -4,
    33357 => -4,
    33358 => -4,
    33359 => -4,
    33360 => -4,
    33361 => -4,
    33362 => -4,
    33363 => -4,
    33364 => -4,
    33365 => -4,
    33366 => -4,
    33367 => -4,
    33368 => -4,
    33369 => -4,
    33370 => -4,
    33371 => -4,
    33372 => -4,
    33373 => -4,
    33374 => -4,
    33375 => -4,
    33376 => -4,
    33377 => -4,
    33378 => -4,
    33379 => -4,
    33380 => -4,
    33381 => -4,
    33382 => -4,
    33383 => -4,
    33384 => -4,
    33385 => -4,
    33386 => -4,
    33387 => -4,
    33388 => -4,
    33389 => -4,
    33390 => -4,
    33391 => -4,
    33392 => -4,
    33393 => -4,
    33394 => -4,
    33395 => -4,
    33396 => -4,
    33397 => -4,
    33398 => -4,
    33399 => -4,
    33400 => -4,
    33401 => -4,
    33402 => -4,
    33403 => -4,
    33404 => -4,
    33405 => -4,
    33406 => -4,
    33407 => -4,
    33408 => -4,
    33409 => -4,
    33410 => -4,
    33411 => -4,
    33412 => -4,
    33413 => -4,
    33414 => -4,
    33415 => -4,
    33416 => -4,
    33417 => -4,
    33418 => -4,
    33419 => -4,
    33420 => -4,
    33421 => -4,
    33422 => -4,
    33423 => -4,
    33424 => -4,
    33425 => -4,
    33426 => -4,
    33427 => -4,
    33428 => -4,
    33429 => -4,
    33430 => -4,
    33431 => -4,
    33432 => -4,
    33433 => -4,
    33434 => -4,
    33435 => -4,
    33436 => -4,
    33437 => -4,
    33438 => -4,
    33439 => -4,
    33440 => -4,
    33441 => -4,
    33442 => -4,
    33443 => -4,
    33444 => -4,
    33445 => -4,
    33446 => -4,
    33447 => -4,
    33448 => -4,
    33449 => -4,
    33450 => -4,
    33451 => -4,
    33452 => -4,
    33453 => -4,
    33454 => -4,
    33455 => -4,
    33456 => -4,
    33457 => -4,
    33458 => -4,
    33459 => -4,
    33460 => -4,
    33461 => -4,
    33462 => -4,
    33463 => -4,
    33464 => -4,
    33465 => -4,
    33466 => -4,
    33467 => -4,
    33468 => -4,
    33469 => -4,
    33470 => -4,
    33471 => -4,
    33472 => -4,
    33473 => -4,
    33474 => -4,
    33475 => -4,
    33476 => -4,
    33477 => -4,
    33478 => -4,
    33479 => -4,
    33480 => -4,
    33481 => -4,
    33482 => -4,
    33483 => -4,
    33484 => -4,
    33485 => -4,
    33486 => -4,
    33487 => -4,
    33488 => -4,
    33489 => -4,
    33490 => -4,
    33491 => -4,
    33492 => -4,
    33493 => -4,
    33494 => -4,
    33495 => -4,
    33496 => -4,
    33497 => -4,
    33498 => -4,
    33499 => -4,
    33500 => -4,
    33501 => -4,
    33502 => -4,
    33503 => -4,
    33504 => -4,
    33505 => -4,
    33506 => -4,
    33507 => -4,
    33508 => -4,
    33509 => -4,
    33510 => -4,
    33511 => -4,
    33512 => -4,
    33513 => -4,
    33514 => -5,
    33515 => -5,
    33516 => -5,
    33517 => -5,
    33518 => -5,
    33519 => -5,
    33520 => -5,
    33521 => -5,
    33522 => -5,
    33523 => -5,
    33524 => -5,
    33525 => -5,
    33526 => -5,
    33527 => -5,
    33528 => -5,
    33529 => -5,
    33530 => -5,
    33531 => -5,
    33532 => -5,
    33533 => -5,
    33534 => -5,
    33535 => -5,
    33536 => -5,
    33537 => -5,
    33538 => -5,
    33539 => -5,
    33540 => -5,
    33541 => -5,
    33542 => -5,
    33543 => -5,
    33544 => -5,
    33545 => -5,
    33546 => -5,
    33547 => -5,
    33548 => -5,
    33549 => -5,
    33550 => -5,
    33551 => -5,
    33552 => -5,
    33553 => -5,
    33554 => -5,
    33555 => -5,
    33556 => -5,
    33557 => -5,
    33558 => -5,
    33559 => -5,
    33560 => -5,
    33561 => -5,
    33562 => -5,
    33563 => -5,
    33564 => -5,
    33565 => -5,
    33566 => -5,
    33567 => -5,
    33568 => -5,
    33569 => -5,
    33570 => -5,
    33571 => -5,
    33572 => -5,
    33573 => -5,
    33574 => -5,
    33575 => -5,
    33576 => -5,
    33577 => -5,
    33578 => -5,
    33579 => -5,
    33580 => -5,
    33581 => -5,
    33582 => -5,
    33583 => -5,
    33584 => -5,
    33585 => -5,
    33586 => -5,
    33587 => -5,
    33588 => -5,
    33589 => -5,
    33590 => -5,
    33591 => -5,
    33592 => -5,
    33593 => -5,
    33594 => -5,
    33595 => -5,
    33596 => -5,
    33597 => -5,
    33598 => -5,
    33599 => -5,
    33600 => -5,
    33601 => -5,
    33602 => -5,
    33603 => -5,
    33604 => -5,
    33605 => -5,
    33606 => -5,
    33607 => -5,
    33608 => -5,
    33609 => -5,
    33610 => -5,
    33611 => -5,
    33612 => -5,
    33613 => -5,
    33614 => -5,
    33615 => -5,
    33616 => -5,
    33617 => -5,
    33618 => -5,
    33619 => -5,
    33620 => -5,
    33621 => -5,
    33622 => -5,
    33623 => -5,
    33624 => -5,
    33625 => -5,
    33626 => -5,
    33627 => -5,
    33628 => -5,
    33629 => -5,
    33630 => -5,
    33631 => -5,
    33632 => -5,
    33633 => -5,
    33634 => -5,
    33635 => -5,
    33636 => -5,
    33637 => -5,
    33638 => -5,
    33639 => -5,
    33640 => -5,
    33641 => -5,
    33642 => -5,
    33643 => -5,
    33644 => -5,
    33645 => -5,
    33646 => -5,
    33647 => -5,
    33648 => -5,
    33649 => -5,
    33650 => -5,
    33651 => -5,
    33652 => -5,
    33653 => -5,
    33654 => -5,
    33655 => -5,
    33656 => -5,
    33657 => -5,
    33658 => -5,
    33659 => -5,
    33660 => -5,
    33661 => -5,
    33662 => -5,
    33663 => -5,
    33664 => -5,
    33665 => -5,
    33666 => -5,
    33667 => -5,
    33668 => -5,
    33669 => -5,
    33670 => -5,
    33671 => -5,
    33672 => -5,
    33673 => -5,
    33674 => -5,
    33675 => -5,
    33676 => -5,
    33677 => -5,
    33678 => -5,
    33679 => -5,
    33680 => -6,
    33681 => -6,
    33682 => -6,
    33683 => -6,
    33684 => -6,
    33685 => -6,
    33686 => -6,
    33687 => -6,
    33688 => -6,
    33689 => -6,
    33690 => -6,
    33691 => -6,
    33692 => -6,
    33693 => -6,
    33694 => -6,
    33695 => -6,
    33696 => -6,
    33697 => -6,
    33698 => -6,
    33699 => -6,
    33700 => -6,
    33701 => -6,
    33702 => -6,
    33703 => -6,
    33704 => -6,
    33705 => -6,
    33706 => -6,
    33707 => -6,
    33708 => -6,
    33709 => -6,
    33710 => -6,
    33711 => -6,
    33712 => -6,
    33713 => -6,
    33714 => -6,
    33715 => -6,
    33716 => -6,
    33717 => -6,
    33718 => -6,
    33719 => -6,
    33720 => -6,
    33721 => -6,
    33722 => -6,
    33723 => -6,
    33724 => -6,
    33725 => -6,
    33726 => -6,
    33727 => -6,
    33728 => -6,
    33729 => -6,
    33730 => -6,
    33731 => -6,
    33732 => -6,
    33733 => -6,
    33734 => -6,
    33735 => -6,
    33736 => -6,
    33737 => -6,
    33738 => -6,
    33739 => -6,
    33740 => -6,
    33741 => -6,
    33742 => -6,
    33743 => -6,
    33744 => -6,
    33745 => -6,
    33746 => -6,
    33747 => -6,
    33748 => -6,
    33749 => -6,
    33750 => -6,
    33751 => -6,
    33752 => -6,
    33753 => -6,
    33754 => -6,
    33755 => -6,
    33756 => -6,
    33757 => -6,
    33758 => -6,
    33759 => -6,
    33760 => -6,
    33761 => -6,
    33762 => -6,
    33763 => -6,
    33764 => -6,
    33765 => -6,
    33766 => -6,
    33767 => -6,
    33768 => -6,
    33769 => -6,
    33770 => -6,
    33771 => -6,
    33772 => -6,
    33773 => -6,
    33774 => -6,
    33775 => -6,
    33776 => -6,
    33777 => -6,
    33778 => -6,
    33779 => -6,
    33780 => -6,
    33781 => -6,
    33782 => -6,
    33783 => -6,
    33784 => -6,
    33785 => -6,
    33786 => -6,
    33787 => -6,
    33788 => -6,
    33789 => -6,
    33790 => -6,
    33791 => -6,
    33792 => -6,
    33793 => -6,
    33794 => -6,
    33795 => -6,
    33796 => -6,
    33797 => -6,
    33798 => -6,
    33799 => -6,
    33800 => -6,
    33801 => -6,
    33802 => -6,
    33803 => -6,
    33804 => -6,
    33805 => -6,
    33806 => -6,
    33807 => -6,
    33808 => -6,
    33809 => -6,
    33810 => -6,
    33811 => -6,
    33812 => -6,
    33813 => -6,
    33814 => -6,
    33815 => -6,
    33816 => -6,
    33817 => -6,
    33818 => -6,
    33819 => -6,
    33820 => -6,
    33821 => -6,
    33822 => -6,
    33823 => -6,
    33824 => -6,
    33825 => -6,
    33826 => -6,
    33827 => -6,
    33828 => -6,
    33829 => -6,
    33830 => -6,
    33831 => -6,
    33832 => -6,
    33833 => -6,
    33834 => -6,
    33835 => -6,
    33836 => -6,
    33837 => -6,
    33838 => -6,
    33839 => -6,
    33840 => -6,
    33841 => -6,
    33842 => -6,
    33843 => -6,
    33844 => -6,
    33845 => -6,
    33846 => -6,
    33847 => -7,
    33848 => -7,
    33849 => -7,
    33850 => -7,
    33851 => -7,
    33852 => -7,
    33853 => -7,
    33854 => -7,
    33855 => -7,
    33856 => -7,
    33857 => -7,
    33858 => -7,
    33859 => -7,
    33860 => -7,
    33861 => -7,
    33862 => -7,
    33863 => -7,
    33864 => -7,
    33865 => -7,
    33866 => -7,
    33867 => -7,
    33868 => -7,
    33869 => -7,
    33870 => -7,
    33871 => -7,
    33872 => -7,
    33873 => -7,
    33874 => -7,
    33875 => -7,
    33876 => -7,
    33877 => -7,
    33878 => -7,
    33879 => -7,
    33880 => -7,
    33881 => -7,
    33882 => -7,
    33883 => -7,
    33884 => -7,
    33885 => -7,
    33886 => -7,
    33887 => -7,
    33888 => -7,
    33889 => -7,
    33890 => -7,
    33891 => -7,
    33892 => -7,
    33893 => -7,
    33894 => -7,
    33895 => -7,
    33896 => -7,
    33897 => -7,
    33898 => -7,
    33899 => -7,
    33900 => -7,
    33901 => -7,
    33902 => -7,
    33903 => -7,
    33904 => -7,
    33905 => -7,
    33906 => -7,
    33907 => -7,
    33908 => -7,
    33909 => -7,
    33910 => -7,
    33911 => -7,
    33912 => -7,
    33913 => -7,
    33914 => -7,
    33915 => -7,
    33916 => -7,
    33917 => -7,
    33918 => -7,
    33919 => -7,
    33920 => -7,
    33921 => -7,
    33922 => -7,
    33923 => -7,
    33924 => -7,
    33925 => -7,
    33926 => -7,
    33927 => -7,
    33928 => -7,
    33929 => -7,
    33930 => -7,
    33931 => -7,
    33932 => -7,
    33933 => -7,
    33934 => -7,
    33935 => -7,
    33936 => -7,
    33937 => -7,
    33938 => -7,
    33939 => -7,
    33940 => -7,
    33941 => -7,
    33942 => -7,
    33943 => -7,
    33944 => -7,
    33945 => -7,
    33946 => -7,
    33947 => -7,
    33948 => -7,
    33949 => -7,
    33950 => -7,
    33951 => -7,
    33952 => -7,
    33953 => -7,
    33954 => -7,
    33955 => -7,
    33956 => -7,
    33957 => -7,
    33958 => -7,
    33959 => -7,
    33960 => -7,
    33961 => -7,
    33962 => -7,
    33963 => -7,
    33964 => -7,
    33965 => -7,
    33966 => -7,
    33967 => -7,
    33968 => -7,
    33969 => -7,
    33970 => -7,
    33971 => -7,
    33972 => -7,
    33973 => -7,
    33974 => -7,
    33975 => -7,
    33976 => -7,
    33977 => -7,
    33978 => -7,
    33979 => -7,
    33980 => -7,
    33981 => -7,
    33982 => -7,
    33983 => -7,
    33984 => -7,
    33985 => -7,
    33986 => -7,
    33987 => -7,
    33988 => -7,
    33989 => -7,
    33990 => -7,
    33991 => -7,
    33992 => -7,
    33993 => -7,
    33994 => -7,
    33995 => -7,
    33996 => -7,
    33997 => -7,
    33998 => -7,
    33999 => -7,
    34000 => -7,
    34001 => -7,
    34002 => -7,
    34003 => -7,
    34004 => -7,
    34005 => -7,
    34006 => -7,
    34007 => -7,
    34008 => -7,
    34009 => -7,
    34010 => -7,
    34011 => -7,
    34012 => -7,
    34013 => -8,
    34014 => -8,
    34015 => -8,
    34016 => -8,
    34017 => -8,
    34018 => -8,
    34019 => -8,
    34020 => -8,
    34021 => -8,
    34022 => -8,
    34023 => -8,
    34024 => -8,
    34025 => -8,
    34026 => -8,
    34027 => -8,
    34028 => -8,
    34029 => -8,
    34030 => -8,
    34031 => -8,
    34032 => -8,
    34033 => -8,
    34034 => -8,
    34035 => -8,
    34036 => -8,
    34037 => -8,
    34038 => -8,
    34039 => -8,
    34040 => -8,
    34041 => -8,
    34042 => -8,
    34043 => -8,
    34044 => -8,
    34045 => -8,
    34046 => -8,
    34047 => -8,
    34048 => -8,
    34049 => -8,
    34050 => -8,
    34051 => -8,
    34052 => -8,
    34053 => -8,
    34054 => -8,
    34055 => -8,
    34056 => -8,
    34057 => -8,
    34058 => -8,
    34059 => -8,
    34060 => -8,
    34061 => -8,
    34062 => -8,
    34063 => -8,
    34064 => -8,
    34065 => -8,
    34066 => -8,
    34067 => -8,
    34068 => -8,
    34069 => -8,
    34070 => -8,
    34071 => -8,
    34072 => -8,
    34073 => -8,
    34074 => -8,
    34075 => -8,
    34076 => -8,
    34077 => -8,
    34078 => -8,
    34079 => -8,
    34080 => -8,
    34081 => -8,
    34082 => -8,
    34083 => -8,
    34084 => -8,
    34085 => -8,
    34086 => -8,
    34087 => -8,
    34088 => -8,
    34089 => -8,
    34090 => -8,
    34091 => -8,
    34092 => -8,
    34093 => -8,
    34094 => -8,
    34095 => -8,
    34096 => -8,
    34097 => -8,
    34098 => -8,
    34099 => -8,
    34100 => -8,
    34101 => -8,
    34102 => -8,
    34103 => -8,
    34104 => -8,
    34105 => -8,
    34106 => -8,
    34107 => -8,
    34108 => -8,
    34109 => -8,
    34110 => -8,
    34111 => -8,
    34112 => -8,
    34113 => -8,
    34114 => -8,
    34115 => -8,
    34116 => -8,
    34117 => -8,
    34118 => -8,
    34119 => -8,
    34120 => -8,
    34121 => -8,
    34122 => -8,
    34123 => -8,
    34124 => -8,
    34125 => -8,
    34126 => -8,
    34127 => -8,
    34128 => -8,
    34129 => -8,
    34130 => -8,
    34131 => -8,
    34132 => -8,
    34133 => -8,
    34134 => -8,
    34135 => -8,
    34136 => -8,
    34137 => -8,
    34138 => -8,
    34139 => -8,
    34140 => -8,
    34141 => -8,
    34142 => -8,
    34143 => -8,
    34144 => -8,
    34145 => -8,
    34146 => -8,
    34147 => -8,
    34148 => -8,
    34149 => -8,
    34150 => -8,
    34151 => -8,
    34152 => -8,
    34153 => -8,
    34154 => -8,
    34155 => -8,
    34156 => -8,
    34157 => -8,
    34158 => -8,
    34159 => -8,
    34160 => -8,
    34161 => -8,
    34162 => -8,
    34163 => -8,
    34164 => -8,
    34165 => -8,
    34166 => -8,
    34167 => -8,
    34168 => -8,
    34169 => -8,
    34170 => -8,
    34171 => -8,
    34172 => -8,
    34173 => -8,
    34174 => -8,
    34175 => -8,
    34176 => -8,
    34177 => -8,
    34178 => -8,
    34179 => -8,
    34180 => -9,
    34181 => -9,
    34182 => -9,
    34183 => -9,
    34184 => -9,
    34185 => -9,
    34186 => -9,
    34187 => -9,
    34188 => -9,
    34189 => -9,
    34190 => -9,
    34191 => -9,
    34192 => -9,
    34193 => -9,
    34194 => -9,
    34195 => -9,
    34196 => -9,
    34197 => -9,
    34198 => -9,
    34199 => -9,
    34200 => -9,
    34201 => -9,
    34202 => -9,
    34203 => -9,
    34204 => -9,
    34205 => -9,
    34206 => -9,
    34207 => -9,
    34208 => -9,
    34209 => -9,
    34210 => -9,
    34211 => -9,
    34212 => -9,
    34213 => -9,
    34214 => -9,
    34215 => -9,
    34216 => -9,
    34217 => -9,
    34218 => -9,
    34219 => -9,
    34220 => -9,
    34221 => -9,
    34222 => -9,
    34223 => -9,
    34224 => -9,
    34225 => -9,
    34226 => -9,
    34227 => -9,
    34228 => -9,
    34229 => -9,
    34230 => -9,
    34231 => -9,
    34232 => -9,
    34233 => -9,
    34234 => -9,
    34235 => -9,
    34236 => -9,
    34237 => -9,
    34238 => -9,
    34239 => -9,
    34240 => -9,
    34241 => -9,
    34242 => -9,
    34243 => -9,
    34244 => -9,
    34245 => -9,
    34246 => -9,
    34247 => -9,
    34248 => -9,
    34249 => -9,
    34250 => -9,
    34251 => -9,
    34252 => -9,
    34253 => -9,
    34254 => -9,
    34255 => -9,
    34256 => -9,
    34257 => -9,
    34258 => -9,
    34259 => -9,
    34260 => -9,
    34261 => -9,
    34262 => -9,
    34263 => -9,
    34264 => -9,
    34265 => -9,
    34266 => -9,
    34267 => -9,
    34268 => -9,
    34269 => -9,
    34270 => -9,
    34271 => -9,
    34272 => -9,
    34273 => -9,
    34274 => -9,
    34275 => -9,
    34276 => -9,
    34277 => -9,
    34278 => -9,
    34279 => -9,
    34280 => -9,
    34281 => -9,
    34282 => -9,
    34283 => -9,
    34284 => -9,
    34285 => -9,
    34286 => -9,
    34287 => -9,
    34288 => -9,
    34289 => -9,
    34290 => -9,
    34291 => -9,
    34292 => -9,
    34293 => -9,
    34294 => -9,
    34295 => -9,
    34296 => -9,
    34297 => -9,
    34298 => -9,
    34299 => -9,
    34300 => -9,
    34301 => -9,
    34302 => -9,
    34303 => -9,
    34304 => -9,
    34305 => -9,
    34306 => -9,
    34307 => -9,
    34308 => -9,
    34309 => -9,
    34310 => -9,
    34311 => -9,
    34312 => -9,
    34313 => -9,
    34314 => -9,
    34315 => -9,
    34316 => -9,
    34317 => -9,
    34318 => -9,
    34319 => -9,
    34320 => -9,
    34321 => -9,
    34322 => -9,
    34323 => -9,
    34324 => -9,
    34325 => -9,
    34326 => -9,
    34327 => -9,
    34328 => -9,
    34329 => -9,
    34330 => -9,
    34331 => -9,
    34332 => -9,
    34333 => -9,
    34334 => -9,
    34335 => -9,
    34336 => -9,
    34337 => -9,
    34338 => -9,
    34339 => -9,
    34340 => -9,
    34341 => -9,
    34342 => -9,
    34343 => -9,
    34344 => -9,
    34345 => -9,
    34346 => -9,
    34347 => -10,
    34348 => -10,
    34349 => -10,
    34350 => -10,
    34351 => -10,
    34352 => -10,
    34353 => -10,
    34354 => -10,
    34355 => -10,
    34356 => -10,
    34357 => -10,
    34358 => -10,
    34359 => -10,
    34360 => -10,
    34361 => -10,
    34362 => -10,
    34363 => -10,
    34364 => -10,
    34365 => -10,
    34366 => -10,
    34367 => -10,
    34368 => -10,
    34369 => -10,
    34370 => -10,
    34371 => -10,
    34372 => -10,
    34373 => -10,
    34374 => -10,
    34375 => -10,
    34376 => -10,
    34377 => -10,
    34378 => -10,
    34379 => -10,
    34380 => -10,
    34381 => -10,
    34382 => -10,
    34383 => -10,
    34384 => -10,
    34385 => -10,
    34386 => -10,
    34387 => -10,
    34388 => -10,
    34389 => -10,
    34390 => -10,
    34391 => -10,
    34392 => -10,
    34393 => -10,
    34394 => -10,
    34395 => -10,
    34396 => -10,
    34397 => -10,
    34398 => -10,
    34399 => -10,
    34400 => -10,
    34401 => -10,
    34402 => -10,
    34403 => -10,
    34404 => -10,
    34405 => -10,
    34406 => -10,
    34407 => -10,
    34408 => -10,
    34409 => -10,
    34410 => -10,
    34411 => -10,
    34412 => -10,
    34413 => -10,
    34414 => -10,
    34415 => -10,
    34416 => -10,
    34417 => -10,
    34418 => -10,
    34419 => -10,
    34420 => -10,
    34421 => -10,
    34422 => -10,
    34423 => -10,
    34424 => -10,
    34425 => -10,
    34426 => -10,
    34427 => -10,
    34428 => -10,
    34429 => -10,
    34430 => -10,
    34431 => -10,
    34432 => -10,
    34433 => -10,
    34434 => -10,
    34435 => -10,
    34436 => -10,
    34437 => -10,
    34438 => -10,
    34439 => -10,
    34440 => -10,
    34441 => -10,
    34442 => -10,
    34443 => -10,
    34444 => -10,
    34445 => -10,
    34446 => -10,
    34447 => -10,
    34448 => -10,
    34449 => -10,
    34450 => -10,
    34451 => -10,
    34452 => -10,
    34453 => -10,
    34454 => -10,
    34455 => -10,
    34456 => -10,
    34457 => -10,
    34458 => -10,
    34459 => -10,
    34460 => -10,
    34461 => -10,
    34462 => -10,
    34463 => -10,
    34464 => -10,
    34465 => -10,
    34466 => -10,
    34467 => -10,
    34468 => -10,
    34469 => -10,
    34470 => -10,
    34471 => -10,
    34472 => -10,
    34473 => -10,
    34474 => -10,
    34475 => -10,
    34476 => -10,
    34477 => -10,
    34478 => -10,
    34479 => -10,
    34480 => -10,
    34481 => -10,
    34482 => -10,
    34483 => -10,
    34484 => -10,
    34485 => -10,
    34486 => -10,
    34487 => -10,
    34488 => -10,
    34489 => -10,
    34490 => -10,
    34491 => -10,
    34492 => -10,
    34493 => -10,
    34494 => -10,
    34495 => -10,
    34496 => -10,
    34497 => -10,
    34498 => -10,
    34499 => -10,
    34500 => -10,
    34501 => -10,
    34502 => -10,
    34503 => -10,
    34504 => -10,
    34505 => -10,
    34506 => -10,
    34507 => -10,
    34508 => -10,
    34509 => -10,
    34510 => -10,
    34511 => -10,
    34512 => -10,
    34513 => -10,
    34514 => -10,
    34515 => -11,
    34516 => -11,
    34517 => -11,
    34518 => -11,
    34519 => -11,
    34520 => -11,
    34521 => -11,
    34522 => -11,
    34523 => -11,
    34524 => -11,
    34525 => -11,
    34526 => -11,
    34527 => -11,
    34528 => -11,
    34529 => -11,
    34530 => -11,
    34531 => -11,
    34532 => -11,
    34533 => -11,
    34534 => -11,
    34535 => -11,
    34536 => -11,
    34537 => -11,
    34538 => -11,
    34539 => -11,
    34540 => -11,
    34541 => -11,
    34542 => -11,
    34543 => -11,
    34544 => -11,
    34545 => -11,
    34546 => -11,
    34547 => -11,
    34548 => -11,
    34549 => -11,
    34550 => -11,
    34551 => -11,
    34552 => -11,
    34553 => -11,
    34554 => -11,
    34555 => -11,
    34556 => -11,
    34557 => -11,
    34558 => -11,
    34559 => -11,
    34560 => -11,
    34561 => -11,
    34562 => -11,
    34563 => -11,
    34564 => -11,
    34565 => -11,
    34566 => -11,
    34567 => -11,
    34568 => -11,
    34569 => -11,
    34570 => -11,
    34571 => -11,
    34572 => -11,
    34573 => -11,
    34574 => -11,
    34575 => -11,
    34576 => -11,
    34577 => -11,
    34578 => -11,
    34579 => -11,
    34580 => -11,
    34581 => -11,
    34582 => -11,
    34583 => -11,
    34584 => -11,
    34585 => -11,
    34586 => -11,
    34587 => -11,
    34588 => -11,
    34589 => -11,
    34590 => -11,
    34591 => -11,
    34592 => -11,
    34593 => -11,
    34594 => -11,
    34595 => -11,
    34596 => -11,
    34597 => -11,
    34598 => -11,
    34599 => -11,
    34600 => -11,
    34601 => -11,
    34602 => -11,
    34603 => -11,
    34604 => -11,
    34605 => -11,
    34606 => -11,
    34607 => -11,
    34608 => -11,
    34609 => -11,
    34610 => -11,
    34611 => -11,
    34612 => -11,
    34613 => -11,
    34614 => -11,
    34615 => -11,
    34616 => -11,
    34617 => -11,
    34618 => -11,
    34619 => -11,
    34620 => -11,
    34621 => -11,
    34622 => -11,
    34623 => -11,
    34624 => -11,
    34625 => -11,
    34626 => -11,
    34627 => -11,
    34628 => -11,
    34629 => -11,
    34630 => -11,
    34631 => -11,
    34632 => -11,
    34633 => -11,
    34634 => -11,
    34635 => -11,
    34636 => -11,
    34637 => -11,
    34638 => -11,
    34639 => -11,
    34640 => -11,
    34641 => -11,
    34642 => -11,
    34643 => -11,
    34644 => -11,
    34645 => -11,
    34646 => -11,
    34647 => -11,
    34648 => -11,
    34649 => -11,
    34650 => -11,
    34651 => -11,
    34652 => -11,
    34653 => -11,
    34654 => -11,
    34655 => -11,
    34656 => -11,
    34657 => -11,
    34658 => -11,
    34659 => -11,
    34660 => -11,
    34661 => -11,
    34662 => -11,
    34663 => -11,
    34664 => -11,
    34665 => -11,
    34666 => -11,
    34667 => -11,
    34668 => -11,
    34669 => -11,
    34670 => -11,
    34671 => -11,
    34672 => -11,
    34673 => -11,
    34674 => -11,
    34675 => -11,
    34676 => -11,
    34677 => -11,
    34678 => -11,
    34679 => -11,
    34680 => -11,
    34681 => -11,
    34682 => -11,
    34683 => -12,
    34684 => -12,
    34685 => -12,
    34686 => -12,
    34687 => -12,
    34688 => -12,
    34689 => -12,
    34690 => -12,
    34691 => -12,
    34692 => -12,
    34693 => -12,
    34694 => -12,
    34695 => -12,
    34696 => -12,
    34697 => -12,
    34698 => -12,
    34699 => -12,
    34700 => -12,
    34701 => -12,
    34702 => -12,
    34703 => -12,
    34704 => -12,
    34705 => -12,
    34706 => -12,
    34707 => -12,
    34708 => -12,
    34709 => -12,
    34710 => -12,
    34711 => -12,
    34712 => -12,
    34713 => -12,
    34714 => -12,
    34715 => -12,
    34716 => -12,
    34717 => -12,
    34718 => -12,
    34719 => -12,
    34720 => -12,
    34721 => -12,
    34722 => -12,
    34723 => -12,
    34724 => -12,
    34725 => -12,
    34726 => -12,
    34727 => -12,
    34728 => -12,
    34729 => -12,
    34730 => -12,
    34731 => -12,
    34732 => -12,
    34733 => -12,
    34734 => -12,
    34735 => -12,
    34736 => -12,
    34737 => -12,
    34738 => -12,
    34739 => -12,
    34740 => -12,
    34741 => -12,
    34742 => -12,
    34743 => -12,
    34744 => -12,
    34745 => -12,
    34746 => -12,
    34747 => -12,
    34748 => -12,
    34749 => -12,
    34750 => -12,
    34751 => -12,
    34752 => -12,
    34753 => -12,
    34754 => -12,
    34755 => -12,
    34756 => -12,
    34757 => -12,
    34758 => -12,
    34759 => -12,
    34760 => -12,
    34761 => -12,
    34762 => -12,
    34763 => -12,
    34764 => -12,
    34765 => -12,
    34766 => -12,
    34767 => -12,
    34768 => -12,
    34769 => -12,
    34770 => -12,
    34771 => -12,
    34772 => -12,
    34773 => -12,
    34774 => -12,
    34775 => -12,
    34776 => -12,
    34777 => -12,
    34778 => -12,
    34779 => -12,
    34780 => -12,
    34781 => -12,
    34782 => -12,
    34783 => -12,
    34784 => -12,
    34785 => -12,
    34786 => -12,
    34787 => -12,
    34788 => -12,
    34789 => -12,
    34790 => -12,
    34791 => -12,
    34792 => -12,
    34793 => -12,
    34794 => -12,
    34795 => -12,
    34796 => -12,
    34797 => -12,
    34798 => -12,
    34799 => -12,
    34800 => -12,
    34801 => -12,
    34802 => -12,
    34803 => -12,
    34804 => -12,
    34805 => -12,
    34806 => -12,
    34807 => -12,
    34808 => -12,
    34809 => -12,
    34810 => -12,
    34811 => -12,
    34812 => -12,
    34813 => -12,
    34814 => -12,
    34815 => -12,
    34816 => -12,
    34817 => -12,
    34818 => -12,
    34819 => -12,
    34820 => -12,
    34821 => -12,
    34822 => -12,
    34823 => -12,
    34824 => -12,
    34825 => -12,
    34826 => -12,
    34827 => -12,
    34828 => -12,
    34829 => -12,
    34830 => -12,
    34831 => -12,
    34832 => -12,
    34833 => -12,
    34834 => -12,
    34835 => -12,
    34836 => -12,
    34837 => -12,
    34838 => -12,
    34839 => -12,
    34840 => -12,
    34841 => -12,
    34842 => -12,
    34843 => -12,
    34844 => -12,
    34845 => -12,
    34846 => -12,
    34847 => -12,
    34848 => -12,
    34849 => -12,
    34850 => -12,
    34851 => -12,
    34852 => -13,
    34853 => -13,
    34854 => -13,
    34855 => -13,
    34856 => -13,
    34857 => -13,
    34858 => -13,
    34859 => -13,
    34860 => -13,
    34861 => -13,
    34862 => -13,
    34863 => -13,
    34864 => -13,
    34865 => -13,
    34866 => -13,
    34867 => -13,
    34868 => -13,
    34869 => -13,
    34870 => -13,
    34871 => -13,
    34872 => -13,
    34873 => -13,
    34874 => -13,
    34875 => -13,
    34876 => -13,
    34877 => -13,
    34878 => -13,
    34879 => -13,
    34880 => -13,
    34881 => -13,
    34882 => -13,
    34883 => -13,
    34884 => -13,
    34885 => -13,
    34886 => -13,
    34887 => -13,
    34888 => -13,
    34889 => -13,
    34890 => -13,
    34891 => -13,
    34892 => -13,
    34893 => -13,
    34894 => -13,
    34895 => -13,
    34896 => -13,
    34897 => -13,
    34898 => -13,
    34899 => -13,
    34900 => -13,
    34901 => -13,
    34902 => -13,
    34903 => -13,
    34904 => -13,
    34905 => -13,
    34906 => -13,
    34907 => -13,
    34908 => -13,
    34909 => -13,
    34910 => -13,
    34911 => -13,
    34912 => -13,
    34913 => -13,
    34914 => -13,
    34915 => -13,
    34916 => -13,
    34917 => -13,
    34918 => -13,
    34919 => -13,
    34920 => -13,
    34921 => -13,
    34922 => -13,
    34923 => -13,
    34924 => -13,
    34925 => -13,
    34926 => -13,
    34927 => -13,
    34928 => -13,
    34929 => -13,
    34930 => -13,
    34931 => -13,
    34932 => -13,
    34933 => -13,
    34934 => -13,
    34935 => -13,
    34936 => -13,
    34937 => -13,
    34938 => -13,
    34939 => -13,
    34940 => -13,
    34941 => -13,
    34942 => -13,
    34943 => -13,
    34944 => -13,
    34945 => -13,
    34946 => -13,
    34947 => -13,
    34948 => -13,
    34949 => -13,
    34950 => -13,
    34951 => -13,
    34952 => -13,
    34953 => -13,
    34954 => -13,
    34955 => -13,
    34956 => -13,
    34957 => -13,
    34958 => -13,
    34959 => -13,
    34960 => -13,
    34961 => -13,
    34962 => -13,
    34963 => -13,
    34964 => -13,
    34965 => -13,
    34966 => -13,
    34967 => -13,
    34968 => -13,
    34969 => -13,
    34970 => -13,
    34971 => -13,
    34972 => -13,
    34973 => -13,
    34974 => -13,
    34975 => -13,
    34976 => -13,
    34977 => -13,
    34978 => -13,
    34979 => -13,
    34980 => -13,
    34981 => -13,
    34982 => -13,
    34983 => -13,
    34984 => -13,
    34985 => -13,
    34986 => -13,
    34987 => -13,
    34988 => -13,
    34989 => -13,
    34990 => -13,
    34991 => -13,
    34992 => -13,
    34993 => -13,
    34994 => -13,
    34995 => -13,
    34996 => -13,
    34997 => -13,
    34998 => -13,
    34999 => -13,
    35000 => -13,
    35001 => -13,
    35002 => -13,
    35003 => -13,
    35004 => -13,
    35005 => -13,
    35006 => -13,
    35007 => -13,
    35008 => -13,
    35009 => -13,
    35010 => -13,
    35011 => -13,
    35012 => -13,
    35013 => -13,
    35014 => -13,
    35015 => -13,
    35016 => -13,
    35017 => -13,
    35018 => -13,
    35019 => -13,
    35020 => -13,
    35021 => -14,
    35022 => -14,
    35023 => -14,
    35024 => -14,
    35025 => -14,
    35026 => -14,
    35027 => -14,
    35028 => -14,
    35029 => -14,
    35030 => -14,
    35031 => -14,
    35032 => -14,
    35033 => -14,
    35034 => -14,
    35035 => -14,
    35036 => -14,
    35037 => -14,
    35038 => -14,
    35039 => -14,
    35040 => -14,
    35041 => -14,
    35042 => -14,
    35043 => -14,
    35044 => -14,
    35045 => -14,
    35046 => -14,
    35047 => -14,
    35048 => -14,
    35049 => -14,
    35050 => -14,
    35051 => -14,
    35052 => -14,
    35053 => -14,
    35054 => -14,
    35055 => -14,
    35056 => -14,
    35057 => -14,
    35058 => -14,
    35059 => -14,
    35060 => -14,
    35061 => -14,
    35062 => -14,
    35063 => -14,
    35064 => -14,
    35065 => -14,
    35066 => -14,
    35067 => -14,
    35068 => -14,
    35069 => -14,
    35070 => -14,
    35071 => -14,
    35072 => -14,
    35073 => -14,
    35074 => -14,
    35075 => -14,
    35076 => -14,
    35077 => -14,
    35078 => -14,
    35079 => -14,
    35080 => -14,
    35081 => -14,
    35082 => -14,
    35083 => -14,
    35084 => -14,
    35085 => -14,
    35086 => -14,
    35087 => -14,
    35088 => -14,
    35089 => -14,
    35090 => -14,
    35091 => -14,
    35092 => -14,
    35093 => -14,
    35094 => -14,
    35095 => -14,
    35096 => -14,
    35097 => -14,
    35098 => -14,
    35099 => -14,
    35100 => -14,
    35101 => -14,
    35102 => -14,
    35103 => -14,
    35104 => -14,
    35105 => -14,
    35106 => -14,
    35107 => -14,
    35108 => -14,
    35109 => -14,
    35110 => -14,
    35111 => -14,
    35112 => -14,
    35113 => -14,
    35114 => -14,
    35115 => -14,
    35116 => -14,
    35117 => -14,
    35118 => -14,
    35119 => -14,
    35120 => -14,
    35121 => -14,
    35122 => -14,
    35123 => -14,
    35124 => -14,
    35125 => -14,
    35126 => -14,
    35127 => -14,
    35128 => -14,
    35129 => -14,
    35130 => -14,
    35131 => -14,
    35132 => -14,
    35133 => -14,
    35134 => -14,
    35135 => -14,
    35136 => -14,
    35137 => -14,
    35138 => -14,
    35139 => -14,
    35140 => -14,
    35141 => -14,
    35142 => -14,
    35143 => -14,
    35144 => -14,
    35145 => -14,
    35146 => -14,
    35147 => -14,
    35148 => -14,
    35149 => -14,
    35150 => -14,
    35151 => -14,
    35152 => -14,
    35153 => -14,
    35154 => -14,
    35155 => -14,
    35156 => -14,
    35157 => -14,
    35158 => -14,
    35159 => -14,
    35160 => -14,
    35161 => -14,
    35162 => -14,
    35163 => -14,
    35164 => -14,
    35165 => -14,
    35166 => -14,
    35167 => -14,
    35168 => -14,
    35169 => -14,
    35170 => -14,
    35171 => -14,
    35172 => -14,
    35173 => -14,
    35174 => -14,
    35175 => -14,
    35176 => -14,
    35177 => -14,
    35178 => -14,
    35179 => -14,
    35180 => -14,
    35181 => -14,
    35182 => -14,
    35183 => -14,
    35184 => -14,
    35185 => -14,
    35186 => -14,
    35187 => -14,
    35188 => -14,
    35189 => -14,
    35190 => -14,
    35191 => -15,
    35192 => -15,
    35193 => -15,
    35194 => -15,
    35195 => -15,
    35196 => -15,
    35197 => -15,
    35198 => -15,
    35199 => -15,
    35200 => -15,
    35201 => -15,
    35202 => -15,
    35203 => -15,
    35204 => -15,
    35205 => -15,
    35206 => -15,
    35207 => -15,
    35208 => -15,
    35209 => -15,
    35210 => -15,
    35211 => -15,
    35212 => -15,
    35213 => -15,
    35214 => -15,
    35215 => -15,
    35216 => -15,
    35217 => -15,
    35218 => -15,
    35219 => -15,
    35220 => -15,
    35221 => -15,
    35222 => -15,
    35223 => -15,
    35224 => -15,
    35225 => -15,
    35226 => -15,
    35227 => -15,
    35228 => -15,
    35229 => -15,
    35230 => -15,
    35231 => -15,
    35232 => -15,
    35233 => -15,
    35234 => -15,
    35235 => -15,
    35236 => -15,
    35237 => -15,
    35238 => -15,
    35239 => -15,
    35240 => -15,
    35241 => -15,
    35242 => -15,
    35243 => -15,
    35244 => -15,
    35245 => -15,
    35246 => -15,
    35247 => -15,
    35248 => -15,
    35249 => -15,
    35250 => -15,
    35251 => -15,
    35252 => -15,
    35253 => -15,
    35254 => -15,
    35255 => -15,
    35256 => -15,
    35257 => -15,
    35258 => -15,
    35259 => -15,
    35260 => -15,
    35261 => -15,
    35262 => -15,
    35263 => -15,
    35264 => -15,
    35265 => -15,
    35266 => -15,
    35267 => -15,
    35268 => -15,
    35269 => -15,
    35270 => -15,
    35271 => -15,
    35272 => -15,
    35273 => -15,
    35274 => -15,
    35275 => -15,
    35276 => -15,
    35277 => -15,
    35278 => -15,
    35279 => -15,
    35280 => -15,
    35281 => -15,
    35282 => -15,
    35283 => -15,
    35284 => -15,
    35285 => -15,
    35286 => -15,
    35287 => -15,
    35288 => -15,
    35289 => -15,
    35290 => -15,
    35291 => -15,
    35292 => -15,
    35293 => -15,
    35294 => -15,
    35295 => -15,
    35296 => -15,
    35297 => -15,
    35298 => -15,
    35299 => -15,
    35300 => -15,
    35301 => -15,
    35302 => -15,
    35303 => -15,
    35304 => -15,
    35305 => -15,
    35306 => -15,
    35307 => -15,
    35308 => -15,
    35309 => -15,
    35310 => -15,
    35311 => -15,
    35312 => -15,
    35313 => -15,
    35314 => -15,
    35315 => -15,
    35316 => -15,
    35317 => -15,
    35318 => -15,
    35319 => -15,
    35320 => -15,
    35321 => -15,
    35322 => -15,
    35323 => -15,
    35324 => -15,
    35325 => -15,
    35326 => -15,
    35327 => -15,
    35328 => -15,
    35329 => -15,
    35330 => -15,
    35331 => -15,
    35332 => -15,
    35333 => -15,
    35334 => -15,
    35335 => -15,
    35336 => -15,
    35337 => -15,
    35338 => -15,
    35339 => -15,
    35340 => -15,
    35341 => -15,
    35342 => -15,
    35343 => -15,
    35344 => -15,
    35345 => -15,
    35346 => -15,
    35347 => -15,
    35348 => -15,
    35349 => -15,
    35350 => -15,
    35351 => -15,
    35352 => -15,
    35353 => -15,
    35354 => -15,
    35355 => -15,
    35356 => -15,
    35357 => -15,
    35358 => -15,
    35359 => -15,
    35360 => -15,
    35361 => -16,
    35362 => -16,
    35363 => -16,
    35364 => -16,
    35365 => -16,
    35366 => -16,
    35367 => -16,
    35368 => -16,
    35369 => -16,
    35370 => -16,
    35371 => -16,
    35372 => -16,
    35373 => -16,
    35374 => -16,
    35375 => -16,
    35376 => -16,
    35377 => -16,
    35378 => -16,
    35379 => -16,
    35380 => -16,
    35381 => -16,
    35382 => -16,
    35383 => -16,
    35384 => -16,
    35385 => -16,
    35386 => -16,
    35387 => -16,
    35388 => -16,
    35389 => -16,
    35390 => -16,
    35391 => -16,
    35392 => -16,
    35393 => -16,
    35394 => -16,
    35395 => -16,
    35396 => -16,
    35397 => -16,
    35398 => -16,
    35399 => -16,
    35400 => -16,
    35401 => -16,
    35402 => -16,
    35403 => -16,
    35404 => -16,
    35405 => -16,
    35406 => -16,
    35407 => -16,
    35408 => -16,
    35409 => -16,
    35410 => -16,
    35411 => -16,
    35412 => -16,
    35413 => -16,
    35414 => -16,
    35415 => -16,
    35416 => -16,
    35417 => -16,
    35418 => -16,
    35419 => -16,
    35420 => -16,
    35421 => -16,
    35422 => -16,
    35423 => -16,
    35424 => -16,
    35425 => -16,
    35426 => -16,
    35427 => -16,
    35428 => -16,
    35429 => -16,
    35430 => -16,
    35431 => -16,
    35432 => -16,
    35433 => -16,
    35434 => -16,
    35435 => -16,
    35436 => -16,
    35437 => -16,
    35438 => -16,
    35439 => -16,
    35440 => -16,
    35441 => -16,
    35442 => -16,
    35443 => -16,
    35444 => -16,
    35445 => -16,
    35446 => -16,
    35447 => -16,
    35448 => -16,
    35449 => -16,
    35450 => -16,
    35451 => -16,
    35452 => -16,
    35453 => -16,
    35454 => -16,
    35455 => -16,
    35456 => -16,
    35457 => -16,
    35458 => -16,
    35459 => -16,
    35460 => -16,
    35461 => -16,
    35462 => -16,
    35463 => -16,
    35464 => -16,
    35465 => -16,
    35466 => -16,
    35467 => -16,
    35468 => -16,
    35469 => -16,
    35470 => -16,
    35471 => -16,
    35472 => -16,
    35473 => -16,
    35474 => -16,
    35475 => -16,
    35476 => -16,
    35477 => -16,
    35478 => -16,
    35479 => -16,
    35480 => -16,
    35481 => -16,
    35482 => -16,
    35483 => -16,
    35484 => -16,
    35485 => -16,
    35486 => -16,
    35487 => -16,
    35488 => -16,
    35489 => -16,
    35490 => -16,
    35491 => -16,
    35492 => -16,
    35493 => -16,
    35494 => -16,
    35495 => -16,
    35496 => -16,
    35497 => -16,
    35498 => -16,
    35499 => -16,
    35500 => -16,
    35501 => -16,
    35502 => -16,
    35503 => -16,
    35504 => -16,
    35505 => -16,
    35506 => -16,
    35507 => -16,
    35508 => -16,
    35509 => -16,
    35510 => -16,
    35511 => -16,
    35512 => -16,
    35513 => -16,
    35514 => -16,
    35515 => -16,
    35516 => -16,
    35517 => -16,
    35518 => -16,
    35519 => -16,
    35520 => -16,
    35521 => -16,
    35522 => -16,
    35523 => -16,
    35524 => -16,
    35525 => -16,
    35526 => -16,
    35527 => -16,
    35528 => -16,
    35529 => -16,
    35530 => -16,
    35531 => -16,
    35532 => -16,
    35533 => -17,
    35534 => -17,
    35535 => -17,
    35536 => -17,
    35537 => -17,
    35538 => -17,
    35539 => -17,
    35540 => -17,
    35541 => -17,
    35542 => -17,
    35543 => -17,
    35544 => -17,
    35545 => -17,
    35546 => -17,
    35547 => -17,
    35548 => -17,
    35549 => -17,
    35550 => -17,
    35551 => -17,
    35552 => -17,
    35553 => -17,
    35554 => -17,
    35555 => -17,
    35556 => -17,
    35557 => -17,
    35558 => -17,
    35559 => -17,
    35560 => -17,
    35561 => -17,
    35562 => -17,
    35563 => -17,
    35564 => -17,
    35565 => -17,
    35566 => -17,
    35567 => -17,
    35568 => -17,
    35569 => -17,
    35570 => -17,
    35571 => -17,
    35572 => -17,
    35573 => -17,
    35574 => -17,
    35575 => -17,
    35576 => -17,
    35577 => -17,
    35578 => -17,
    35579 => -17,
    35580 => -17,
    35581 => -17,
    35582 => -17,
    35583 => -17,
    35584 => -17,
    35585 => -17,
    35586 => -17,
    35587 => -17,
    35588 => -17,
    35589 => -17,
    35590 => -17,
    35591 => -17,
    35592 => -17,
    35593 => -17,
    35594 => -17,
    35595 => -17,
    35596 => -17,
    35597 => -17,
    35598 => -17,
    35599 => -17,
    35600 => -17,
    35601 => -17,
    35602 => -17,
    35603 => -17,
    35604 => -17,
    35605 => -17,
    35606 => -17,
    35607 => -17,
    35608 => -17,
    35609 => -17,
    35610 => -17,
    35611 => -17,
    35612 => -17,
    35613 => -17,
    35614 => -17,
    35615 => -17,
    35616 => -17,
    35617 => -17,
    35618 => -17,
    35619 => -17,
    35620 => -17,
    35621 => -17,
    35622 => -17,
    35623 => -17,
    35624 => -17,
    35625 => -17,
    35626 => -17,
    35627 => -17,
    35628 => -17,
    35629 => -17,
    35630 => -17,
    35631 => -17,
    35632 => -17,
    35633 => -17,
    35634 => -17,
    35635 => -17,
    35636 => -17,
    35637 => -17,
    35638 => -17,
    35639 => -17,
    35640 => -17,
    35641 => -17,
    35642 => -17,
    35643 => -17,
    35644 => -17,
    35645 => -17,
    35646 => -17,
    35647 => -17,
    35648 => -17,
    35649 => -17,
    35650 => -17,
    35651 => -17,
    35652 => -17,
    35653 => -17,
    35654 => -17,
    35655 => -17,
    35656 => -17,
    35657 => -17,
    35658 => -17,
    35659 => -17,
    35660 => -17,
    35661 => -17,
    35662 => -17,
    35663 => -17,
    35664 => -17,
    35665 => -17,
    35666 => -17,
    35667 => -17,
    35668 => -17,
    35669 => -17,
    35670 => -17,
    35671 => -17,
    35672 => -17,
    35673 => -17,
    35674 => -17,
    35675 => -17,
    35676 => -17,
    35677 => -17,
    35678 => -17,
    35679 => -17,
    35680 => -17,
    35681 => -17,
    35682 => -17,
    35683 => -17,
    35684 => -17,
    35685 => -17,
    35686 => -17,
    35687 => -17,
    35688 => -17,
    35689 => -17,
    35690 => -17,
    35691 => -17,
    35692 => -17,
    35693 => -17,
    35694 => -17,
    35695 => -17,
    35696 => -17,
    35697 => -17,
    35698 => -17,
    35699 => -17,
    35700 => -17,
    35701 => -17,
    35702 => -17,
    35703 => -17,
    35704 => -18,
    35705 => -18,
    35706 => -18,
    35707 => -18,
    35708 => -18,
    35709 => -18,
    35710 => -18,
    35711 => -18,
    35712 => -18,
    35713 => -18,
    35714 => -18,
    35715 => -18,
    35716 => -18,
    35717 => -18,
    35718 => -18,
    35719 => -18,
    35720 => -18,
    35721 => -18,
    35722 => -18,
    35723 => -18,
    35724 => -18,
    35725 => -18,
    35726 => -18,
    35727 => -18,
    35728 => -18,
    35729 => -18,
    35730 => -18,
    35731 => -18,
    35732 => -18,
    35733 => -18,
    35734 => -18,
    35735 => -18,
    35736 => -18,
    35737 => -18,
    35738 => -18,
    35739 => -18,
    35740 => -18,
    35741 => -18,
    35742 => -18,
    35743 => -18,
    35744 => -18,
    35745 => -18,
    35746 => -18,
    35747 => -18,
    35748 => -18,
    35749 => -18,
    35750 => -18,
    35751 => -18,
    35752 => -18,
    35753 => -18,
    35754 => -18,
    35755 => -18,
    35756 => -18,
    35757 => -18,
    35758 => -18,
    35759 => -18,
    35760 => -18,
    35761 => -18,
    35762 => -18,
    35763 => -18,
    35764 => -18,
    35765 => -18,
    35766 => -18,
    35767 => -18,
    35768 => -18,
    35769 => -18,
    35770 => -18,
    35771 => -18,
    35772 => -18,
    35773 => -18,
    35774 => -18,
    35775 => -18,
    35776 => -18,
    35777 => -18,
    35778 => -18,
    35779 => -18,
    35780 => -18,
    35781 => -18,
    35782 => -18,
    35783 => -18,
    35784 => -18,
    35785 => -18,
    35786 => -18,
    35787 => -18,
    35788 => -18,
    35789 => -18,
    35790 => -18,
    35791 => -18,
    35792 => -18,
    35793 => -18,
    35794 => -18,
    35795 => -18,
    35796 => -18,
    35797 => -18,
    35798 => -18,
    35799 => -18,
    35800 => -18,
    35801 => -18,
    35802 => -18,
    35803 => -18,
    35804 => -18,
    35805 => -18,
    35806 => -18,
    35807 => -18,
    35808 => -18,
    35809 => -18,
    35810 => -18,
    35811 => -18,
    35812 => -18,
    35813 => -18,
    35814 => -18,
    35815 => -18,
    35816 => -18,
    35817 => -18,
    35818 => -18,
    35819 => -18,
    35820 => -18,
    35821 => -18,
    35822 => -18,
    35823 => -18,
    35824 => -18,
    35825 => -18,
    35826 => -18,
    35827 => -18,
    35828 => -18,
    35829 => -18,
    35830 => -18,
    35831 => -18,
    35832 => -18,
    35833 => -18,
    35834 => -18,
    35835 => -18,
    35836 => -18,
    35837 => -18,
    35838 => -18,
    35839 => -18,
    35840 => -18,
    35841 => -18,
    35842 => -18,
    35843 => -18,
    35844 => -18,
    35845 => -18,
    35846 => -18,
    35847 => -18,
    35848 => -18,
    35849 => -18,
    35850 => -18,
    35851 => -18,
    35852 => -18,
    35853 => -18,
    35854 => -18,
    35855 => -18,
    35856 => -18,
    35857 => -18,
    35858 => -18,
    35859 => -18,
    35860 => -18,
    35861 => -18,
    35862 => -18,
    35863 => -18,
    35864 => -18,
    35865 => -18,
    35866 => -18,
    35867 => -18,
    35868 => -18,
    35869 => -18,
    35870 => -18,
    35871 => -18,
    35872 => -18,
    35873 => -18,
    35874 => -18,
    35875 => -18,
    35876 => -18,
    35877 => -19,
    35878 => -19,
    35879 => -19,
    35880 => -19,
    35881 => -19,
    35882 => -19,
    35883 => -19,
    35884 => -19,
    35885 => -19,
    35886 => -19,
    35887 => -19,
    35888 => -19,
    35889 => -19,
    35890 => -19,
    35891 => -19,
    35892 => -19,
    35893 => -19,
    35894 => -19,
    35895 => -19,
    35896 => -19,
    35897 => -19,
    35898 => -19,
    35899 => -19,
    35900 => -19,
    35901 => -19,
    35902 => -19,
    35903 => -19,
    35904 => -19,
    35905 => -19,
    35906 => -19,
    35907 => -19,
    35908 => -19,
    35909 => -19,
    35910 => -19,
    35911 => -19,
    35912 => -19,
    35913 => -19,
    35914 => -19,
    35915 => -19,
    35916 => -19,
    35917 => -19,
    35918 => -19,
    35919 => -19,
    35920 => -19,
    35921 => -19,
    35922 => -19,
    35923 => -19,
    35924 => -19,
    35925 => -19,
    35926 => -19,
    35927 => -19,
    35928 => -19,
    35929 => -19,
    35930 => -19,
    35931 => -19,
    35932 => -19,
    35933 => -19,
    35934 => -19,
    35935 => -19,
    35936 => -19,
    35937 => -19,
    35938 => -19,
    35939 => -19,
    35940 => -19,
    35941 => -19,
    35942 => -19,
    35943 => -19,
    35944 => -19,
    35945 => -19,
    35946 => -19,
    35947 => -19,
    35948 => -19,
    35949 => -19,
    35950 => -19,
    35951 => -19,
    35952 => -19,
    35953 => -19,
    35954 => -19,
    35955 => -19,
    35956 => -19,
    35957 => -19,
    35958 => -19,
    35959 => -19,
    35960 => -19,
    35961 => -19,
    35962 => -19,
    35963 => -19,
    35964 => -19,
    35965 => -19,
    35966 => -19,
    35967 => -19,
    35968 => -19,
    35969 => -19,
    35970 => -19,
    35971 => -19,
    35972 => -19,
    35973 => -19,
    35974 => -19,
    35975 => -19,
    35976 => -19,
    35977 => -19,
    35978 => -19,
    35979 => -19,
    35980 => -19,
    35981 => -19,
    35982 => -19,
    35983 => -19,
    35984 => -19,
    35985 => -19,
    35986 => -19,
    35987 => -19,
    35988 => -19,
    35989 => -19,
    35990 => -19,
    35991 => -19,
    35992 => -19,
    35993 => -19,
    35994 => -19,
    35995 => -19,
    35996 => -19,
    35997 => -19,
    35998 => -19,
    35999 => -19,
    36000 => -19,
    36001 => -19,
    36002 => -19,
    36003 => -19,
    36004 => -19,
    36005 => -19,
    36006 => -19,
    36007 => -19,
    36008 => -19,
    36009 => -19,
    36010 => -19,
    36011 => -19,
    36012 => -19,
    36013 => -19,
    36014 => -19,
    36015 => -19,
    36016 => -19,
    36017 => -19,
    36018 => -19,
    36019 => -19,
    36020 => -19,
    36021 => -19,
    36022 => -19,
    36023 => -19,
    36024 => -19,
    36025 => -19,
    36026 => -19,
    36027 => -19,
    36028 => -19,
    36029 => -19,
    36030 => -19,
    36031 => -19,
    36032 => -19,
    36033 => -19,
    36034 => -19,
    36035 => -19,
    36036 => -19,
    36037 => -19,
    36038 => -19,
    36039 => -19,
    36040 => -19,
    36041 => -19,
    36042 => -19,
    36043 => -19,
    36044 => -19,
    36045 => -19,
    36046 => -19,
    36047 => -19,
    36048 => -19,
    36049 => -19,
    36050 => -19,
    36051 => -20,
    36052 => -20,
    36053 => -20,
    36054 => -20,
    36055 => -20,
    36056 => -20,
    36057 => -20,
    36058 => -20,
    36059 => -20,
    36060 => -20,
    36061 => -20,
    36062 => -20,
    36063 => -20,
    36064 => -20,
    36065 => -20,
    36066 => -20,
    36067 => -20,
    36068 => -20,
    36069 => -20,
    36070 => -20,
    36071 => -20,
    36072 => -20,
    36073 => -20,
    36074 => -20,
    36075 => -20,
    36076 => -20,
    36077 => -20,
    36078 => -20,
    36079 => -20,
    36080 => -20,
    36081 => -20,
    36082 => -20,
    36083 => -20,
    36084 => -20,
    36085 => -20,
    36086 => -20,
    36087 => -20,
    36088 => -20,
    36089 => -20,
    36090 => -20,
    36091 => -20,
    36092 => -20,
    36093 => -20,
    36094 => -20,
    36095 => -20,
    36096 => -20,
    36097 => -20,
    36098 => -20,
    36099 => -20,
    36100 => -20,
    36101 => -20,
    36102 => -20,
    36103 => -20,
    36104 => -20,
    36105 => -20,
    36106 => -20,
    36107 => -20,
    36108 => -20,
    36109 => -20,
    36110 => -20,
    36111 => -20,
    36112 => -20,
    36113 => -20,
    36114 => -20,
    36115 => -20,
    36116 => -20,
    36117 => -20,
    36118 => -20,
    36119 => -20,
    36120 => -20,
    36121 => -20,
    36122 => -20,
    36123 => -20,
    36124 => -20,
    36125 => -20,
    36126 => -20,
    36127 => -20,
    36128 => -20,
    36129 => -20,
    36130 => -20,
    36131 => -20,
    36132 => -20,
    36133 => -20,
    36134 => -20,
    36135 => -20,
    36136 => -20,
    36137 => -20,
    36138 => -20,
    36139 => -20,
    36140 => -20,
    36141 => -20,
    36142 => -20,
    36143 => -20,
    36144 => -20,
    36145 => -20,
    36146 => -20,
    36147 => -20,
    36148 => -20,
    36149 => -20,
    36150 => -20,
    36151 => -20,
    36152 => -20,
    36153 => -20,
    36154 => -20,
    36155 => -20,
    36156 => -20,
    36157 => -20,
    36158 => -20,
    36159 => -20,
    36160 => -20,
    36161 => -20,
    36162 => -20,
    36163 => -20,
    36164 => -20,
    36165 => -20,
    36166 => -20,
    36167 => -20,
    36168 => -20,
    36169 => -20,
    36170 => -20,
    36171 => -20,
    36172 => -20,
    36173 => -20,
    36174 => -20,
    36175 => -20,
    36176 => -20,
    36177 => -20,
    36178 => -20,
    36179 => -20,
    36180 => -20,
    36181 => -20,
    36182 => -20,
    36183 => -20,
    36184 => -20,
    36185 => -20,
    36186 => -20,
    36187 => -20,
    36188 => -20,
    36189 => -20,
    36190 => -20,
    36191 => -20,
    36192 => -20,
    36193 => -20,
    36194 => -20,
    36195 => -20,
    36196 => -20,
    36197 => -20,
    36198 => -20,
    36199 => -20,
    36200 => -20,
    36201 => -20,
    36202 => -20,
    36203 => -20,
    36204 => -20,
    36205 => -20,
    36206 => -20,
    36207 => -20,
    36208 => -20,
    36209 => -20,
    36210 => -20,
    36211 => -20,
    36212 => -20,
    36213 => -20,
    36214 => -20,
    36215 => -20,
    36216 => -20,
    36217 => -20,
    36218 => -20,
    36219 => -20,
    36220 => -20,
    36221 => -20,
    36222 => -20,
    36223 => -20,
    36224 => -20,
    36225 => -21,
    36226 => -21,
    36227 => -21,
    36228 => -21,
    36229 => -21,
    36230 => -21,
    36231 => -21,
    36232 => -21,
    36233 => -21,
    36234 => -21,
    36235 => -21,
    36236 => -21,
    36237 => -21,
    36238 => -21,
    36239 => -21,
    36240 => -21,
    36241 => -21,
    36242 => -21,
    36243 => -21,
    36244 => -21,
    36245 => -21,
    36246 => -21,
    36247 => -21,
    36248 => -21,
    36249 => -21,
    36250 => -21,
    36251 => -21,
    36252 => -21,
    36253 => -21,
    36254 => -21,
    36255 => -21,
    36256 => -21,
    36257 => -21,
    36258 => -21,
    36259 => -21,
    36260 => -21,
    36261 => -21,
    36262 => -21,
    36263 => -21,
    36264 => -21,
    36265 => -21,
    36266 => -21,
    36267 => -21,
    36268 => -21,
    36269 => -21,
    36270 => -21,
    36271 => -21,
    36272 => -21,
    36273 => -21,
    36274 => -21,
    36275 => -21,
    36276 => -21,
    36277 => -21,
    36278 => -21,
    36279 => -21,
    36280 => -21,
    36281 => -21,
    36282 => -21,
    36283 => -21,
    36284 => -21,
    36285 => -21,
    36286 => -21,
    36287 => -21,
    36288 => -21,
    36289 => -21,
    36290 => -21,
    36291 => -21,
    36292 => -21,
    36293 => -21,
    36294 => -21,
    36295 => -21,
    36296 => -21,
    36297 => -21,
    36298 => -21,
    36299 => -21,
    36300 => -21,
    36301 => -21,
    36302 => -21,
    36303 => -21,
    36304 => -21,
    36305 => -21,
    36306 => -21,
    36307 => -21,
    36308 => -21,
    36309 => -21,
    36310 => -21,
    36311 => -21,
    36312 => -21,
    36313 => -21,
    36314 => -21,
    36315 => -21,
    36316 => -21,
    36317 => -21,
    36318 => -21,
    36319 => -21,
    36320 => -21,
    36321 => -21,
    36322 => -21,
    36323 => -21,
    36324 => -21,
    36325 => -21,
    36326 => -21,
    36327 => -21,
    36328 => -21,
    36329 => -21,
    36330 => -21,
    36331 => -21,
    36332 => -21,
    36333 => -21,
    36334 => -21,
    36335 => -21,
    36336 => -21,
    36337 => -21,
    36338 => -21,
    36339 => -21,
    36340 => -21,
    36341 => -21,
    36342 => -21,
    36343 => -21,
    36344 => -21,
    36345 => -21,
    36346 => -21,
    36347 => -21,
    36348 => -21,
    36349 => -21,
    36350 => -21,
    36351 => -21,
    36352 => -21,
    36353 => -21,
    36354 => -21,
    36355 => -21,
    36356 => -21,
    36357 => -21,
    36358 => -21,
    36359 => -21,
    36360 => -21,
    36361 => -21,
    36362 => -21,
    36363 => -21,
    36364 => -21,
    36365 => -21,
    36366 => -21,
    36367 => -21,
    36368 => -21,
    36369 => -21,
    36370 => -21,
    36371 => -21,
    36372 => -21,
    36373 => -21,
    36374 => -21,
    36375 => -21,
    36376 => -21,
    36377 => -21,
    36378 => -21,
    36379 => -21,
    36380 => -21,
    36381 => -21,
    36382 => -21,
    36383 => -21,
    36384 => -21,
    36385 => -21,
    36386 => -21,
    36387 => -21,
    36388 => -21,
    36389 => -21,
    36390 => -21,
    36391 => -21,
    36392 => -21,
    36393 => -21,
    36394 => -21,
    36395 => -21,
    36396 => -21,
    36397 => -21,
    36398 => -21,
    36399 => -21,
    36400 => -21,
    36401 => -22,
    36402 => -22,
    36403 => -22,
    36404 => -22,
    36405 => -22,
    36406 => -22,
    36407 => -22,
    36408 => -22,
    36409 => -22,
    36410 => -22,
    36411 => -22,
    36412 => -22,
    36413 => -22,
    36414 => -22,
    36415 => -22,
    36416 => -22,
    36417 => -22,
    36418 => -22,
    36419 => -22,
    36420 => -22,
    36421 => -22,
    36422 => -22,
    36423 => -22,
    36424 => -22,
    36425 => -22,
    36426 => -22,
    36427 => -22,
    36428 => -22,
    36429 => -22,
    36430 => -22,
    36431 => -22,
    36432 => -22,
    36433 => -22,
    36434 => -22,
    36435 => -22,
    36436 => -22,
    36437 => -22,
    36438 => -22,
    36439 => -22,
    36440 => -22,
    36441 => -22,
    36442 => -22,
    36443 => -22,
    36444 => -22,
    36445 => -22,
    36446 => -22,
    36447 => -22,
    36448 => -22,
    36449 => -22,
    36450 => -22,
    36451 => -22,
    36452 => -22,
    36453 => -22,
    36454 => -22,
    36455 => -22,
    36456 => -22,
    36457 => -22,
    36458 => -22,
    36459 => -22,
    36460 => -22,
    36461 => -22,
    36462 => -22,
    36463 => -22,
    36464 => -22,
    36465 => -22,
    36466 => -22,
    36467 => -22,
    36468 => -22,
    36469 => -22,
    36470 => -22,
    36471 => -22,
    36472 => -22,
    36473 => -22,
    36474 => -22,
    36475 => -22,
    36476 => -22,
    36477 => -22,
    36478 => -22,
    36479 => -22,
    36480 => -22,
    36481 => -22,
    36482 => -22,
    36483 => -22,
    36484 => -22,
    36485 => -22,
    36486 => -22,
    36487 => -22,
    36488 => -22,
    36489 => -22,
    36490 => -22,
    36491 => -22,
    36492 => -22,
    36493 => -22,
    36494 => -22,
    36495 => -22,
    36496 => -22,
    36497 => -22,
    36498 => -22,
    36499 => -22,
    36500 => -22,
    36501 => -22,
    36502 => -22,
    36503 => -22,
    36504 => -22,
    36505 => -22,
    36506 => -22,
    36507 => -22,
    36508 => -22,
    36509 => -22,
    36510 => -22,
    36511 => -22,
    36512 => -22,
    36513 => -22,
    36514 => -22,
    36515 => -22,
    36516 => -22,
    36517 => -22,
    36518 => -22,
    36519 => -22,
    36520 => -22,
    36521 => -22,
    36522 => -22,
    36523 => -22,
    36524 => -22,
    36525 => -22,
    36526 => -22,
    36527 => -22,
    36528 => -22,
    36529 => -22,
    36530 => -22,
    36531 => -22,
    36532 => -22,
    36533 => -22,
    36534 => -22,
    36535 => -22,
    36536 => -22,
    36537 => -22,
    36538 => -22,
    36539 => -22,
    36540 => -22,
    36541 => -22,
    36542 => -22,
    36543 => -22,
    36544 => -22,
    36545 => -22,
    36546 => -22,
    36547 => -22,
    36548 => -22,
    36549 => -22,
    36550 => -22,
    36551 => -22,
    36552 => -22,
    36553 => -22,
    36554 => -22,
    36555 => -22,
    36556 => -22,
    36557 => -22,
    36558 => -22,
    36559 => -22,
    36560 => -22,
    36561 => -22,
    36562 => -22,
    36563 => -22,
    36564 => -22,
    36565 => -22,
    36566 => -22,
    36567 => -22,
    36568 => -22,
    36569 => -22,
    36570 => -22,
    36571 => -22,
    36572 => -22,
    36573 => -22,
    36574 => -22,
    36575 => -22,
    36576 => -22,
    36577 => -22,
    36578 => -23,
    36579 => -23,
    36580 => -23,
    36581 => -23,
    36582 => -23,
    36583 => -23,
    36584 => -23,
    36585 => -23,
    36586 => -23,
    36587 => -23,
    36588 => -23,
    36589 => -23,
    36590 => -23,
    36591 => -23,
    36592 => -23,
    36593 => -23,
    36594 => -23,
    36595 => -23,
    36596 => -23,
    36597 => -23,
    36598 => -23,
    36599 => -23,
    36600 => -23,
    36601 => -23,
    36602 => -23,
    36603 => -23,
    36604 => -23,
    36605 => -23,
    36606 => -23,
    36607 => -23,
    36608 => -23,
    36609 => -23,
    36610 => -23,
    36611 => -23,
    36612 => -23,
    36613 => -23,
    36614 => -23,
    36615 => -23,
    36616 => -23,
    36617 => -23,
    36618 => -23,
    36619 => -23,
    36620 => -23,
    36621 => -23,
    36622 => -23,
    36623 => -23,
    36624 => -23,
    36625 => -23,
    36626 => -23,
    36627 => -23,
    36628 => -23,
    36629 => -23,
    36630 => -23,
    36631 => -23,
    36632 => -23,
    36633 => -23,
    36634 => -23,
    36635 => -23,
    36636 => -23,
    36637 => -23,
    36638 => -23,
    36639 => -23,
    36640 => -23,
    36641 => -23,
    36642 => -23,
    36643 => -23,
    36644 => -23,
    36645 => -23,
    36646 => -23,
    36647 => -23,
    36648 => -23,
    36649 => -23,
    36650 => -23,
    36651 => -23,
    36652 => -23,
    36653 => -23,
    36654 => -23,
    36655 => -23,
    36656 => -23,
    36657 => -23,
    36658 => -23,
    36659 => -23,
    36660 => -23,
    36661 => -23,
    36662 => -23,
    36663 => -23,
    36664 => -23,
    36665 => -23,
    36666 => -23,
    36667 => -23,
    36668 => -23,
    36669 => -23,
    36670 => -23,
    36671 => -23,
    36672 => -23,
    36673 => -23,
    36674 => -23,
    36675 => -23,
    36676 => -23,
    36677 => -23,
    36678 => -23,
    36679 => -23,
    36680 => -23,
    36681 => -23,
    36682 => -23,
    36683 => -23,
    36684 => -23,
    36685 => -23,
    36686 => -23,
    36687 => -23,
    36688 => -23,
    36689 => -23,
    36690 => -23,
    36691 => -23,
    36692 => -23,
    36693 => -23,
    36694 => -23,
    36695 => -23,
    36696 => -23,
    36697 => -23,
    36698 => -23,
    36699 => -23,
    36700 => -23,
    36701 => -23,
    36702 => -23,
    36703 => -23,
    36704 => -23,
    36705 => -23,
    36706 => -23,
    36707 => -23,
    36708 => -23,
    36709 => -23,
    36710 => -23,
    36711 => -23,
    36712 => -23,
    36713 => -23,
    36714 => -23,
    36715 => -23,
    36716 => -23,
    36717 => -23,
    36718 => -23,
    36719 => -23,
    36720 => -23,
    36721 => -23,
    36722 => -23,
    36723 => -23,
    36724 => -23,
    36725 => -23,
    36726 => -23,
    36727 => -23,
    36728 => -23,
    36729 => -23,
    36730 => -23,
    36731 => -23,
    36732 => -23,
    36733 => -23,
    36734 => -23,
    36735 => -23,
    36736 => -23,
    36737 => -23,
    36738 => -23,
    36739 => -23,
    36740 => -23,
    36741 => -23,
    36742 => -23,
    36743 => -23,
    36744 => -23,
    36745 => -23,
    36746 => -23,
    36747 => -23,
    36748 => -23,
    36749 => -23,
    36750 => -23,
    36751 => -23,
    36752 => -23,
    36753 => -23,
    36754 => -23,
    36755 => -23,
    36756 => -24,
    36757 => -24,
    36758 => -24,
    36759 => -24,
    36760 => -24,
    36761 => -24,
    36762 => -24,
    36763 => -24,
    36764 => -24,
    36765 => -24,
    36766 => -24,
    36767 => -24,
    36768 => -24,
    36769 => -24,
    36770 => -24,
    36771 => -24,
    36772 => -24,
    36773 => -24,
    36774 => -24,
    36775 => -24,
    36776 => -24,
    36777 => -24,
    36778 => -24,
    36779 => -24,
    36780 => -24,
    36781 => -24,
    36782 => -24,
    36783 => -24,
    36784 => -24,
    36785 => -24,
    36786 => -24,
    36787 => -24,
    36788 => -24,
    36789 => -24,
    36790 => -24,
    36791 => -24,
    36792 => -24,
    36793 => -24,
    36794 => -24,
    36795 => -24,
    36796 => -24,
    36797 => -24,
    36798 => -24,
    36799 => -24,
    36800 => -24,
    36801 => -24,
    36802 => -24,
    36803 => -24,
    36804 => -24,
    36805 => -24,
    36806 => -24,
    36807 => -24,
    36808 => -24,
    36809 => -24,
    36810 => -24,
    36811 => -24,
    36812 => -24,
    36813 => -24,
    36814 => -24,
    36815 => -24,
    36816 => -24,
    36817 => -24,
    36818 => -24,
    36819 => -24,
    36820 => -24,
    36821 => -24,
    36822 => -24,
    36823 => -24,
    36824 => -24,
    36825 => -24,
    36826 => -24,
    36827 => -24,
    36828 => -24,
    36829 => -24,
    36830 => -24,
    36831 => -24,
    36832 => -24,
    36833 => -24,
    36834 => -24,
    36835 => -24,
    36836 => -24,
    36837 => -24,
    36838 => -24,
    36839 => -24,
    36840 => -24,
    36841 => -24,
    36842 => -24,
    36843 => -24,
    36844 => -24,
    36845 => -24,
    36846 => -24,
    36847 => -24,
    36848 => -24,
    36849 => -24,
    36850 => -24,
    36851 => -24,
    36852 => -24,
    36853 => -24,
    36854 => -24,
    36855 => -24,
    36856 => -24,
    36857 => -24,
    36858 => -24,
    36859 => -24,
    36860 => -24,
    36861 => -24,
    36862 => -24,
    36863 => -24,
    36864 => -24,
    36865 => -24,
    36866 => -24,
    36867 => -24,
    36868 => -24,
    36869 => -24,
    36870 => -24,
    36871 => -24,
    36872 => -24,
    36873 => -24,
    36874 => -24,
    36875 => -24,
    36876 => -24,
    36877 => -24,
    36878 => -24,
    36879 => -24,
    36880 => -24,
    36881 => -24,
    36882 => -24,
    36883 => -24,
    36884 => -24,
    36885 => -24,
    36886 => -24,
    36887 => -24,
    36888 => -24,
    36889 => -24,
    36890 => -24,
    36891 => -24,
    36892 => -24,
    36893 => -24,
    36894 => -24,
    36895 => -24,
    36896 => -24,
    36897 => -24,
    36898 => -24,
    36899 => -24,
    36900 => -24,
    36901 => -24,
    36902 => -24,
    36903 => -24,
    36904 => -24,
    36905 => -24,
    36906 => -24,
    36907 => -24,
    36908 => -24,
    36909 => -24,
    36910 => -24,
    36911 => -24,
    36912 => -24,
    36913 => -24,
    36914 => -24,
    36915 => -24,
    36916 => -24,
    36917 => -24,
    36918 => -24,
    36919 => -24,
    36920 => -24,
    36921 => -24,
    36922 => -24,
    36923 => -24,
    36924 => -24,
    36925 => -24,
    36926 => -24,
    36927 => -24,
    36928 => -24,
    36929 => -24,
    36930 => -24,
    36931 => -24,
    36932 => -24,
    36933 => -24,
    36934 => -24,
    36935 => -25,
    36936 => -25,
    36937 => -25,
    36938 => -25,
    36939 => -25,
    36940 => -25,
    36941 => -25,
    36942 => -25,
    36943 => -25,
    36944 => -25,
    36945 => -25,
    36946 => -25,
    36947 => -25,
    36948 => -25,
    36949 => -25,
    36950 => -25,
    36951 => -25,
    36952 => -25,
    36953 => -25,
    36954 => -25,
    36955 => -25,
    36956 => -25,
    36957 => -25,
    36958 => -25,
    36959 => -25,
    36960 => -25,
    36961 => -25,
    36962 => -25,
    36963 => -25,
    36964 => -25,
    36965 => -25,
    36966 => -25,
    36967 => -25,
    36968 => -25,
    36969 => -25,
    36970 => -25,
    36971 => -25,
    36972 => -25,
    36973 => -25,
    36974 => -25,
    36975 => -25,
    36976 => -25,
    36977 => -25,
    36978 => -25,
    36979 => -25,
    36980 => -25,
    36981 => -25,
    36982 => -25,
    36983 => -25,
    36984 => -25,
    36985 => -25,
    36986 => -25,
    36987 => -25,
    36988 => -25,
    36989 => -25,
    36990 => -25,
    36991 => -25,
    36992 => -25,
    36993 => -25,
    36994 => -25,
    36995 => -25,
    36996 => -25,
    36997 => -25,
    36998 => -25,
    36999 => -25,
    37000 => -25,
    37001 => -25,
    37002 => -25,
    37003 => -25,
    37004 => -25,
    37005 => -25,
    37006 => -25,
    37007 => -25,
    37008 => -25,
    37009 => -25,
    37010 => -25,
    37011 => -25,
    37012 => -25,
    37013 => -25,
    37014 => -25,
    37015 => -25,
    37016 => -25,
    37017 => -25,
    37018 => -25,
    37019 => -25,
    37020 => -25,
    37021 => -25,
    37022 => -25,
    37023 => -25,
    37024 => -25,
    37025 => -25,
    37026 => -25,
    37027 => -25,
    37028 => -25,
    37029 => -25,
    37030 => -25,
    37031 => -25,
    37032 => -25,
    37033 => -25,
    37034 => -25,
    37035 => -25,
    37036 => -25,
    37037 => -25,
    37038 => -25,
    37039 => -25,
    37040 => -25,
    37041 => -25,
    37042 => -25,
    37043 => -25,
    37044 => -25,
    37045 => -25,
    37046 => -25,
    37047 => -25,
    37048 => -25,
    37049 => -25,
    37050 => -25,
    37051 => -25,
    37052 => -25,
    37053 => -25,
    37054 => -25,
    37055 => -25,
    37056 => -25,
    37057 => -25,
    37058 => -25,
    37059 => -25,
    37060 => -25,
    37061 => -25,
    37062 => -25,
    37063 => -25,
    37064 => -25,
    37065 => -25,
    37066 => -25,
    37067 => -25,
    37068 => -25,
    37069 => -25,
    37070 => -25,
    37071 => -25,
    37072 => -25,
    37073 => -25,
    37074 => -25,
    37075 => -25,
    37076 => -25,
    37077 => -25,
    37078 => -25,
    37079 => -25,
    37080 => -25,
    37081 => -25,
    37082 => -25,
    37083 => -25,
    37084 => -25,
    37085 => -25,
    37086 => -25,
    37087 => -25,
    37088 => -25,
    37089 => -25,
    37090 => -25,
    37091 => -25,
    37092 => -25,
    37093 => -25,
    37094 => -25,
    37095 => -25,
    37096 => -25,
    37097 => -25,
    37098 => -25,
    37099 => -25,
    37100 => -25,
    37101 => -25,
    37102 => -25,
    37103 => -25,
    37104 => -25,
    37105 => -25,
    37106 => -25,
    37107 => -25,
    37108 => -25,
    37109 => -25,
    37110 => -25,
    37111 => -25,
    37112 => -25,
    37113 => -25,
    37114 => -25,
    37115 => -26,
    37116 => -26,
    37117 => -26,
    37118 => -26,
    37119 => -26,
    37120 => -26,
    37121 => -26,
    37122 => -26,
    37123 => -26,
    37124 => -26,
    37125 => -26,
    37126 => -26,
    37127 => -26,
    37128 => -26,
    37129 => -26,
    37130 => -26,
    37131 => -26,
    37132 => -26,
    37133 => -26,
    37134 => -26,
    37135 => -26,
    37136 => -26,
    37137 => -26,
    37138 => -26,
    37139 => -26,
    37140 => -26,
    37141 => -26,
    37142 => -26,
    37143 => -26,
    37144 => -26,
    37145 => -26,
    37146 => -26,
    37147 => -26,
    37148 => -26,
    37149 => -26,
    37150 => -26,
    37151 => -26,
    37152 => -26,
    37153 => -26,
    37154 => -26,
    37155 => -26,
    37156 => -26,
    37157 => -26,
    37158 => -26,
    37159 => -26,
    37160 => -26,
    37161 => -26,
    37162 => -26,
    37163 => -26,
    37164 => -26,
    37165 => -26,
    37166 => -26,
    37167 => -26,
    37168 => -26,
    37169 => -26,
    37170 => -26,
    37171 => -26,
    37172 => -26,
    37173 => -26,
    37174 => -26,
    37175 => -26,
    37176 => -26,
    37177 => -26,
    37178 => -26,
    37179 => -26,
    37180 => -26,
    37181 => -26,
    37182 => -26,
    37183 => -26,
    37184 => -26,
    37185 => -26,
    37186 => -26,
    37187 => -26,
    37188 => -26,
    37189 => -26,
    37190 => -26,
    37191 => -26,
    37192 => -26,
    37193 => -26,
    37194 => -26,
    37195 => -26,
    37196 => -26,
    37197 => -26,
    37198 => -26,
    37199 => -26,
    37200 => -26,
    37201 => -26,
    37202 => -26,
    37203 => -26,
    37204 => -26,
    37205 => -26,
    37206 => -26,
    37207 => -26,
    37208 => -26,
    37209 => -26,
    37210 => -26,
    37211 => -26,
    37212 => -26,
    37213 => -26,
    37214 => -26,
    37215 => -26,
    37216 => -26,
    37217 => -26,
    37218 => -26,
    37219 => -26,
    37220 => -26,
    37221 => -26,
    37222 => -26,
    37223 => -26,
    37224 => -26,
    37225 => -26,
    37226 => -26,
    37227 => -26,
    37228 => -26,
    37229 => -26,
    37230 => -26,
    37231 => -26,
    37232 => -26,
    37233 => -26,
    37234 => -26,
    37235 => -26,
    37236 => -26,
    37237 => -26,
    37238 => -26,
    37239 => -26,
    37240 => -26,
    37241 => -26,
    37242 => -26,
    37243 => -26,
    37244 => -26,
    37245 => -26,
    37246 => -26,
    37247 => -26,
    37248 => -26,
    37249 => -26,
    37250 => -26,
    37251 => -26,
    37252 => -26,
    37253 => -26,
    37254 => -26,
    37255 => -26,
    37256 => -26,
    37257 => -26,
    37258 => -26,
    37259 => -26,
    37260 => -26,
    37261 => -26,
    37262 => -26,
    37263 => -26,
    37264 => -26,
    37265 => -26,
    37266 => -26,
    37267 => -26,
    37268 => -26,
    37269 => -26,
    37270 => -26,
    37271 => -26,
    37272 => -26,
    37273 => -26,
    37274 => -26,
    37275 => -26,
    37276 => -26,
    37277 => -26,
    37278 => -26,
    37279 => -26,
    37280 => -26,
    37281 => -26,
    37282 => -26,
    37283 => -26,
    37284 => -26,
    37285 => -26,
    37286 => -26,
    37287 => -26,
    37288 => -26,
    37289 => -26,
    37290 => -26,
    37291 => -26,
    37292 => -26,
    37293 => -26,
    37294 => -26,
    37295 => -26,
    37296 => -26,
    37297 => -27,
    37298 => -27,
    37299 => -27,
    37300 => -27,
    37301 => -27,
    37302 => -27,
    37303 => -27,
    37304 => -27,
    37305 => -27,
    37306 => -27,
    37307 => -27,
    37308 => -27,
    37309 => -27,
    37310 => -27,
    37311 => -27,
    37312 => -27,
    37313 => -27,
    37314 => -27,
    37315 => -27,
    37316 => -27,
    37317 => -27,
    37318 => -27,
    37319 => -27,
    37320 => -27,
    37321 => -27,
    37322 => -27,
    37323 => -27,
    37324 => -27,
    37325 => -27,
    37326 => -27,
    37327 => -27,
    37328 => -27,
    37329 => -27,
    37330 => -27,
    37331 => -27,
    37332 => -27,
    37333 => -27,
    37334 => -27,
    37335 => -27,
    37336 => -27,
    37337 => -27,
    37338 => -27,
    37339 => -27,
    37340 => -27,
    37341 => -27,
    37342 => -27,
    37343 => -27,
    37344 => -27,
    37345 => -27,
    37346 => -27,
    37347 => -27,
    37348 => -27,
    37349 => -27,
    37350 => -27,
    37351 => -27,
    37352 => -27,
    37353 => -27,
    37354 => -27,
    37355 => -27,
    37356 => -27,
    37357 => -27,
    37358 => -27,
    37359 => -27,
    37360 => -27,
    37361 => -27,
    37362 => -27,
    37363 => -27,
    37364 => -27,
    37365 => -27,
    37366 => -27,
    37367 => -27,
    37368 => -27,
    37369 => -27,
    37370 => -27,
    37371 => -27,
    37372 => -27,
    37373 => -27,
    37374 => -27,
    37375 => -27,
    37376 => -27,
    37377 => -27,
    37378 => -27,
    37379 => -27,
    37380 => -27,
    37381 => -27,
    37382 => -27,
    37383 => -27,
    37384 => -27,
    37385 => -27,
    37386 => -27,
    37387 => -27,
    37388 => -27,
    37389 => -27,
    37390 => -27,
    37391 => -27,
    37392 => -27,
    37393 => -27,
    37394 => -27,
    37395 => -27,
    37396 => -27,
    37397 => -27,
    37398 => -27,
    37399 => -27,
    37400 => -27,
    37401 => -27,
    37402 => -27,
    37403 => -27,
    37404 => -27,
    37405 => -27,
    37406 => -27,
    37407 => -27,
    37408 => -27,
    37409 => -27,
    37410 => -27,
    37411 => -27,
    37412 => -27,
    37413 => -27,
    37414 => -27,
    37415 => -27,
    37416 => -27,
    37417 => -27,
    37418 => -27,
    37419 => -27,
    37420 => -27,
    37421 => -27,
    37422 => -27,
    37423 => -27,
    37424 => -27,
    37425 => -27,
    37426 => -27,
    37427 => -27,
    37428 => -27,
    37429 => -27,
    37430 => -27,
    37431 => -27,
    37432 => -27,
    37433 => -27,
    37434 => -27,
    37435 => -27,
    37436 => -27,
    37437 => -27,
    37438 => -27,
    37439 => -27,
    37440 => -27,
    37441 => -27,
    37442 => -27,
    37443 => -27,
    37444 => -27,
    37445 => -27,
    37446 => -27,
    37447 => -27,
    37448 => -27,
    37449 => -27,
    37450 => -27,
    37451 => -27,
    37452 => -27,
    37453 => -27,
    37454 => -27,
    37455 => -27,
    37456 => -27,
    37457 => -27,
    37458 => -27,
    37459 => -27,
    37460 => -27,
    37461 => -27,
    37462 => -27,
    37463 => -27,
    37464 => -27,
    37465 => -27,
    37466 => -27,
    37467 => -27,
    37468 => -27,
    37469 => -27,
    37470 => -27,
    37471 => -27,
    37472 => -27,
    37473 => -27,
    37474 => -27,
    37475 => -27,
    37476 => -27,
    37477 => -27,
    37478 => -27,
    37479 => -27,
    37480 => -28,
    37481 => -28,
    37482 => -28,
    37483 => -28,
    37484 => -28,
    37485 => -28,
    37486 => -28,
    37487 => -28,
    37488 => -28,
    37489 => -28,
    37490 => -28,
    37491 => -28,
    37492 => -28,
    37493 => -28,
    37494 => -28,
    37495 => -28,
    37496 => -28,
    37497 => -28,
    37498 => -28,
    37499 => -28,
    37500 => -28,
    37501 => -28,
    37502 => -28,
    37503 => -28,
    37504 => -28,
    37505 => -28,
    37506 => -28,
    37507 => -28,
    37508 => -28,
    37509 => -28,
    37510 => -28,
    37511 => -28,
    37512 => -28,
    37513 => -28,
    37514 => -28,
    37515 => -28,
    37516 => -28,
    37517 => -28,
    37518 => -28,
    37519 => -28,
    37520 => -28,
    37521 => -28,
    37522 => -28,
    37523 => -28,
    37524 => -28,
    37525 => -28,
    37526 => -28,
    37527 => -28,
    37528 => -28,
    37529 => -28,
    37530 => -28,
    37531 => -28,
    37532 => -28,
    37533 => -28,
    37534 => -28,
    37535 => -28,
    37536 => -28,
    37537 => -28,
    37538 => -28,
    37539 => -28,
    37540 => -28,
    37541 => -28,
    37542 => -28,
    37543 => -28,
    37544 => -28,
    37545 => -28,
    37546 => -28,
    37547 => -28,
    37548 => -28,
    37549 => -28,
    37550 => -28,
    37551 => -28,
    37552 => -28,
    37553 => -28,
    37554 => -28,
    37555 => -28,
    37556 => -28,
    37557 => -28,
    37558 => -28,
    37559 => -28,
    37560 => -28,
    37561 => -28,
    37562 => -28,
    37563 => -28,
    37564 => -28,
    37565 => -28,
    37566 => -28,
    37567 => -28,
    37568 => -28,
    37569 => -28,
    37570 => -28,
    37571 => -28,
    37572 => -28,
    37573 => -28,
    37574 => -28,
    37575 => -28,
    37576 => -28,
    37577 => -28,
    37578 => -28,
    37579 => -28,
    37580 => -28,
    37581 => -28,
    37582 => -28,
    37583 => -28,
    37584 => -28,
    37585 => -28,
    37586 => -28,
    37587 => -28,
    37588 => -28,
    37589 => -28,
    37590 => -28,
    37591 => -28,
    37592 => -28,
    37593 => -28,
    37594 => -28,
    37595 => -28,
    37596 => -28,
    37597 => -28,
    37598 => -28,
    37599 => -28,
    37600 => -28,
    37601 => -28,
    37602 => -28,
    37603 => -28,
    37604 => -28,
    37605 => -28,
    37606 => -28,
    37607 => -28,
    37608 => -28,
    37609 => -28,
    37610 => -28,
    37611 => -28,
    37612 => -28,
    37613 => -28,
    37614 => -28,
    37615 => -28,
    37616 => -28,
    37617 => -28,
    37618 => -28,
    37619 => -28,
    37620 => -28,
    37621 => -28,
    37622 => -28,
    37623 => -28,
    37624 => -28,
    37625 => -28,
    37626 => -28,
    37627 => -28,
    37628 => -28,
    37629 => -28,
    37630 => -28,
    37631 => -28,
    37632 => -28,
    37633 => -28,
    37634 => -28,
    37635 => -28,
    37636 => -28,
    37637 => -28,
    37638 => -28,
    37639 => -28,
    37640 => -28,
    37641 => -28,
    37642 => -28,
    37643 => -28,
    37644 => -28,
    37645 => -28,
    37646 => -28,
    37647 => -28,
    37648 => -28,
    37649 => -28,
    37650 => -28,
    37651 => -28,
    37652 => -28,
    37653 => -28,
    37654 => -28,
    37655 => -28,
    37656 => -28,
    37657 => -28,
    37658 => -28,
    37659 => -28,
    37660 => -28,
    37661 => -28,
    37662 => -28,
    37663 => -28,
    37664 => -28,
    37665 => -29,
    37666 => -29,
    37667 => -29,
    37668 => -29,
    37669 => -29,
    37670 => -29,
    37671 => -29,
    37672 => -29,
    37673 => -29,
    37674 => -29,
    37675 => -29,
    37676 => -29,
    37677 => -29,
    37678 => -29,
    37679 => -29,
    37680 => -29,
    37681 => -29,
    37682 => -29,
    37683 => -29,
    37684 => -29,
    37685 => -29,
    37686 => -29,
    37687 => -29,
    37688 => -29,
    37689 => -29,
    37690 => -29,
    37691 => -29,
    37692 => -29,
    37693 => -29,
    37694 => -29,
    37695 => -29,
    37696 => -29,
    37697 => -29,
    37698 => -29,
    37699 => -29,
    37700 => -29,
    37701 => -29,
    37702 => -29,
    37703 => -29,
    37704 => -29,
    37705 => -29,
    37706 => -29,
    37707 => -29,
    37708 => -29,
    37709 => -29,
    37710 => -29,
    37711 => -29,
    37712 => -29,
    37713 => -29,
    37714 => -29,
    37715 => -29,
    37716 => -29,
    37717 => -29,
    37718 => -29,
    37719 => -29,
    37720 => -29,
    37721 => -29,
    37722 => -29,
    37723 => -29,
    37724 => -29,
    37725 => -29,
    37726 => -29,
    37727 => -29,
    37728 => -29,
    37729 => -29,
    37730 => -29,
    37731 => -29,
    37732 => -29,
    37733 => -29,
    37734 => -29,
    37735 => -29,
    37736 => -29,
    37737 => -29,
    37738 => -29,
    37739 => -29,
    37740 => -29,
    37741 => -29,
    37742 => -29,
    37743 => -29,
    37744 => -29,
    37745 => -29,
    37746 => -29,
    37747 => -29,
    37748 => -29,
    37749 => -29,
    37750 => -29,
    37751 => -29,
    37752 => -29,
    37753 => -29,
    37754 => -29,
    37755 => -29,
    37756 => -29,
    37757 => -29,
    37758 => -29,
    37759 => -29,
    37760 => -29,
    37761 => -29,
    37762 => -29,
    37763 => -29,
    37764 => -29,
    37765 => -29,
    37766 => -29,
    37767 => -29,
    37768 => -29,
    37769 => -29,
    37770 => -29,
    37771 => -29,
    37772 => -29,
    37773 => -29,
    37774 => -29,
    37775 => -29,
    37776 => -29,
    37777 => -29,
    37778 => -29,
    37779 => -29,
    37780 => -29,
    37781 => -29,
    37782 => -29,
    37783 => -29,
    37784 => -29,
    37785 => -29,
    37786 => -29,
    37787 => -29,
    37788 => -29,
    37789 => -29,
    37790 => -29,
    37791 => -29,
    37792 => -29,
    37793 => -29,
    37794 => -29,
    37795 => -29,
    37796 => -29,
    37797 => -29,
    37798 => -29,
    37799 => -29,
    37800 => -29,
    37801 => -29,
    37802 => -29,
    37803 => -29,
    37804 => -29,
    37805 => -29,
    37806 => -29,
    37807 => -29,
    37808 => -29,
    37809 => -29,
    37810 => -29,
    37811 => -29,
    37812 => -29,
    37813 => -29,
    37814 => -29,
    37815 => -29,
    37816 => -29,
    37817 => -29,
    37818 => -29,
    37819 => -29,
    37820 => -29,
    37821 => -29,
    37822 => -29,
    37823 => -29,
    37824 => -29,
    37825 => -29,
    37826 => -29,
    37827 => -29,
    37828 => -29,
    37829 => -29,
    37830 => -29,
    37831 => -29,
    37832 => -29,
    37833 => -29,
    37834 => -29,
    37835 => -29,
    37836 => -29,
    37837 => -29,
    37838 => -29,
    37839 => -29,
    37840 => -29,
    37841 => -29,
    37842 => -29,
    37843 => -29,
    37844 => -29,
    37845 => -29,
    37846 => -29,
    37847 => -29,
    37848 => -29,
    37849 => -29,
    37850 => -29,
    37851 => -30,
    37852 => -30,
    37853 => -30,
    37854 => -30,
    37855 => -30,
    37856 => -30,
    37857 => -30,
    37858 => -30,
    37859 => -30,
    37860 => -30,
    37861 => -30,
    37862 => -30,
    37863 => -30,
    37864 => -30,
    37865 => -30,
    37866 => -30,
    37867 => -30,
    37868 => -30,
    37869 => -30,
    37870 => -30,
    37871 => -30,
    37872 => -30,
    37873 => -30,
    37874 => -30,
    37875 => -30,
    37876 => -30,
    37877 => -30,
    37878 => -30,
    37879 => -30,
    37880 => -30,
    37881 => -30,
    37882 => -30,
    37883 => -30,
    37884 => -30,
    37885 => -30,
    37886 => -30,
    37887 => -30,
    37888 => -30,
    37889 => -30,
    37890 => -30,
    37891 => -30,
    37892 => -30,
    37893 => -30,
    37894 => -30,
    37895 => -30,
    37896 => -30,
    37897 => -30,
    37898 => -30,
    37899 => -30,
    37900 => -30,
    37901 => -30,
    37902 => -30,
    37903 => -30,
    37904 => -30,
    37905 => -30,
    37906 => -30,
    37907 => -30,
    37908 => -30,
    37909 => -30,
    37910 => -30,
    37911 => -30,
    37912 => -30,
    37913 => -30,
    37914 => -30,
    37915 => -30,
    37916 => -30,
    37917 => -30,
    37918 => -30,
    37919 => -30,
    37920 => -30,
    37921 => -30,
    37922 => -30,
    37923 => -30,
    37924 => -30,
    37925 => -30,
    37926 => -30,
    37927 => -30,
    37928 => -30,
    37929 => -30,
    37930 => -30,
    37931 => -30,
    37932 => -30,
    37933 => -30,
    37934 => -30,
    37935 => -30,
    37936 => -30,
    37937 => -30,
    37938 => -30,
    37939 => -30,
    37940 => -30,
    37941 => -30,
    37942 => -30,
    37943 => -30,
    37944 => -30,
    37945 => -30,
    37946 => -30,
    37947 => -30,
    37948 => -30,
    37949 => -30,
    37950 => -30,
    37951 => -30,
    37952 => -30,
    37953 => -30,
    37954 => -30,
    37955 => -30,
    37956 => -30,
    37957 => -30,
    37958 => -30,
    37959 => -30,
    37960 => -30,
    37961 => -30,
    37962 => -30,
    37963 => -30,
    37964 => -30,
    37965 => -30,
    37966 => -30,
    37967 => -30,
    37968 => -30,
    37969 => -30,
    37970 => -30,
    37971 => -30,
    37972 => -30,
    37973 => -30,
    37974 => -30,
    37975 => -30,
    37976 => -30,
    37977 => -30,
    37978 => -30,
    37979 => -30,
    37980 => -30,
    37981 => -30,
    37982 => -30,
    37983 => -30,
    37984 => -30,
    37985 => -30,
    37986 => -30,
    37987 => -30,
    37988 => -30,
    37989 => -30,
    37990 => -30,
    37991 => -30,
    37992 => -30,
    37993 => -30,
    37994 => -30,
    37995 => -30,
    37996 => -30,
    37997 => -30,
    37998 => -30,
    37999 => -30,
    38000 => -30,
    38001 => -30,
    38002 => -30,
    38003 => -30,
    38004 => -30,
    38005 => -30,
    38006 => -30,
    38007 => -30,
    38008 => -30,
    38009 => -30,
    38010 => -30,
    38011 => -30,
    38012 => -30,
    38013 => -30,
    38014 => -30,
    38015 => -30,
    38016 => -30,
    38017 => -30,
    38018 => -30,
    38019 => -30,
    38020 => -30,
    38021 => -30,
    38022 => -30,
    38023 => -30,
    38024 => -30,
    38025 => -30,
    38026 => -30,
    38027 => -30,
    38028 => -30,
    38029 => -30,
    38030 => -30,
    38031 => -30,
    38032 => -30,
    38033 => -30,
    38034 => -30,
    38035 => -30,
    38036 => -30,
    38037 => -30,
    38038 => -30,
    38039 => -30,
    38040 => -31,
    38041 => -31,
    38042 => -31,
    38043 => -31,
    38044 => -31,
    38045 => -31,
    38046 => -31,
    38047 => -31,
    38048 => -31,
    38049 => -31,
    38050 => -31,
    38051 => -31,
    38052 => -31,
    38053 => -31,
    38054 => -31,
    38055 => -31,
    38056 => -31,
    38057 => -31,
    38058 => -31,
    38059 => -31,
    38060 => -31,
    38061 => -31,
    38062 => -31,
    38063 => -31,
    38064 => -31,
    38065 => -31,
    38066 => -31,
    38067 => -31,
    38068 => -31,
    38069 => -31,
    38070 => -31,
    38071 => -31,
    38072 => -31,
    38073 => -31,
    38074 => -31,
    38075 => -31,
    38076 => -31,
    38077 => -31,
    38078 => -31,
    38079 => -31,
    38080 => -31,
    38081 => -31,
    38082 => -31,
    38083 => -31,
    38084 => -31,
    38085 => -31,
    38086 => -31,
    38087 => -31,
    38088 => -31,
    38089 => -31,
    38090 => -31,
    38091 => -31,
    38092 => -31,
    38093 => -31,
    38094 => -31,
    38095 => -31,
    38096 => -31,
    38097 => -31,
    38098 => -31,
    38099 => -31,
    38100 => -31,
    38101 => -31,
    38102 => -31,
    38103 => -31,
    38104 => -31,
    38105 => -31,
    38106 => -31,
    38107 => -31,
    38108 => -31,
    38109 => -31,
    38110 => -31,
    38111 => -31,
    38112 => -31,
    38113 => -31,
    38114 => -31,
    38115 => -31,
    38116 => -31,
    38117 => -31,
    38118 => -31,
    38119 => -31,
    38120 => -31,
    38121 => -31,
    38122 => -31,
    38123 => -31,
    38124 => -31,
    38125 => -31,
    38126 => -31,
    38127 => -31,
    38128 => -31,
    38129 => -31,
    38130 => -31,
    38131 => -31,
    38132 => -31,
    38133 => -31,
    38134 => -31,
    38135 => -31,
    38136 => -31,
    38137 => -31,
    38138 => -31,
    38139 => -31,
    38140 => -31,
    38141 => -31,
    38142 => -31,
    38143 => -31,
    38144 => -31,
    38145 => -31,
    38146 => -31,
    38147 => -31,
    38148 => -31,
    38149 => -31,
    38150 => -31,
    38151 => -31,
    38152 => -31,
    38153 => -31,
    38154 => -31,
    38155 => -31,
    38156 => -31,
    38157 => -31,
    38158 => -31,
    38159 => -31,
    38160 => -31,
    38161 => -31,
    38162 => -31,
    38163 => -31,
    38164 => -31,
    38165 => -31,
    38166 => -31,
    38167 => -31,
    38168 => -31,
    38169 => -31,
    38170 => -31,
    38171 => -31,
    38172 => -31,
    38173 => -31,
    38174 => -31,
    38175 => -31,
    38176 => -31,
    38177 => -31,
    38178 => -31,
    38179 => -31,
    38180 => -31,
    38181 => -31,
    38182 => -31,
    38183 => -31,
    38184 => -31,
    38185 => -31,
    38186 => -31,
    38187 => -31,
    38188 => -31,
    38189 => -31,
    38190 => -31,
    38191 => -31,
    38192 => -31,
    38193 => -31,
    38194 => -31,
    38195 => -31,
    38196 => -31,
    38197 => -31,
    38198 => -31,
    38199 => -31,
    38200 => -31,
    38201 => -31,
    38202 => -31,
    38203 => -31,
    38204 => -31,
    38205 => -31,
    38206 => -31,
    38207 => -31,
    38208 => -31,
    38209 => -31,
    38210 => -31,
    38211 => -31,
    38212 => -31,
    38213 => -31,
    38214 => -31,
    38215 => -31,
    38216 => -31,
    38217 => -31,
    38218 => -31,
    38219 => -31,
    38220 => -31,
    38221 => -31,
    38222 => -31,
    38223 => -31,
    38224 => -31,
    38225 => -31,
    38226 => -31,
    38227 => -31,
    38228 => -31,
    38229 => -31,
    38230 => -32,
    38231 => -32,
    38232 => -32,
    38233 => -32,
    38234 => -32,
    38235 => -32,
    38236 => -32,
    38237 => -32,
    38238 => -32,
    38239 => -32,
    38240 => -32,
    38241 => -32,
    38242 => -32,
    38243 => -32,
    38244 => -32,
    38245 => -32,
    38246 => -32,
    38247 => -32,
    38248 => -32,
    38249 => -32,
    38250 => -32,
    38251 => -32,
    38252 => -32,
    38253 => -32,
    38254 => -32,
    38255 => -32,
    38256 => -32,
    38257 => -32,
    38258 => -32,
    38259 => -32,
    38260 => -32,
    38261 => -32,
    38262 => -32,
    38263 => -32,
    38264 => -32,
    38265 => -32,
    38266 => -32,
    38267 => -32,
    38268 => -32,
    38269 => -32,
    38270 => -32,
    38271 => -32,
    38272 => -32,
    38273 => -32,
    38274 => -32,
    38275 => -32,
    38276 => -32,
    38277 => -32,
    38278 => -32,
    38279 => -32,
    38280 => -32,
    38281 => -32,
    38282 => -32,
    38283 => -32,
    38284 => -32,
    38285 => -32,
    38286 => -32,
    38287 => -32,
    38288 => -32,
    38289 => -32,
    38290 => -32,
    38291 => -32,
    38292 => -32,
    38293 => -32,
    38294 => -32,
    38295 => -32,
    38296 => -32,
    38297 => -32,
    38298 => -32,
    38299 => -32,
    38300 => -32,
    38301 => -32,
    38302 => -32,
    38303 => -32,
    38304 => -32,
    38305 => -32,
    38306 => -32,
    38307 => -32,
    38308 => -32,
    38309 => -32,
    38310 => -32,
    38311 => -32,
    38312 => -32,
    38313 => -32,
    38314 => -32,
    38315 => -32,
    38316 => -32,
    38317 => -32,
    38318 => -32,
    38319 => -32,
    38320 => -32,
    38321 => -32,
    38322 => -32,
    38323 => -32,
    38324 => -32,
    38325 => -32,
    38326 => -32,
    38327 => -32,
    38328 => -32,
    38329 => -32,
    38330 => -32,
    38331 => -32,
    38332 => -32,
    38333 => -32,
    38334 => -32,
    38335 => -32,
    38336 => -32,
    38337 => -32,
    38338 => -32,
    38339 => -32,
    38340 => -32,
    38341 => -32,
    38342 => -32,
    38343 => -32,
    38344 => -32,
    38345 => -32,
    38346 => -32,
    38347 => -32,
    38348 => -32,
    38349 => -32,
    38350 => -32,
    38351 => -32,
    38352 => -32,
    38353 => -32,
    38354 => -32,
    38355 => -32,
    38356 => -32,
    38357 => -32,
    38358 => -32,
    38359 => -32,
    38360 => -32,
    38361 => -32,
    38362 => -32,
    38363 => -32,
    38364 => -32,
    38365 => -32,
    38366 => -32,
    38367 => -32,
    38368 => -32,
    38369 => -32,
    38370 => -32,
    38371 => -32,
    38372 => -32,
    38373 => -32,
    38374 => -32,
    38375 => -32,
    38376 => -32,
    38377 => -32,
    38378 => -32,
    38379 => -32,
    38380 => -32,
    38381 => -32,
    38382 => -32,
    38383 => -32,
    38384 => -32,
    38385 => -32,
    38386 => -32,
    38387 => -32,
    38388 => -32,
    38389 => -32,
    38390 => -32,
    38391 => -32,
    38392 => -32,
    38393 => -32,
    38394 => -32,
    38395 => -32,
    38396 => -32,
    38397 => -32,
    38398 => -32,
    38399 => -32,
    38400 => -32,
    38401 => -32,
    38402 => -32,
    38403 => -32,
    38404 => -32,
    38405 => -32,
    38406 => -32,
    38407 => -32,
    38408 => -32,
    38409 => -32,
    38410 => -32,
    38411 => -32,
    38412 => -32,
    38413 => -32,
    38414 => -32,
    38415 => -32,
    38416 => -32,
    38417 => -32,
    38418 => -32,
    38419 => -32,
    38420 => -32,
    38421 => -32,
    38422 => -33,
    38423 => -33,
    38424 => -33,
    38425 => -33,
    38426 => -33,
    38427 => -33,
    38428 => -33,
    38429 => -33,
    38430 => -33,
    38431 => -33,
    38432 => -33,
    38433 => -33,
    38434 => -33,
    38435 => -33,
    38436 => -33,
    38437 => -33,
    38438 => -33,
    38439 => -33,
    38440 => -33,
    38441 => -33,
    38442 => -33,
    38443 => -33,
    38444 => -33,
    38445 => -33,
    38446 => -33,
    38447 => -33,
    38448 => -33,
    38449 => -33,
    38450 => -33,
    38451 => -33,
    38452 => -33,
    38453 => -33,
    38454 => -33,
    38455 => -33,
    38456 => -33,
    38457 => -33,
    38458 => -33,
    38459 => -33,
    38460 => -33,
    38461 => -33,
    38462 => -33,
    38463 => -33,
    38464 => -33,
    38465 => -33,
    38466 => -33,
    38467 => -33,
    38468 => -33,
    38469 => -33,
    38470 => -33,
    38471 => -33,
    38472 => -33,
    38473 => -33,
    38474 => -33,
    38475 => -33,
    38476 => -33,
    38477 => -33,
    38478 => -33,
    38479 => -33,
    38480 => -33,
    38481 => -33,
    38482 => -33,
    38483 => -33,
    38484 => -33,
    38485 => -33,
    38486 => -33,
    38487 => -33,
    38488 => -33,
    38489 => -33,
    38490 => -33,
    38491 => -33,
    38492 => -33,
    38493 => -33,
    38494 => -33,
    38495 => -33,
    38496 => -33,
    38497 => -33,
    38498 => -33,
    38499 => -33,
    38500 => -33,
    38501 => -33,
    38502 => -33,
    38503 => -33,
    38504 => -33,
    38505 => -33,
    38506 => -33,
    38507 => -33,
    38508 => -33,
    38509 => -33,
    38510 => -33,
    38511 => -33,
    38512 => -33,
    38513 => -33,
    38514 => -33,
    38515 => -33,
    38516 => -33,
    38517 => -33,
    38518 => -33,
    38519 => -33,
    38520 => -33,
    38521 => -33,
    38522 => -33,
    38523 => -33,
    38524 => -33,
    38525 => -33,
    38526 => -33,
    38527 => -33,
    38528 => -33,
    38529 => -33,
    38530 => -33,
    38531 => -33,
    38532 => -33,
    38533 => -33,
    38534 => -33,
    38535 => -33,
    38536 => -33,
    38537 => -33,
    38538 => -33,
    38539 => -33,
    38540 => -33,
    38541 => -33,
    38542 => -33,
    38543 => -33,
    38544 => -33,
    38545 => -33,
    38546 => -33,
    38547 => -33,
    38548 => -33,
    38549 => -33,
    38550 => -33,
    38551 => -33,
    38552 => -33,
    38553 => -33,
    38554 => -33,
    38555 => -33,
    38556 => -33,
    38557 => -33,
    38558 => -33,
    38559 => -33,
    38560 => -33,
    38561 => -33,
    38562 => -33,
    38563 => -33,
    38564 => -33,
    38565 => -33,
    38566 => -33,
    38567 => -33,
    38568 => -33,
    38569 => -33,
    38570 => -33,
    38571 => -33,
    38572 => -33,
    38573 => -33,
    38574 => -33,
    38575 => -33,
    38576 => -33,
    38577 => -33,
    38578 => -33,
    38579 => -33,
    38580 => -33,
    38581 => -33,
    38582 => -33,
    38583 => -33,
    38584 => -33,
    38585 => -33,
    38586 => -33,
    38587 => -33,
    38588 => -33,
    38589 => -33,
    38590 => -33,
    38591 => -33,
    38592 => -33,
    38593 => -33,
    38594 => -33,
    38595 => -33,
    38596 => -33,
    38597 => -33,
    38598 => -33,
    38599 => -33,
    38600 => -33,
    38601 => -33,
    38602 => -33,
    38603 => -33,
    38604 => -33,
    38605 => -33,
    38606 => -33,
    38607 => -33,
    38608 => -33,
    38609 => -33,
    38610 => -33,
    38611 => -33,
    38612 => -33,
    38613 => -33,
    38614 => -33,
    38615 => -33,
    38616 => -34,
    38617 => -34,
    38618 => -34,
    38619 => -34,
    38620 => -34,
    38621 => -34,
    38622 => -34,
    38623 => -34,
    38624 => -34,
    38625 => -34,
    38626 => -34,
    38627 => -34,
    38628 => -34,
    38629 => -34,
    38630 => -34,
    38631 => -34,
    38632 => -34,
    38633 => -34,
    38634 => -34,
    38635 => -34,
    38636 => -34,
    38637 => -34,
    38638 => -34,
    38639 => -34,
    38640 => -34,
    38641 => -34,
    38642 => -34,
    38643 => -34,
    38644 => -34,
    38645 => -34,
    38646 => -34,
    38647 => -34,
    38648 => -34,
    38649 => -34,
    38650 => -34,
    38651 => -34,
    38652 => -34,
    38653 => -34,
    38654 => -34,
    38655 => -34,
    38656 => -34,
    38657 => -34,
    38658 => -34,
    38659 => -34,
    38660 => -34,
    38661 => -34,
    38662 => -34,
    38663 => -34,
    38664 => -34,
    38665 => -34,
    38666 => -34,
    38667 => -34,
    38668 => -34,
    38669 => -34,
    38670 => -34,
    38671 => -34,
    38672 => -34,
    38673 => -34,
    38674 => -34,
    38675 => -34,
    38676 => -34,
    38677 => -34,
    38678 => -34,
    38679 => -34,
    38680 => -34,
    38681 => -34,
    38682 => -34,
    38683 => -34,
    38684 => -34,
    38685 => -34,
    38686 => -34,
    38687 => -34,
    38688 => -34,
    38689 => -34,
    38690 => -34,
    38691 => -34,
    38692 => -34,
    38693 => -34,
    38694 => -34,
    38695 => -34,
    38696 => -34,
    38697 => -34,
    38698 => -34,
    38699 => -34,
    38700 => -34,
    38701 => -34,
    38702 => -34,
    38703 => -34,
    38704 => -34,
    38705 => -34,
    38706 => -34,
    38707 => -34,
    38708 => -34,
    38709 => -34,
    38710 => -34,
    38711 => -34,
    38712 => -34,
    38713 => -34,
    38714 => -34,
    38715 => -34,
    38716 => -34,
    38717 => -34,
    38718 => -34,
    38719 => -34,
    38720 => -34,
    38721 => -34,
    38722 => -34,
    38723 => -34,
    38724 => -34,
    38725 => -34,
    38726 => -34,
    38727 => -34,
    38728 => -34,
    38729 => -34,
    38730 => -34,
    38731 => -34,
    38732 => -34,
    38733 => -34,
    38734 => -34,
    38735 => -34,
    38736 => -34,
    38737 => -34,
    38738 => -34,
    38739 => -34,
    38740 => -34,
    38741 => -34,
    38742 => -34,
    38743 => -34,
    38744 => -34,
    38745 => -34,
    38746 => -34,
    38747 => -34,
    38748 => -34,
    38749 => -34,
    38750 => -34,
    38751 => -34,
    38752 => -34,
    38753 => -34,
    38754 => -34,
    38755 => -34,
    38756 => -34,
    38757 => -34,
    38758 => -34,
    38759 => -34,
    38760 => -34,
    38761 => -34,
    38762 => -34,
    38763 => -34,
    38764 => -34,
    38765 => -34,
    38766 => -34,
    38767 => -34,
    38768 => -34,
    38769 => -34,
    38770 => -34,
    38771 => -34,
    38772 => -34,
    38773 => -34,
    38774 => -34,
    38775 => -34,
    38776 => -34,
    38777 => -34,
    38778 => -34,
    38779 => -34,
    38780 => -34,
    38781 => -34,
    38782 => -34,
    38783 => -34,
    38784 => -34,
    38785 => -34,
    38786 => -34,
    38787 => -34,
    38788 => -34,
    38789 => -34,
    38790 => -34,
    38791 => -34,
    38792 => -34,
    38793 => -34,
    38794 => -34,
    38795 => -34,
    38796 => -34,
    38797 => -34,
    38798 => -34,
    38799 => -34,
    38800 => -34,
    38801 => -34,
    38802 => -34,
    38803 => -34,
    38804 => -34,
    38805 => -34,
    38806 => -34,
    38807 => -34,
    38808 => -34,
    38809 => -34,
    38810 => -34,
    38811 => -34,
    38812 => -34,
    38813 => -35,
    38814 => -35,
    38815 => -35,
    38816 => -35,
    38817 => -35,
    38818 => -35,
    38819 => -35,
    38820 => -35,
    38821 => -35,
    38822 => -35,
    38823 => -35,
    38824 => -35,
    38825 => -35,
    38826 => -35,
    38827 => -35,
    38828 => -35,
    38829 => -35,
    38830 => -35,
    38831 => -35,
    38832 => -35,
    38833 => -35,
    38834 => -35,
    38835 => -35,
    38836 => -35,
    38837 => -35,
    38838 => -35,
    38839 => -35,
    38840 => -35,
    38841 => -35,
    38842 => -35,
    38843 => -35,
    38844 => -35,
    38845 => -35,
    38846 => -35,
    38847 => -35,
    38848 => -35,
    38849 => -35,
    38850 => -35,
    38851 => -35,
    38852 => -35,
    38853 => -35,
    38854 => -35,
    38855 => -35,
    38856 => -35,
    38857 => -35,
    38858 => -35,
    38859 => -35,
    38860 => -35,
    38861 => -35,
    38862 => -35,
    38863 => -35,
    38864 => -35,
    38865 => -35,
    38866 => -35,
    38867 => -35,
    38868 => -35,
    38869 => -35,
    38870 => -35,
    38871 => -35,
    38872 => -35,
    38873 => -35,
    38874 => -35,
    38875 => -35,
    38876 => -35,
    38877 => -35,
    38878 => -35,
    38879 => -35,
    38880 => -35,
    38881 => -35,
    38882 => -35,
    38883 => -35,
    38884 => -35,
    38885 => -35,
    38886 => -35,
    38887 => -35,
    38888 => -35,
    38889 => -35,
    38890 => -35,
    38891 => -35,
    38892 => -35,
    38893 => -35,
    38894 => -35,
    38895 => -35,
    38896 => -35,
    38897 => -35,
    38898 => -35,
    38899 => -35,
    38900 => -35,
    38901 => -35,
    38902 => -35,
    38903 => -35,
    38904 => -35,
    38905 => -35,
    38906 => -35,
    38907 => -35,
    38908 => -35,
    38909 => -35,
    38910 => -35,
    38911 => -35,
    38912 => -35,
    38913 => -35,
    38914 => -35,
    38915 => -35,
    38916 => -35,
    38917 => -35,
    38918 => -35,
    38919 => -35,
    38920 => -35,
    38921 => -35,
    38922 => -35,
    38923 => -35,
    38924 => -35,
    38925 => -35,
    38926 => -35,
    38927 => -35,
    38928 => -35,
    38929 => -35,
    38930 => -35,
    38931 => -35,
    38932 => -35,
    38933 => -35,
    38934 => -35,
    38935 => -35,
    38936 => -35,
    38937 => -35,
    38938 => -35,
    38939 => -35,
    38940 => -35,
    38941 => -35,
    38942 => -35,
    38943 => -35,
    38944 => -35,
    38945 => -35,
    38946 => -35,
    38947 => -35,
    38948 => -35,
    38949 => -35,
    38950 => -35,
    38951 => -35,
    38952 => -35,
    38953 => -35,
    38954 => -35,
    38955 => -35,
    38956 => -35,
    38957 => -35,
    38958 => -35,
    38959 => -35,
    38960 => -35,
    38961 => -35,
    38962 => -35,
    38963 => -35,
    38964 => -35,
    38965 => -35,
    38966 => -35,
    38967 => -35,
    38968 => -35,
    38969 => -35,
    38970 => -35,
    38971 => -35,
    38972 => -35,
    38973 => -35,
    38974 => -35,
    38975 => -35,
    38976 => -35,
    38977 => -35,
    38978 => -35,
    38979 => -35,
    38980 => -35,
    38981 => -35,
    38982 => -35,
    38983 => -35,
    38984 => -35,
    38985 => -35,
    38986 => -35,
    38987 => -35,
    38988 => -35,
    38989 => -35,
    38990 => -35,
    38991 => -35,
    38992 => -35,
    38993 => -35,
    38994 => -35,
    38995 => -35,
    38996 => -35,
    38997 => -35,
    38998 => -35,
    38999 => -35,
    39000 => -35,
    39001 => -35,
    39002 => -35,
    39003 => -35,
    39004 => -35,
    39005 => -35,
    39006 => -35,
    39007 => -35,
    39008 => -35,
    39009 => -35,
    39010 => -35,
    39011 => -35,
    39012 => -36,
    39013 => -36,
    39014 => -36,
    39015 => -36,
    39016 => -36,
    39017 => -36,
    39018 => -36,
    39019 => -36,
    39020 => -36,
    39021 => -36,
    39022 => -36,
    39023 => -36,
    39024 => -36,
    39025 => -36,
    39026 => -36,
    39027 => -36,
    39028 => -36,
    39029 => -36,
    39030 => -36,
    39031 => -36,
    39032 => -36,
    39033 => -36,
    39034 => -36,
    39035 => -36,
    39036 => -36,
    39037 => -36,
    39038 => -36,
    39039 => -36,
    39040 => -36,
    39041 => -36,
    39042 => -36,
    39043 => -36,
    39044 => -36,
    39045 => -36,
    39046 => -36,
    39047 => -36,
    39048 => -36,
    39049 => -36,
    39050 => -36,
    39051 => -36,
    39052 => -36,
    39053 => -36,
    39054 => -36,
    39055 => -36,
    39056 => -36,
    39057 => -36,
    39058 => -36,
    39059 => -36,
    39060 => -36,
    39061 => -36,
    39062 => -36,
    39063 => -36,
    39064 => -36,
    39065 => -36,
    39066 => -36,
    39067 => -36,
    39068 => -36,
    39069 => -36,
    39070 => -36,
    39071 => -36,
    39072 => -36,
    39073 => -36,
    39074 => -36,
    39075 => -36,
    39076 => -36,
    39077 => -36,
    39078 => -36,
    39079 => -36,
    39080 => -36,
    39081 => -36,
    39082 => -36,
    39083 => -36,
    39084 => -36,
    39085 => -36,
    39086 => -36,
    39087 => -36,
    39088 => -36,
    39089 => -36,
    39090 => -36,
    39091 => -36,
    39092 => -36,
    39093 => -36,
    39094 => -36,
    39095 => -36,
    39096 => -36,
    39097 => -36,
    39098 => -36,
    39099 => -36,
    39100 => -36,
    39101 => -36,
    39102 => -36,
    39103 => -36,
    39104 => -36,
    39105 => -36,
    39106 => -36,
    39107 => -36,
    39108 => -36,
    39109 => -36,
    39110 => -36,
    39111 => -36,
    39112 => -36,
    39113 => -36,
    39114 => -36,
    39115 => -36,
    39116 => -36,
    39117 => -36,
    39118 => -36,
    39119 => -36,
    39120 => -36,
    39121 => -36,
    39122 => -36,
    39123 => -36,
    39124 => -36,
    39125 => -36,
    39126 => -36,
    39127 => -36,
    39128 => -36,
    39129 => -36,
    39130 => -36,
    39131 => -36,
    39132 => -36,
    39133 => -36,
    39134 => -36,
    39135 => -36,
    39136 => -36,
    39137 => -36,
    39138 => -36,
    39139 => -36,
    39140 => -36,
    39141 => -36,
    39142 => -36,
    39143 => -36,
    39144 => -36,
    39145 => -36,
    39146 => -36,
    39147 => -36,
    39148 => -36,
    39149 => -36,
    39150 => -36,
    39151 => -36,
    39152 => -36,
    39153 => -36,
    39154 => -36,
    39155 => -36,
    39156 => -36,
    39157 => -36,
    39158 => -36,
    39159 => -36,
    39160 => -36,
    39161 => -36,
    39162 => -36,
    39163 => -36,
    39164 => -36,
    39165 => -36,
    39166 => -36,
    39167 => -36,
    39168 => -36,
    39169 => -36,
    39170 => -36,
    39171 => -36,
    39172 => -36,
    39173 => -36,
    39174 => -36,
    39175 => -36,
    39176 => -36,
    39177 => -36,
    39178 => -36,
    39179 => -36,
    39180 => -36,
    39181 => -36,
    39182 => -36,
    39183 => -36,
    39184 => -36,
    39185 => -36,
    39186 => -36,
    39187 => -36,
    39188 => -36,
    39189 => -36,
    39190 => -36,
    39191 => -36,
    39192 => -36,
    39193 => -36,
    39194 => -36,
    39195 => -36,
    39196 => -36,
    39197 => -36,
    39198 => -36,
    39199 => -36,
    39200 => -36,
    39201 => -36,
    39202 => -36,
    39203 => -36,
    39204 => -36,
    39205 => -36,
    39206 => -36,
    39207 => -36,
    39208 => -36,
    39209 => -36,
    39210 => -36,
    39211 => -36,
    39212 => -36,
    39213 => -36,
    39214 => -37,
    39215 => -37,
    39216 => -37,
    39217 => -37,
    39218 => -37,
    39219 => -37,
    39220 => -37,
    39221 => -37,
    39222 => -37,
    39223 => -37,
    39224 => -37,
    39225 => -37,
    39226 => -37,
    39227 => -37,
    39228 => -37,
    39229 => -37,
    39230 => -37,
    39231 => -37,
    39232 => -37,
    39233 => -37,
    39234 => -37,
    39235 => -37,
    39236 => -37,
    39237 => -37,
    39238 => -37,
    39239 => -37,
    39240 => -37,
    39241 => -37,
    39242 => -37,
    39243 => -37,
    39244 => -37,
    39245 => -37,
    39246 => -37,
    39247 => -37,
    39248 => -37,
    39249 => -37,
    39250 => -37,
    39251 => -37,
    39252 => -37,
    39253 => -37,
    39254 => -37,
    39255 => -37,
    39256 => -37,
    39257 => -37,
    39258 => -37,
    39259 => -37,
    39260 => -37,
    39261 => -37,
    39262 => -37,
    39263 => -37,
    39264 => -37,
    39265 => -37,
    39266 => -37,
    39267 => -37,
    39268 => -37,
    39269 => -37,
    39270 => -37,
    39271 => -37,
    39272 => -37,
    39273 => -37,
    39274 => -37,
    39275 => -37,
    39276 => -37,
    39277 => -37,
    39278 => -37,
    39279 => -37,
    39280 => -37,
    39281 => -37,
    39282 => -37,
    39283 => -37,
    39284 => -37,
    39285 => -37,
    39286 => -37,
    39287 => -37,
    39288 => -37,
    39289 => -37,
    39290 => -37,
    39291 => -37,
    39292 => -37,
    39293 => -37,
    39294 => -37,
    39295 => -37,
    39296 => -37,
    39297 => -37,
    39298 => -37,
    39299 => -37,
    39300 => -37,
    39301 => -37,
    39302 => -37,
    39303 => -37,
    39304 => -37,
    39305 => -37,
    39306 => -37,
    39307 => -37,
    39308 => -37,
    39309 => -37,
    39310 => -37,
    39311 => -37,
    39312 => -37,
    39313 => -37,
    39314 => -37,
    39315 => -37,
    39316 => -37,
    39317 => -37,
    39318 => -37,
    39319 => -37,
    39320 => -37,
    39321 => -37,
    39322 => -37,
    39323 => -37,
    39324 => -37,
    39325 => -37,
    39326 => -37,
    39327 => -37,
    39328 => -37,
    39329 => -37,
    39330 => -37,
    39331 => -37,
    39332 => -37,
    39333 => -37,
    39334 => -37,
    39335 => -37,
    39336 => -37,
    39337 => -37,
    39338 => -37,
    39339 => -37,
    39340 => -37,
    39341 => -37,
    39342 => -37,
    39343 => -37,
    39344 => -37,
    39345 => -37,
    39346 => -37,
    39347 => -37,
    39348 => -37,
    39349 => -37,
    39350 => -37,
    39351 => -37,
    39352 => -37,
    39353 => -37,
    39354 => -37,
    39355 => -37,
    39356 => -37,
    39357 => -37,
    39358 => -37,
    39359 => -37,
    39360 => -37,
    39361 => -37,
    39362 => -37,
    39363 => -37,
    39364 => -37,
    39365 => -37,
    39366 => -37,
    39367 => -37,
    39368 => -37,
    39369 => -37,
    39370 => -37,
    39371 => -37,
    39372 => -37,
    39373 => -37,
    39374 => -37,
    39375 => -37,
    39376 => -37,
    39377 => -37,
    39378 => -37,
    39379 => -37,
    39380 => -37,
    39381 => -37,
    39382 => -37,
    39383 => -37,
    39384 => -37,
    39385 => -37,
    39386 => -37,
    39387 => -37,
    39388 => -37,
    39389 => -37,
    39390 => -37,
    39391 => -37,
    39392 => -37,
    39393 => -37,
    39394 => -37,
    39395 => -37,
    39396 => -37,
    39397 => -37,
    39398 => -37,
    39399 => -37,
    39400 => -37,
    39401 => -37,
    39402 => -37,
    39403 => -37,
    39404 => -37,
    39405 => -37,
    39406 => -37,
    39407 => -37,
    39408 => -37,
    39409 => -37,
    39410 => -37,
    39411 => -37,
    39412 => -37,
    39413 => -37,
    39414 => -37,
    39415 => -37,
    39416 => -37,
    39417 => -37,
    39418 => -37,
    39419 => -38,
    39420 => -38,
    39421 => -38,
    39422 => -38,
    39423 => -38,
    39424 => -38,
    39425 => -38,
    39426 => -38,
    39427 => -38,
    39428 => -38,
    39429 => -38,
    39430 => -38,
    39431 => -38,
    39432 => -38,
    39433 => -38,
    39434 => -38,
    39435 => -38,
    39436 => -38,
    39437 => -38,
    39438 => -38,
    39439 => -38,
    39440 => -38,
    39441 => -38,
    39442 => -38,
    39443 => -38,
    39444 => -38,
    39445 => -38,
    39446 => -38,
    39447 => -38,
    39448 => -38,
    39449 => -38,
    39450 => -38,
    39451 => -38,
    39452 => -38,
    39453 => -38,
    39454 => -38,
    39455 => -38,
    39456 => -38,
    39457 => -38,
    39458 => -38,
    39459 => -38,
    39460 => -38,
    39461 => -38,
    39462 => -38,
    39463 => -38,
    39464 => -38,
    39465 => -38,
    39466 => -38,
    39467 => -38,
    39468 => -38,
    39469 => -38,
    39470 => -38,
    39471 => -38,
    39472 => -38,
    39473 => -38,
    39474 => -38,
    39475 => -38,
    39476 => -38,
    39477 => -38,
    39478 => -38,
    39479 => -38,
    39480 => -38,
    39481 => -38,
    39482 => -38,
    39483 => -38,
    39484 => -38,
    39485 => -38,
    39486 => -38,
    39487 => -38,
    39488 => -38,
    39489 => -38,
    39490 => -38,
    39491 => -38,
    39492 => -38,
    39493 => -38,
    39494 => -38,
    39495 => -38,
    39496 => -38,
    39497 => -38,
    39498 => -38,
    39499 => -38,
    39500 => -38,
    39501 => -38,
    39502 => -38,
    39503 => -38,
    39504 => -38,
    39505 => -38,
    39506 => -38,
    39507 => -38,
    39508 => -38,
    39509 => -38,
    39510 => -38,
    39511 => -38,
    39512 => -38,
    39513 => -38,
    39514 => -38,
    39515 => -38,
    39516 => -38,
    39517 => -38,
    39518 => -38,
    39519 => -38,
    39520 => -38,
    39521 => -38,
    39522 => -38,
    39523 => -38,
    39524 => -38,
    39525 => -38,
    39526 => -38,
    39527 => -38,
    39528 => -38,
    39529 => -38,
    39530 => -38,
    39531 => -38,
    39532 => -38,
    39533 => -38,
    39534 => -38,
    39535 => -38,
    39536 => -38,
    39537 => -38,
    39538 => -38,
    39539 => -38,
    39540 => -38,
    39541 => -38,
    39542 => -38,
    39543 => -38,
    39544 => -38,
    39545 => -38,
    39546 => -38,
    39547 => -38,
    39548 => -38,
    39549 => -38,
    39550 => -38,
    39551 => -38,
    39552 => -38,
    39553 => -38,
    39554 => -38,
    39555 => -38,
    39556 => -38,
    39557 => -38,
    39558 => -38,
    39559 => -38,
    39560 => -38,
    39561 => -38,
    39562 => -38,
    39563 => -38,
    39564 => -38,
    39565 => -38,
    39566 => -38,
    39567 => -38,
    39568 => -38,
    39569 => -38,
    39570 => -38,
    39571 => -38,
    39572 => -38,
    39573 => -38,
    39574 => -38,
    39575 => -38,
    39576 => -38,
    39577 => -38,
    39578 => -38,
    39579 => -38,
    39580 => -38,
    39581 => -38,
    39582 => -38,
    39583 => -38,
    39584 => -38,
    39585 => -38,
    39586 => -38,
    39587 => -38,
    39588 => -38,
    39589 => -38,
    39590 => -38,
    39591 => -38,
    39592 => -38,
    39593 => -38,
    39594 => -38,
    39595 => -38,
    39596 => -38,
    39597 => -38,
    39598 => -38,
    39599 => -38,
    39600 => -38,
    39601 => -38,
    39602 => -38,
    39603 => -38,
    39604 => -38,
    39605 => -38,
    39606 => -38,
    39607 => -38,
    39608 => -38,
    39609 => -38,
    39610 => -38,
    39611 => -38,
    39612 => -38,
    39613 => -38,
    39614 => -38,
    39615 => -38,
    39616 => -38,
    39617 => -38,
    39618 => -38,
    39619 => -38,
    39620 => -38,
    39621 => -38,
    39622 => -38,
    39623 => -38,
    39624 => -38,
    39625 => -38,
    39626 => -39,
    39627 => -39,
    39628 => -39,
    39629 => -39,
    39630 => -39,
    39631 => -39,
    39632 => -39,
    39633 => -39,
    39634 => -39,
    39635 => -39,
    39636 => -39,
    39637 => -39,
    39638 => -39,
    39639 => -39,
    39640 => -39,
    39641 => -39,
    39642 => -39,
    39643 => -39,
    39644 => -39,
    39645 => -39,
    39646 => -39,
    39647 => -39,
    39648 => -39,
    39649 => -39,
    39650 => -39,
    39651 => -39,
    39652 => -39,
    39653 => -39,
    39654 => -39,
    39655 => -39,
    39656 => -39,
    39657 => -39,
    39658 => -39,
    39659 => -39,
    39660 => -39,
    39661 => -39,
    39662 => -39,
    39663 => -39,
    39664 => -39,
    39665 => -39,
    39666 => -39,
    39667 => -39,
    39668 => -39,
    39669 => -39,
    39670 => -39,
    39671 => -39,
    39672 => -39,
    39673 => -39,
    39674 => -39,
    39675 => -39,
    39676 => -39,
    39677 => -39,
    39678 => -39,
    39679 => -39,
    39680 => -39,
    39681 => -39,
    39682 => -39,
    39683 => -39,
    39684 => -39,
    39685 => -39,
    39686 => -39,
    39687 => -39,
    39688 => -39,
    39689 => -39,
    39690 => -39,
    39691 => -39,
    39692 => -39,
    39693 => -39,
    39694 => -39,
    39695 => -39,
    39696 => -39,
    39697 => -39,
    39698 => -39,
    39699 => -39,
    39700 => -39,
    39701 => -39,
    39702 => -39,
    39703 => -39,
    39704 => -39,
    39705 => -39,
    39706 => -39,
    39707 => -39,
    39708 => -39,
    39709 => -39,
    39710 => -39,
    39711 => -39,
    39712 => -39,
    39713 => -39,
    39714 => -39,
    39715 => -39,
    39716 => -39,
    39717 => -39,
    39718 => -39,
    39719 => -39,
    39720 => -39,
    39721 => -39,
    39722 => -39,
    39723 => -39,
    39724 => -39,
    39725 => -39,
    39726 => -39,
    39727 => -39,
    39728 => -39,
    39729 => -39,
    39730 => -39,
    39731 => -39,
    39732 => -39,
    39733 => -39,
    39734 => -39,
    39735 => -39,
    39736 => -39,
    39737 => -39,
    39738 => -39,
    39739 => -39,
    39740 => -39,
    39741 => -39,
    39742 => -39,
    39743 => -39,
    39744 => -39,
    39745 => -39,
    39746 => -39,
    39747 => -39,
    39748 => -39,
    39749 => -39,
    39750 => -39,
    39751 => -39,
    39752 => -39,
    39753 => -39,
    39754 => -39,
    39755 => -39,
    39756 => -39,
    39757 => -39,
    39758 => -39,
    39759 => -39,
    39760 => -39,
    39761 => -39,
    39762 => -39,
    39763 => -39,
    39764 => -39,
    39765 => -39,
    39766 => -39,
    39767 => -39,
    39768 => -39,
    39769 => -39,
    39770 => -39,
    39771 => -39,
    39772 => -39,
    39773 => -39,
    39774 => -39,
    39775 => -39,
    39776 => -39,
    39777 => -39,
    39778 => -39,
    39779 => -39,
    39780 => -39,
    39781 => -39,
    39782 => -39,
    39783 => -39,
    39784 => -39,
    39785 => -39,
    39786 => -39,
    39787 => -39,
    39788 => -39,
    39789 => -39,
    39790 => -39,
    39791 => -39,
    39792 => -39,
    39793 => -39,
    39794 => -39,
    39795 => -39,
    39796 => -39,
    39797 => -39,
    39798 => -39,
    39799 => -39,
    39800 => -39,
    39801 => -39,
    39802 => -39,
    39803 => -39,
    39804 => -39,
    39805 => -39,
    39806 => -39,
    39807 => -39,
    39808 => -39,
    39809 => -39,
    39810 => -39,
    39811 => -39,
    39812 => -39,
    39813 => -39,
    39814 => -39,
    39815 => -39,
    39816 => -39,
    39817 => -39,
    39818 => -39,
    39819 => -39,
    39820 => -39,
    39821 => -39,
    39822 => -39,
    39823 => -39,
    39824 => -39,
    39825 => -39,
    39826 => -39,
    39827 => -39,
    39828 => -39,
    39829 => -39,
    39830 => -39,
    39831 => -39,
    39832 => -39,
    39833 => -39,
    39834 => -39,
    39835 => -39,
    39836 => -39,
    39837 => -40,
    39838 => -40,
    39839 => -40,
    39840 => -40,
    39841 => -40,
    39842 => -40,
    39843 => -40,
    39844 => -40,
    39845 => -40,
    39846 => -40,
    39847 => -40,
    39848 => -40,
    39849 => -40,
    39850 => -40,
    39851 => -40,
    39852 => -40,
    39853 => -40,
    39854 => -40,
    39855 => -40,
    39856 => -40,
    39857 => -40,
    39858 => -40,
    39859 => -40,
    39860 => -40,
    39861 => -40,
    39862 => -40,
    39863 => -40,
    39864 => -40,
    39865 => -40,
    39866 => -40,
    39867 => -40,
    39868 => -40,
    39869 => -40,
    39870 => -40,
    39871 => -40,
    39872 => -40,
    39873 => -40,
    39874 => -40,
    39875 => -40,
    39876 => -40,
    39877 => -40,
    39878 => -40,
    39879 => -40,
    39880 => -40,
    39881 => -40,
    39882 => -40,
    39883 => -40,
    39884 => -40,
    39885 => -40,
    39886 => -40,
    39887 => -40,
    39888 => -40,
    39889 => -40,
    39890 => -40,
    39891 => -40,
    39892 => -40,
    39893 => -40,
    39894 => -40,
    39895 => -40,
    39896 => -40,
    39897 => -40,
    39898 => -40,
    39899 => -40,
    39900 => -40,
    39901 => -40,
    39902 => -40,
    39903 => -40,
    39904 => -40,
    39905 => -40,
    39906 => -40,
    39907 => -40,
    39908 => -40,
    39909 => -40,
    39910 => -40,
    39911 => -40,
    39912 => -40,
    39913 => -40,
    39914 => -40,
    39915 => -40,
    39916 => -40,
    39917 => -40,
    39918 => -40,
    39919 => -40,
    39920 => -40,
    39921 => -40,
    39922 => -40,
    39923 => -40,
    39924 => -40,
    39925 => -40,
    39926 => -40,
    39927 => -40,
    39928 => -40,
    39929 => -40,
    39930 => -40,
    39931 => -40,
    39932 => -40,
    39933 => -40,
    39934 => -40,
    39935 => -40,
    39936 => -40,
    39937 => -40,
    39938 => -40,
    39939 => -40,
    39940 => -40,
    39941 => -40,
    39942 => -40,
    39943 => -40,
    39944 => -40,
    39945 => -40,
    39946 => -40,
    39947 => -40,
    39948 => -40,
    39949 => -40,
    39950 => -40,
    39951 => -40,
    39952 => -40,
    39953 => -40,
    39954 => -40,
    39955 => -40,
    39956 => -40,
    39957 => -40,
    39958 => -40,
    39959 => -40,
    39960 => -40,
    39961 => -40,
    39962 => -40,
    39963 => -40,
    39964 => -40,
    39965 => -40,
    39966 => -40,
    39967 => -40,
    39968 => -40,
    39969 => -40,
    39970 => -40,
    39971 => -40,
    39972 => -40,
    39973 => -40,
    39974 => -40,
    39975 => -40,
    39976 => -40,
    39977 => -40,
    39978 => -40,
    39979 => -40,
    39980 => -40,
    39981 => -40,
    39982 => -40,
    39983 => -40,
    39984 => -40,
    39985 => -40,
    39986 => -40,
    39987 => -40,
    39988 => -40,
    39989 => -40,
    39990 => -40,
    39991 => -40,
    39992 => -40,
    39993 => -40,
    39994 => -40,
    39995 => -40,
    39996 => -40,
    39997 => -40,
    39998 => -40,
    39999 => -40,
    40000 => -40,
    40001 => -40,
    40002 => -40,
    40003 => -40,
    40004 => -40,
    40005 => -40,
    40006 => -40,
    40007 => -40,
    40008 => -40,
    40009 => -40,
    40010 => -40,
    40011 => -40,
    40012 => -40,
    40013 => -40,
    40014 => -40,
    40015 => -40,
    40016 => -40,
    40017 => -40,
    40018 => -40,
    40019 => -40,
    40020 => -40,
    40021 => -40,
    40022 => -40,
    40023 => -40,
    40024 => -40,
    40025 => -40,
    40026 => -40,
    40027 => -40,
    40028 => -40,
    40029 => -40,
    40030 => -40,
    40031 => -40,
    40032 => -40,
    40033 => -40,
    40034 => -40,
    40035 => -40,
    40036 => -40,
    40037 => -40,
    40038 => -40,
    40039 => -40,
    40040 => -40,
    40041 => -40,
    40042 => -40,
    40043 => -40,
    40044 => -40,
    40045 => -40,
    40046 => -40,
    40047 => -40,
    40048 => -40,
    40049 => -40,
    40050 => -40,
    40051 => -41,
    40052 => -41,
    40053 => -41,
    40054 => -41,
    40055 => -41,
    40056 => -41,
    40057 => -41,
    40058 => -41,
    40059 => -41,
    40060 => -41,
    40061 => -41,
    40062 => -41,
    40063 => -41,
    40064 => -41,
    40065 => -41,
    40066 => -41,
    40067 => -41,
    40068 => -41,
    40069 => -41,
    40070 => -41,
    40071 => -41,
    40072 => -41,
    40073 => -41,
    40074 => -41,
    40075 => -41,
    40076 => -41,
    40077 => -41,
    40078 => -41,
    40079 => -41,
    40080 => -41,
    40081 => -41,
    40082 => -41,
    40083 => -41,
    40084 => -41,
    40085 => -41,
    40086 => -41,
    40087 => -41,
    40088 => -41,
    40089 => -41,
    40090 => -41,
    40091 => -41,
    40092 => -41,
    40093 => -41,
    40094 => -41,
    40095 => -41,
    40096 => -41,
    40097 => -41,
    40098 => -41,
    40099 => -41,
    40100 => -41,
    40101 => -41,
    40102 => -41,
    40103 => -41,
    40104 => -41,
    40105 => -41,
    40106 => -41,
    40107 => -41,
    40108 => -41,
    40109 => -41,
    40110 => -41,
    40111 => -41,
    40112 => -41,
    40113 => -41,
    40114 => -41,
    40115 => -41,
    40116 => -41,
    40117 => -41,
    40118 => -41,
    40119 => -41,
    40120 => -41,
    40121 => -41,
    40122 => -41,
    40123 => -41,
    40124 => -41,
    40125 => -41,
    40126 => -41,
    40127 => -41,
    40128 => -41,
    40129 => -41,
    40130 => -41,
    40131 => -41,
    40132 => -41,
    40133 => -41,
    40134 => -41,
    40135 => -41,
    40136 => -41,
    40137 => -41,
    40138 => -41,
    40139 => -41,
    40140 => -41,
    40141 => -41,
    40142 => -41,
    40143 => -41,
    40144 => -41,
    40145 => -41,
    40146 => -41,
    40147 => -41,
    40148 => -41,
    40149 => -41,
    40150 => -41,
    40151 => -41,
    40152 => -41,
    40153 => -41,
    40154 => -41,
    40155 => -41,
    40156 => -41,
    40157 => -41,
    40158 => -41,
    40159 => -41,
    40160 => -41,
    40161 => -41,
    40162 => -41,
    40163 => -41,
    40164 => -41,
    40165 => -41,
    40166 => -41,
    40167 => -41,
    40168 => -41,
    40169 => -41,
    40170 => -41,
    40171 => -41,
    40172 => -41,
    40173 => -41,
    40174 => -41,
    40175 => -41,
    40176 => -41,
    40177 => -41,
    40178 => -41,
    40179 => -41,
    40180 => -41,
    40181 => -41,
    40182 => -41,
    40183 => -41,
    40184 => -41,
    40185 => -41,
    40186 => -41,
    40187 => -41,
    40188 => -41,
    40189 => -41,
    40190 => -41,
    40191 => -41,
    40192 => -41,
    40193 => -41,
    40194 => -41,
    40195 => -41,
    40196 => -41,
    40197 => -41,
    40198 => -41,
    40199 => -41,
    40200 => -41,
    40201 => -41,
    40202 => -41,
    40203 => -41,
    40204 => -41,
    40205 => -41,
    40206 => -41,
    40207 => -41,
    40208 => -41,
    40209 => -41,
    40210 => -41,
    40211 => -41,
    40212 => -41,
    40213 => -41,
    40214 => -41,
    40215 => -41,
    40216 => -41,
    40217 => -41,
    40218 => -41,
    40219 => -41,
    40220 => -41,
    40221 => -41,
    40222 => -41,
    40223 => -41,
    40224 => -41,
    40225 => -41,
    40226 => -41,
    40227 => -41,
    40228 => -41,
    40229 => -41,
    40230 => -41,
    40231 => -41,
    40232 => -41,
    40233 => -41,
    40234 => -41,
    40235 => -41,
    40236 => -41,
    40237 => -41,
    40238 => -41,
    40239 => -41,
    40240 => -41,
    40241 => -41,
    40242 => -41,
    40243 => -41,
    40244 => -41,
    40245 => -41,
    40246 => -41,
    40247 => -41,
    40248 => -41,
    40249 => -41,
    40250 => -41,
    40251 => -41,
    40252 => -41,
    40253 => -41,
    40254 => -41,
    40255 => -41,
    40256 => -41,
    40257 => -41,
    40258 => -41,
    40259 => -41,
    40260 => -41,
    40261 => -41,
    40262 => -41,
    40263 => -41,
    40264 => -41,
    40265 => -41,
    40266 => -41,
    40267 => -41,
    40268 => -41,
    40269 => -42,
    40270 => -42,
    40271 => -42,
    40272 => -42,
    40273 => -42,
    40274 => -42,
    40275 => -42,
    40276 => -42,
    40277 => -42,
    40278 => -42,
    40279 => -42,
    40280 => -42,
    40281 => -42,
    40282 => -42,
    40283 => -42,
    40284 => -42,
    40285 => -42,
    40286 => -42,
    40287 => -42,
    40288 => -42,
    40289 => -42,
    40290 => -42,
    40291 => -42,
    40292 => -42,
    40293 => -42,
    40294 => -42,
    40295 => -42,
    40296 => -42,
    40297 => -42,
    40298 => -42,
    40299 => -42,
    40300 => -42,
    40301 => -42,
    40302 => -42,
    40303 => -42,
    40304 => -42,
    40305 => -42,
    40306 => -42,
    40307 => -42,
    40308 => -42,
    40309 => -42,
    40310 => -42,
    40311 => -42,
    40312 => -42,
    40313 => -42,
    40314 => -42,
    40315 => -42,
    40316 => -42,
    40317 => -42,
    40318 => -42,
    40319 => -42,
    40320 => -42,
    40321 => -42,
    40322 => -42,
    40323 => -42,
    40324 => -42,
    40325 => -42,
    40326 => -42,
    40327 => -42,
    40328 => -42,
    40329 => -42,
    40330 => -42,
    40331 => -42,
    40332 => -42,
    40333 => -42,
    40334 => -42,
    40335 => -42,
    40336 => -42,
    40337 => -42,
    40338 => -42,
    40339 => -42,
    40340 => -42,
    40341 => -42,
    40342 => -42,
    40343 => -42,
    40344 => -42,
    40345 => -42,
    40346 => -42,
    40347 => -42,
    40348 => -42,
    40349 => -42,
    40350 => -42,
    40351 => -42,
    40352 => -42,
    40353 => -42,
    40354 => -42,
    40355 => -42,
    40356 => -42,
    40357 => -42,
    40358 => -42,
    40359 => -42,
    40360 => -42,
    40361 => -42,
    40362 => -42,
    40363 => -42,
    40364 => -42,
    40365 => -42,
    40366 => -42,
    40367 => -42,
    40368 => -42,
    40369 => -42,
    40370 => -42,
    40371 => -42,
    40372 => -42,
    40373 => -42,
    40374 => -42,
    40375 => -42,
    40376 => -42,
    40377 => -42,
    40378 => -42,
    40379 => -42,
    40380 => -42,
    40381 => -42,
    40382 => -42,
    40383 => -42,
    40384 => -42,
    40385 => -42,
    40386 => -42,
    40387 => -42,
    40388 => -42,
    40389 => -42,
    40390 => -42,
    40391 => -42,
    40392 => -42,
    40393 => -42,
    40394 => -42,
    40395 => -42,
    40396 => -42,
    40397 => -42,
    40398 => -42,
    40399 => -42,
    40400 => -42,
    40401 => -42,
    40402 => -42,
    40403 => -42,
    40404 => -42,
    40405 => -42,
    40406 => -42,
    40407 => -42,
    40408 => -42,
    40409 => -42,
    40410 => -42,
    40411 => -42,
    40412 => -42,
    40413 => -42,
    40414 => -42,
    40415 => -42,
    40416 => -42,
    40417 => -42,
    40418 => -42,
    40419 => -42,
    40420 => -42,
    40421 => -42,
    40422 => -42,
    40423 => -42,
    40424 => -42,
    40425 => -42,
    40426 => -42,
    40427 => -42,
    40428 => -42,
    40429 => -42,
    40430 => -42,
    40431 => -42,
    40432 => -42,
    40433 => -42,
    40434 => -42,
    40435 => -42,
    40436 => -42,
    40437 => -42,
    40438 => -42,
    40439 => -42,
    40440 => -42,
    40441 => -42,
    40442 => -42,
    40443 => -42,
    40444 => -42,
    40445 => -42,
    40446 => -42,
    40447 => -42,
    40448 => -42,
    40449 => -42,
    40450 => -42,
    40451 => -42,
    40452 => -42,
    40453 => -42,
    40454 => -42,
    40455 => -42,
    40456 => -42,
    40457 => -42,
    40458 => -42,
    40459 => -42,
    40460 => -42,
    40461 => -42,
    40462 => -42,
    40463 => -42,
    40464 => -42,
    40465 => -42,
    40466 => -42,
    40467 => -42,
    40468 => -42,
    40469 => -42,
    40470 => -42,
    40471 => -42,
    40472 => -42,
    40473 => -42,
    40474 => -42,
    40475 => -42,
    40476 => -42,
    40477 => -42,
    40478 => -42,
    40479 => -42,
    40480 => -42,
    40481 => -42,
    40482 => -42,
    40483 => -42,
    40484 => -42,
    40485 => -42,
    40486 => -42,
    40487 => -42,
    40488 => -42,
    40489 => -42,
    40490 => -42,
    40491 => -43,
    40492 => -43,
    40493 => -43,
    40494 => -43,
    40495 => -43,
    40496 => -43,
    40497 => -43,
    40498 => -43,
    40499 => -43,
    40500 => -43,
    40501 => -43,
    40502 => -43,
    40503 => -43,
    40504 => -43,
    40505 => -43,
    40506 => -43,
    40507 => -43,
    40508 => -43,
    40509 => -43,
    40510 => -43,
    40511 => -43,
    40512 => -43,
    40513 => -43,
    40514 => -43,
    40515 => -43,
    40516 => -43,
    40517 => -43,
    40518 => -43,
    40519 => -43,
    40520 => -43,
    40521 => -43,
    40522 => -43,
    40523 => -43,
    40524 => -43,
    40525 => -43,
    40526 => -43,
    40527 => -43,
    40528 => -43,
    40529 => -43,
    40530 => -43,
    40531 => -43,
    40532 => -43,
    40533 => -43,
    40534 => -43,
    40535 => -43,
    40536 => -43,
    40537 => -43,
    40538 => -43,
    40539 => -43,
    40540 => -43,
    40541 => -43,
    40542 => -43,
    40543 => -43,
    40544 => -43,
    40545 => -43,
    40546 => -43,
    40547 => -43,
    40548 => -43,
    40549 => -43,
    40550 => -43,
    40551 => -43,
    40552 => -43,
    40553 => -43,
    40554 => -43,
    40555 => -43,
    40556 => -43,
    40557 => -43,
    40558 => -43,
    40559 => -43,
    40560 => -43,
    40561 => -43,
    40562 => -43,
    40563 => -43,
    40564 => -43,
    40565 => -43,
    40566 => -43,
    40567 => -43,
    40568 => -43,
    40569 => -43,
    40570 => -43,
    40571 => -43,
    40572 => -43,
    40573 => -43,
    40574 => -43,
    40575 => -43,
    40576 => -43,
    40577 => -43,
    40578 => -43,
    40579 => -43,
    40580 => -43,
    40581 => -43,
    40582 => -43,
    40583 => -43,
    40584 => -43,
    40585 => -43,
    40586 => -43,
    40587 => -43,
    40588 => -43,
    40589 => -43,
    40590 => -43,
    40591 => -43,
    40592 => -43,
    40593 => -43,
    40594 => -43,
    40595 => -43,
    40596 => -43,
    40597 => -43,
    40598 => -43,
    40599 => -43,
    40600 => -43,
    40601 => -43,
    40602 => -43,
    40603 => -43,
    40604 => -43,
    40605 => -43,
    40606 => -43,
    40607 => -43,
    40608 => -43,
    40609 => -43,
    40610 => -43,
    40611 => -43,
    40612 => -43,
    40613 => -43,
    40614 => -43,
    40615 => -43,
    40616 => -43,
    40617 => -43,
    40618 => -43,
    40619 => -43,
    40620 => -43,
    40621 => -43,
    40622 => -43,
    40623 => -43,
    40624 => -43,
    40625 => -43,
    40626 => -43,
    40627 => -43,
    40628 => -43,
    40629 => -43,
    40630 => -43,
    40631 => -43,
    40632 => -43,
    40633 => -43,
    40634 => -43,
    40635 => -43,
    40636 => -43,
    40637 => -43,
    40638 => -43,
    40639 => -43,
    40640 => -43,
    40641 => -43,
    40642 => -43,
    40643 => -43,
    40644 => -43,
    40645 => -43,
    40646 => -43,
    40647 => -43,
    40648 => -43,
    40649 => -43,
    40650 => -43,
    40651 => -43,
    40652 => -43,
    40653 => -43,
    40654 => -43,
    40655 => -43,
    40656 => -43,
    40657 => -43,
    40658 => -43,
    40659 => -43,
    40660 => -43,
    40661 => -43,
    40662 => -43,
    40663 => -43,
    40664 => -43,
    40665 => -43,
    40666 => -43,
    40667 => -43,
    40668 => -43,
    40669 => -43,
    40670 => -43,
    40671 => -43,
    40672 => -43,
    40673 => -43,
    40674 => -43,
    40675 => -43,
    40676 => -43,
    40677 => -43,
    40678 => -43,
    40679 => -43,
    40680 => -43,
    40681 => -43,
    40682 => -43,
    40683 => -43,
    40684 => -43,
    40685 => -43,
    40686 => -43,
    40687 => -43,
    40688 => -43,
    40689 => -43,
    40690 => -43,
    40691 => -43,
    40692 => -43,
    40693 => -43,
    40694 => -43,
    40695 => -43,
    40696 => -43,
    40697 => -43,
    40698 => -43,
    40699 => -43,
    40700 => -43,
    40701 => -43,
    40702 => -43,
    40703 => -43,
    40704 => -43,
    40705 => -43,
    40706 => -43,
    40707 => -43,
    40708 => -43,
    40709 => -43,
    40710 => -43,
    40711 => -43,
    40712 => -43,
    40713 => -43,
    40714 => -43,
    40715 => -43,
    40716 => -43,
    40717 => -43,
    40718 => -44,
    40719 => -44,
    40720 => -44,
    40721 => -44,
    40722 => -44,
    40723 => -44,
    40724 => -44,
    40725 => -44,
    40726 => -44,
    40727 => -44,
    40728 => -44,
    40729 => -44,
    40730 => -44,
    40731 => -44,
    40732 => -44,
    40733 => -44,
    40734 => -44,
    40735 => -44,
    40736 => -44,
    40737 => -44,
    40738 => -44,
    40739 => -44,
    40740 => -44,
    40741 => -44,
    40742 => -44,
    40743 => -44,
    40744 => -44,
    40745 => -44,
    40746 => -44,
    40747 => -44,
    40748 => -44,
    40749 => -44,
    40750 => -44,
    40751 => -44,
    40752 => -44,
    40753 => -44,
    40754 => -44,
    40755 => -44,
    40756 => -44,
    40757 => -44,
    40758 => -44,
    40759 => -44,
    40760 => -44,
    40761 => -44,
    40762 => -44,
    40763 => -44,
    40764 => -44,
    40765 => -44,
    40766 => -44,
    40767 => -44,
    40768 => -44,
    40769 => -44,
    40770 => -44,
    40771 => -44,
    40772 => -44,
    40773 => -44,
    40774 => -44,
    40775 => -44,
    40776 => -44,
    40777 => -44,
    40778 => -44,
    40779 => -44,
    40780 => -44,
    40781 => -44,
    40782 => -44,
    40783 => -44,
    40784 => -44,
    40785 => -44,
    40786 => -44,
    40787 => -44,
    40788 => -44,
    40789 => -44,
    40790 => -44,
    40791 => -44,
    40792 => -44,
    40793 => -44,
    40794 => -44,
    40795 => -44,
    40796 => -44,
    40797 => -44,
    40798 => -44,
    40799 => -44,
    40800 => -44,
    40801 => -44,
    40802 => -44,
    40803 => -44,
    40804 => -44,
    40805 => -44,
    40806 => -44,
    40807 => -44,
    40808 => -44,
    40809 => -44,
    40810 => -44,
    40811 => -44,
    40812 => -44,
    40813 => -44,
    40814 => -44,
    40815 => -44,
    40816 => -44,
    40817 => -44,
    40818 => -44,
    40819 => -44,
    40820 => -44,
    40821 => -44,
    40822 => -44,
    40823 => -44,
    40824 => -44,
    40825 => -44,
    40826 => -44,
    40827 => -44,
    40828 => -44,
    40829 => -44,
    40830 => -44,
    40831 => -44,
    40832 => -44,
    40833 => -44,
    40834 => -44,
    40835 => -44,
    40836 => -44,
    40837 => -44,
    40838 => -44,
    40839 => -44,
    40840 => -44,
    40841 => -44,
    40842 => -44,
    40843 => -44,
    40844 => -44,
    40845 => -44,
    40846 => -44,
    40847 => -44,
    40848 => -44,
    40849 => -44,
    40850 => -44,
    40851 => -44,
    40852 => -44,
    40853 => -44,
    40854 => -44,
    40855 => -44,
    40856 => -44,
    40857 => -44,
    40858 => -44,
    40859 => -44,
    40860 => -44,
    40861 => -44,
    40862 => -44,
    40863 => -44,
    40864 => -44,
    40865 => -44,
    40866 => -44,
    40867 => -44,
    40868 => -44,
    40869 => -44,
    40870 => -44,
    40871 => -44,
    40872 => -44,
    40873 => -44,
    40874 => -44,
    40875 => -44,
    40876 => -44,
    40877 => -44,
    40878 => -44,
    40879 => -44,
    40880 => -44,
    40881 => -44,
    40882 => -44,
    40883 => -44,
    40884 => -44,
    40885 => -44,
    40886 => -44,
    40887 => -44,
    40888 => -44,
    40889 => -44,
    40890 => -44,
    40891 => -44,
    40892 => -44,
    40893 => -44,
    40894 => -44,
    40895 => -44,
    40896 => -44,
    40897 => -44,
    40898 => -44,
    40899 => -44,
    40900 => -44,
    40901 => -44,
    40902 => -44,
    40903 => -44,
    40904 => -44,
    40905 => -44,
    40906 => -44,
    40907 => -44,
    40908 => -44,
    40909 => -44,
    40910 => -44,
    40911 => -44,
    40912 => -44,
    40913 => -44,
    40914 => -44,
    40915 => -44,
    40916 => -44,
    40917 => -44,
    40918 => -44,
    40919 => -44,
    40920 => -44,
    40921 => -44,
    40922 => -44,
    40923 => -44,
    40924 => -44,
    40925 => -44,
    40926 => -44,
    40927 => -44,
    40928 => -44,
    40929 => -44,
    40930 => -44,
    40931 => -44,
    40932 => -44,
    40933 => -44,
    40934 => -44,
    40935 => -44,
    40936 => -44,
    40937 => -44,
    40938 => -44,
    40939 => -44,
    40940 => -44,
    40941 => -44,
    40942 => -44,
    40943 => -44,
    40944 => -44,
    40945 => -44,
    40946 => -44,
    40947 => -44,
    40948 => -44,
    40949 => -45,
    40950 => -45,
    40951 => -45,
    40952 => -45,
    40953 => -45,
    40954 => -45,
    40955 => -45,
    40956 => -45,
    40957 => -45,
    40958 => -45,
    40959 => -45,
    40960 => -45,
    40961 => -45,
    40962 => -45,
    40963 => -45,
    40964 => -45,
    40965 => -45,
    40966 => -45,
    40967 => -45,
    40968 => -45,
    40969 => -45,
    40970 => -45,
    40971 => -45,
    40972 => -45,
    40973 => -45,
    40974 => -45,
    40975 => -45,
    40976 => -45,
    40977 => -45,
    40978 => -45,
    40979 => -45,
    40980 => -45,
    40981 => -45,
    40982 => -45,
    40983 => -45,
    40984 => -45,
    40985 => -45,
    40986 => -45,
    40987 => -45,
    40988 => -45,
    40989 => -45,
    40990 => -45,
    40991 => -45,
    40992 => -45,
    40993 => -45,
    40994 => -45,
    40995 => -45,
    40996 => -45,
    40997 => -45,
    40998 => -45,
    40999 => -45,
    41000 => -45,
    41001 => -45,
    41002 => -45,
    41003 => -45,
    41004 => -45,
    41005 => -45,
    41006 => -45,
    41007 => -45,
    41008 => -45,
    41009 => -45,
    41010 => -45,
    41011 => -45,
    41012 => -45,
    41013 => -45,
    41014 => -45,
    41015 => -45,
    41016 => -45,
    41017 => -45,
    41018 => -45,
    41019 => -45,
    41020 => -45,
    41021 => -45,
    41022 => -45,
    41023 => -45,
    41024 => -45,
    41025 => -45,
    41026 => -45,
    41027 => -45,
    41028 => -45,
    41029 => -45,
    41030 => -45,
    41031 => -45,
    41032 => -45,
    41033 => -45,
    41034 => -45,
    41035 => -45,
    41036 => -45,
    41037 => -45,
    41038 => -45,
    41039 => -45,
    41040 => -45,
    41041 => -45,
    41042 => -45,
    41043 => -45,
    41044 => -45,
    41045 => -45,
    41046 => -45,
    41047 => -45,
    41048 => -45,
    41049 => -45,
    41050 => -45,
    41051 => -45,
    41052 => -45,
    41053 => -45,
    41054 => -45,
    41055 => -45,
    41056 => -45,
    41057 => -45,
    41058 => -45,
    41059 => -45,
    41060 => -45,
    41061 => -45,
    41062 => -45,
    41063 => -45,
    41064 => -45,
    41065 => -45,
    41066 => -45,
    41067 => -45,
    41068 => -45,
    41069 => -45,
    41070 => -45,
    41071 => -45,
    41072 => -45,
    41073 => -45,
    41074 => -45,
    41075 => -45,
    41076 => -45,
    41077 => -45,
    41078 => -45,
    41079 => -45,
    41080 => -45,
    41081 => -45,
    41082 => -45,
    41083 => -45,
    41084 => -45,
    41085 => -45,
    41086 => -45,
    41087 => -45,
    41088 => -45,
    41089 => -45,
    41090 => -45,
    41091 => -45,
    41092 => -45,
    41093 => -45,
    41094 => -45,
    41095 => -45,
    41096 => -45,
    41097 => -45,
    41098 => -45,
    41099 => -45,
    41100 => -45,
    41101 => -45,
    41102 => -45,
    41103 => -45,
    41104 => -45,
    41105 => -45,
    41106 => -45,
    41107 => -45,
    41108 => -45,
    41109 => -45,
    41110 => -45,
    41111 => -45,
    41112 => -45,
    41113 => -45,
    41114 => -45,
    41115 => -45,
    41116 => -45,
    41117 => -45,
    41118 => -45,
    41119 => -45,
    41120 => -45,
    41121 => -45,
    41122 => -45,
    41123 => -45,
    41124 => -45,
    41125 => -45,
    41126 => -45,
    41127 => -45,
    41128 => -45,
    41129 => -45,
    41130 => -45,
    41131 => -45,
    41132 => -45,
    41133 => -45,
    41134 => -45,
    41135 => -45,
    41136 => -45,
    41137 => -45,
    41138 => -45,
    41139 => -45,
    41140 => -45,
    41141 => -45,
    41142 => -45,
    41143 => -45,
    41144 => -45,
    41145 => -45,
    41146 => -45,
    41147 => -45,
    41148 => -45,
    41149 => -45,
    41150 => -45,
    41151 => -45,
    41152 => -45,
    41153 => -45,
    41154 => -45,
    41155 => -45,
    41156 => -45,
    41157 => -45,
    41158 => -45,
    41159 => -45,
    41160 => -45,
    41161 => -45,
    41162 => -45,
    41163 => -45,
    41164 => -45,
    41165 => -45,
    41166 => -45,
    41167 => -45,
    41168 => -45,
    41169 => -45,
    41170 => -45,
    41171 => -45,
    41172 => -45,
    41173 => -45,
    41174 => -45,
    41175 => -45,
    41176 => -45,
    41177 => -45,
    41178 => -45,
    41179 => -45,
    41180 => -45,
    41181 => -45,
    41182 => -45,
    41183 => -45,
    41184 => -45,
    41185 => -45,
    41186 => -46,
    41187 => -46,
    41188 => -46,
    41189 => -46,
    41190 => -46,
    41191 => -46,
    41192 => -46,
    41193 => -46,
    41194 => -46,
    41195 => -46,
    41196 => -46,
    41197 => -46,
    41198 => -46,
    41199 => -46,
    41200 => -46,
    41201 => -46,
    41202 => -46,
    41203 => -46,
    41204 => -46,
    41205 => -46,
    41206 => -46,
    41207 => -46,
    41208 => -46,
    41209 => -46,
    41210 => -46,
    41211 => -46,
    41212 => -46,
    41213 => -46,
    41214 => -46,
    41215 => -46,
    41216 => -46,
    41217 => -46,
    41218 => -46,
    41219 => -46,
    41220 => -46,
    41221 => -46,
    41222 => -46,
    41223 => -46,
    41224 => -46,
    41225 => -46,
    41226 => -46,
    41227 => -46,
    41228 => -46,
    41229 => -46,
    41230 => -46,
    41231 => -46,
    41232 => -46,
    41233 => -46,
    41234 => -46,
    41235 => -46,
    41236 => -46,
    41237 => -46,
    41238 => -46,
    41239 => -46,
    41240 => -46,
    41241 => -46,
    41242 => -46,
    41243 => -46,
    41244 => -46,
    41245 => -46,
    41246 => -46,
    41247 => -46,
    41248 => -46,
    41249 => -46,
    41250 => -46,
    41251 => -46,
    41252 => -46,
    41253 => -46,
    41254 => -46,
    41255 => -46,
    41256 => -46,
    41257 => -46,
    41258 => -46,
    41259 => -46,
    41260 => -46,
    41261 => -46,
    41262 => -46,
    41263 => -46,
    41264 => -46,
    41265 => -46,
    41266 => -46,
    41267 => -46,
    41268 => -46,
    41269 => -46,
    41270 => -46,
    41271 => -46,
    41272 => -46,
    41273 => -46,
    41274 => -46,
    41275 => -46,
    41276 => -46,
    41277 => -46,
    41278 => -46,
    41279 => -46,
    41280 => -46,
    41281 => -46,
    41282 => -46,
    41283 => -46,
    41284 => -46,
    41285 => -46,
    41286 => -46,
    41287 => -46,
    41288 => -46,
    41289 => -46,
    41290 => -46,
    41291 => -46,
    41292 => -46,
    41293 => -46,
    41294 => -46,
    41295 => -46,
    41296 => -46,
    41297 => -46,
    41298 => -46,
    41299 => -46,
    41300 => -46,
    41301 => -46,
    41302 => -46,
    41303 => -46,
    41304 => -46,
    41305 => -46,
    41306 => -46,
    41307 => -46,
    41308 => -46,
    41309 => -46,
    41310 => -46,
    41311 => -46,
    41312 => -46,
    41313 => -46,
    41314 => -46,
    41315 => -46,
    41316 => -46,
    41317 => -46,
    41318 => -46,
    41319 => -46,
    41320 => -46,
    41321 => -46,
    41322 => -46,
    41323 => -46,
    41324 => -46,
    41325 => -46,
    41326 => -46,
    41327 => -46,
    41328 => -46,
    41329 => -46,
    41330 => -46,
    41331 => -46,
    41332 => -46,
    41333 => -46,
    41334 => -46,
    41335 => -46,
    41336 => -46,
    41337 => -46,
    41338 => -46,
    41339 => -46,
    41340 => -46,
    41341 => -46,
    41342 => -46,
    41343 => -46,
    41344 => -46,
    41345 => -46,
    41346 => -46,
    41347 => -46,
    41348 => -46,
    41349 => -46,
    41350 => -46,
    41351 => -46,
    41352 => -46,
    41353 => -46,
    41354 => -46,
    41355 => -46,
    41356 => -46,
    41357 => -46,
    41358 => -46,
    41359 => -46,
    41360 => -46,
    41361 => -46,
    41362 => -46,
    41363 => -46,
    41364 => -46,
    41365 => -46,
    41366 => -46,
    41367 => -46,
    41368 => -46,
    41369 => -46,
    41370 => -46,
    41371 => -46,
    41372 => -46,
    41373 => -46,
    41374 => -46,
    41375 => -46,
    41376 => -46,
    41377 => -46,
    41378 => -46,
    41379 => -46,
    41380 => -46,
    41381 => -46,
    41382 => -46,
    41383 => -46,
    41384 => -46,
    41385 => -46,
    41386 => -46,
    41387 => -46,
    41388 => -46,
    41389 => -46,
    41390 => -46,
    41391 => -46,
    41392 => -46,
    41393 => -46,
    41394 => -46,
    41395 => -46,
    41396 => -46,
    41397 => -46,
    41398 => -46,
    41399 => -46,
    41400 => -46,
    41401 => -46,
    41402 => -46,
    41403 => -46,
    41404 => -46,
    41405 => -46,
    41406 => -46,
    41407 => -46,
    41408 => -46,
    41409 => -46,
    41410 => -46,
    41411 => -46,
    41412 => -46,
    41413 => -46,
    41414 => -46,
    41415 => -46,
    41416 => -46,
    41417 => -46,
    41418 => -46,
    41419 => -46,
    41420 => -46,
    41421 => -46,
    41422 => -46,
    41423 => -46,
    41424 => -46,
    41425 => -46,
    41426 => -46,
    41427 => -46,
    41428 => -47,
    41429 => -47,
    41430 => -47,
    41431 => -47,
    41432 => -47,
    41433 => -47,
    41434 => -47,
    41435 => -47,
    41436 => -47,
    41437 => -47,
    41438 => -47,
    41439 => -47,
    41440 => -47,
    41441 => -47,
    41442 => -47,
    41443 => -47,
    41444 => -47,
    41445 => -47,
    41446 => -47,
    41447 => -47,
    41448 => -47,
    41449 => -47,
    41450 => -47,
    41451 => -47,
    41452 => -47,
    41453 => -47,
    41454 => -47,
    41455 => -47,
    41456 => -47,
    41457 => -47,
    41458 => -47,
    41459 => -47,
    41460 => -47,
    41461 => -47,
    41462 => -47,
    41463 => -47,
    41464 => -47,
    41465 => -47,
    41466 => -47,
    41467 => -47,
    41468 => -47,
    41469 => -47,
    41470 => -47,
    41471 => -47,
    41472 => -47,
    41473 => -47,
    41474 => -47,
    41475 => -47,
    41476 => -47,
    41477 => -47,
    41478 => -47,
    41479 => -47,
    41480 => -47,
    41481 => -47,
    41482 => -47,
    41483 => -47,
    41484 => -47,
    41485 => -47,
    41486 => -47,
    41487 => -47,
    41488 => -47,
    41489 => -47,
    41490 => -47,
    41491 => -47,
    41492 => -47,
    41493 => -47,
    41494 => -47,
    41495 => -47,
    41496 => -47,
    41497 => -47,
    41498 => -47,
    41499 => -47,
    41500 => -47,
    41501 => -47,
    41502 => -47,
    41503 => -47,
    41504 => -47,
    41505 => -47,
    41506 => -47,
    41507 => -47,
    41508 => -47,
    41509 => -47,
    41510 => -47,
    41511 => -47,
    41512 => -47,
    41513 => -47,
    41514 => -47,
    41515 => -47,
    41516 => -47,
    41517 => -47,
    41518 => -47,
    41519 => -47,
    41520 => -47,
    41521 => -47,
    41522 => -47,
    41523 => -47,
    41524 => -47,
    41525 => -47,
    41526 => -47,
    41527 => -47,
    41528 => -47,
    41529 => -47,
    41530 => -47,
    41531 => -47,
    41532 => -47,
    41533 => -47,
    41534 => -47,
    41535 => -47,
    41536 => -47,
    41537 => -47,
    41538 => -47,
    41539 => -47,
    41540 => -47,
    41541 => -47,
    41542 => -47,
    41543 => -47,
    41544 => -47,
    41545 => -47,
    41546 => -47,
    41547 => -47,
    41548 => -47,
    41549 => -47,
    41550 => -47,
    41551 => -47,
    41552 => -47,
    41553 => -47,
    41554 => -47,
    41555 => -47,
    41556 => -47,
    41557 => -47,
    41558 => -47,
    41559 => -47,
    41560 => -47,
    41561 => -47,
    41562 => -47,
    41563 => -47,
    41564 => -47,
    41565 => -47,
    41566 => -47,
    41567 => -47,
    41568 => -47,
    41569 => -47,
    41570 => -47,
    41571 => -47,
    41572 => -47,
    41573 => -47,
    41574 => -47,
    41575 => -47,
    41576 => -47,
    41577 => -47,
    41578 => -47,
    41579 => -47,
    41580 => -47,
    41581 => -47,
    41582 => -47,
    41583 => -47,
    41584 => -47,
    41585 => -47,
    41586 => -47,
    41587 => -47,
    41588 => -47,
    41589 => -47,
    41590 => -47,
    41591 => -47,
    41592 => -47,
    41593 => -47,
    41594 => -47,
    41595 => -47,
    41596 => -47,
    41597 => -47,
    41598 => -47,
    41599 => -47,
    41600 => -47,
    41601 => -47,
    41602 => -47,
    41603 => -47,
    41604 => -47,
    41605 => -47,
    41606 => -47,
    41607 => -47,
    41608 => -47,
    41609 => -47,
    41610 => -47,
    41611 => -47,
    41612 => -47,
    41613 => -47,
    41614 => -47,
    41615 => -47,
    41616 => -47,
    41617 => -47,
    41618 => -47,
    41619 => -47,
    41620 => -47,
    41621 => -47,
    41622 => -47,
    41623 => -47,
    41624 => -47,
    41625 => -47,
    41626 => -47,
    41627 => -47,
    41628 => -47,
    41629 => -47,
    41630 => -47,
    41631 => -47,
    41632 => -47,
    41633 => -47,
    41634 => -47,
    41635 => -47,
    41636 => -47,
    41637 => -47,
    41638 => -47,
    41639 => -47,
    41640 => -47,
    41641 => -47,
    41642 => -47,
    41643 => -47,
    41644 => -47,
    41645 => -47,
    41646 => -47,
    41647 => -47,
    41648 => -47,
    41649 => -47,
    41650 => -47,
    41651 => -47,
    41652 => -47,
    41653 => -47,
    41654 => -47,
    41655 => -47,
    41656 => -47,
    41657 => -47,
    41658 => -47,
    41659 => -47,
    41660 => -47,
    41661 => -47,
    41662 => -47,
    41663 => -47,
    41664 => -47,
    41665 => -47,
    41666 => -47,
    41667 => -47,
    41668 => -47,
    41669 => -47,
    41670 => -47,
    41671 => -47,
    41672 => -47,
    41673 => -47,
    41674 => -47,
    41675 => -47,
    41676 => -47,
    41677 => -48,
    41678 => -48,
    41679 => -48,
    41680 => -48,
    41681 => -48,
    41682 => -48,
    41683 => -48,
    41684 => -48,
    41685 => -48,
    41686 => -48,
    41687 => -48,
    41688 => -48,
    41689 => -48,
    41690 => -48,
    41691 => -48,
    41692 => -48,
    41693 => -48,
    41694 => -48,
    41695 => -48,
    41696 => -48,
    41697 => -48,
    41698 => -48,
    41699 => -48,
    41700 => -48,
    41701 => -48,
    41702 => -48,
    41703 => -48,
    41704 => -48,
    41705 => -48,
    41706 => -48,
    41707 => -48,
    41708 => -48,
    41709 => -48,
    41710 => -48,
    41711 => -48,
    41712 => -48,
    41713 => -48,
    41714 => -48,
    41715 => -48,
    41716 => -48,
    41717 => -48,
    41718 => -48,
    41719 => -48,
    41720 => -48,
    41721 => -48,
    41722 => -48,
    41723 => -48,
    41724 => -48,
    41725 => -48,
    41726 => -48,
    41727 => -48,
    41728 => -48,
    41729 => -48,
    41730 => -48,
    41731 => -48,
    41732 => -48,
    41733 => -48,
    41734 => -48,
    41735 => -48,
    41736 => -48,
    41737 => -48,
    41738 => -48,
    41739 => -48,
    41740 => -48,
    41741 => -48,
    41742 => -48,
    41743 => -48,
    41744 => -48,
    41745 => -48,
    41746 => -48,
    41747 => -48,
    41748 => -48,
    41749 => -48,
    41750 => -48,
    41751 => -48,
    41752 => -48,
    41753 => -48,
    41754 => -48,
    41755 => -48,
    41756 => -48,
    41757 => -48,
    41758 => -48,
    41759 => -48,
    41760 => -48,
    41761 => -48,
    41762 => -48,
    41763 => -48,
    41764 => -48,
    41765 => -48,
    41766 => -48,
    41767 => -48,
    41768 => -48,
    41769 => -48,
    41770 => -48,
    41771 => -48,
    41772 => -48,
    41773 => -48,
    41774 => -48,
    41775 => -48,
    41776 => -48,
    41777 => -48,
    41778 => -48,
    41779 => -48,
    41780 => -48,
    41781 => -48,
    41782 => -48,
    41783 => -48,
    41784 => -48,
    41785 => -48,
    41786 => -48,
    41787 => -48,
    41788 => -48,
    41789 => -48,
    41790 => -48,
    41791 => -48,
    41792 => -48,
    41793 => -48,
    41794 => -48,
    41795 => -48,
    41796 => -48,
    41797 => -48,
    41798 => -48,
    41799 => -48,
    41800 => -48,
    41801 => -48,
    41802 => -48,
    41803 => -48,
    41804 => -48,
    41805 => -48,
    41806 => -48,
    41807 => -48,
    41808 => -48,
    41809 => -48,
    41810 => -48,
    41811 => -48,
    41812 => -48,
    41813 => -48,
    41814 => -48,
    41815 => -48,
    41816 => -48,
    41817 => -48,
    41818 => -48,
    41819 => -48,
    41820 => -48,
    41821 => -48,
    41822 => -48,
    41823 => -48,
    41824 => -48,
    41825 => -48,
    41826 => -48,
    41827 => -48,
    41828 => -48,
    41829 => -48,
    41830 => -48,
    41831 => -48,
    41832 => -48,
    41833 => -48,
    41834 => -48,
    41835 => -48,
    41836 => -48,
    41837 => -48,
    41838 => -48,
    41839 => -48,
    41840 => -48,
    41841 => -48,
    41842 => -48,
    41843 => -48,
    41844 => -48,
    41845 => -48,
    41846 => -48,
    41847 => -48,
    41848 => -48,
    41849 => -48,
    41850 => -48,
    41851 => -48,
    41852 => -48,
    41853 => -48,
    41854 => -48,
    41855 => -48,
    41856 => -48,
    41857 => -48,
    41858 => -48,
    41859 => -48,
    41860 => -48,
    41861 => -48,
    41862 => -48,
    41863 => -48,
    41864 => -48,
    41865 => -48,
    41866 => -48,
    41867 => -48,
    41868 => -48,
    41869 => -48,
    41870 => -48,
    41871 => -48,
    41872 => -48,
    41873 => -48,
    41874 => -48,
    41875 => -48,
    41876 => -48,
    41877 => -48,
    41878 => -48,
    41879 => -48,
    41880 => -48,
    41881 => -48,
    41882 => -48,
    41883 => -48,
    41884 => -48,
    41885 => -48,
    41886 => -48,
    41887 => -48,
    41888 => -48,
    41889 => -48,
    41890 => -48,
    41891 => -48,
    41892 => -48,
    41893 => -48,
    41894 => -48,
    41895 => -48,
    41896 => -48,
    41897 => -48,
    41898 => -48,
    41899 => -48,
    41900 => -48,
    41901 => -48,
    41902 => -48,
    41903 => -48,
    41904 => -48,
    41905 => -48,
    41906 => -48,
    41907 => -48,
    41908 => -48,
    41909 => -48,
    41910 => -48,
    41911 => -48,
    41912 => -48,
    41913 => -48,
    41914 => -48,
    41915 => -48,
    41916 => -48,
    41917 => -48,
    41918 => -48,
    41919 => -48,
    41920 => -48,
    41921 => -48,
    41922 => -48,
    41923 => -48,
    41924 => -48,
    41925 => -48,
    41926 => -48,
    41927 => -48,
    41928 => -48,
    41929 => -48,
    41930 => -48,
    41931 => -48,
    41932 => -48,
    41933 => -49,
    41934 => -49,
    41935 => -49,
    41936 => -49,
    41937 => -49,
    41938 => -49,
    41939 => -49,
    41940 => -49,
    41941 => -49,
    41942 => -49,
    41943 => -49,
    41944 => -49,
    41945 => -49,
    41946 => -49,
    41947 => -49,
    41948 => -49,
    41949 => -49,
    41950 => -49,
    41951 => -49,
    41952 => -49,
    41953 => -49,
    41954 => -49,
    41955 => -49,
    41956 => -49,
    41957 => -49,
    41958 => -49,
    41959 => -49,
    41960 => -49,
    41961 => -49,
    41962 => -49,
    41963 => -49,
    41964 => -49,
    41965 => -49,
    41966 => -49,
    41967 => -49,
    41968 => -49,
    41969 => -49,
    41970 => -49,
    41971 => -49,
    41972 => -49,
    41973 => -49,
    41974 => -49,
    41975 => -49,
    41976 => -49,
    41977 => -49,
    41978 => -49,
    41979 => -49,
    41980 => -49,
    41981 => -49,
    41982 => -49,
    41983 => -49,
    41984 => -49,
    41985 => -49,
    41986 => -49,
    41987 => -49,
    41988 => -49,
    41989 => -49,
    41990 => -49,
    41991 => -49,
    41992 => -49,
    41993 => -49,
    41994 => -49,
    41995 => -49,
    41996 => -49,
    41997 => -49,
    41998 => -49,
    41999 => -49,
    42000 => -49,
    42001 => -49,
    42002 => -49,
    42003 => -49,
    42004 => -49,
    42005 => -49,
    42006 => -49,
    42007 => -49,
    42008 => -49,
    42009 => -49,
    42010 => -49,
    42011 => -49,
    42012 => -49,
    42013 => -49,
    42014 => -49,
    42015 => -49,
    42016 => -49,
    42017 => -49,
    42018 => -49,
    42019 => -49,
    42020 => -49,
    42021 => -49,
    42022 => -49,
    42023 => -49,
    42024 => -49,
    42025 => -49,
    42026 => -49,
    42027 => -49,
    42028 => -49,
    42029 => -49,
    42030 => -49,
    42031 => -49,
    42032 => -49,
    42033 => -49,
    42034 => -49,
    42035 => -49,
    42036 => -49,
    42037 => -49,
    42038 => -49,
    42039 => -49,
    42040 => -49,
    42041 => -49,
    42042 => -49,
    42043 => -49,
    42044 => -49,
    42045 => -49,
    42046 => -49,
    42047 => -49,
    42048 => -49,
    42049 => -49,
    42050 => -49,
    42051 => -49,
    42052 => -49,
    42053 => -49,
    42054 => -49,
    42055 => -49,
    42056 => -49,
    42057 => -49,
    42058 => -49,
    42059 => -49,
    42060 => -49,
    42061 => -49,
    42062 => -49,
    42063 => -49,
    42064 => -49,
    42065 => -49,
    42066 => -49,
    42067 => -49,
    42068 => -49,
    42069 => -49,
    42070 => -49,
    42071 => -49,
    42072 => -49,
    42073 => -49,
    42074 => -49,
    42075 => -49,
    42076 => -49,
    42077 => -49,
    42078 => -49,
    42079 => -49,
    42080 => -49,
    42081 => -49,
    42082 => -49,
    42083 => -49,
    42084 => -49,
    42085 => -49,
    42086 => -49,
    42087 => -49,
    42088 => -49,
    42089 => -49,
    42090 => -49,
    42091 => -49,
    42092 => -49,
    42093 => -49,
    42094 => -49,
    42095 => -49,
    42096 => -49,
    42097 => -49,
    42098 => -49,
    42099 => -49,
    42100 => -49,
    42101 => -49,
    42102 => -49,
    42103 => -49,
    42104 => -49,
    42105 => -49,
    42106 => -49,
    42107 => -49,
    42108 => -49,
    42109 => -49,
    42110 => -49,
    42111 => -49,
    42112 => -49,
    42113 => -49,
    42114 => -49,
    42115 => -49,
    42116 => -49,
    42117 => -49,
    42118 => -49,
    42119 => -49,
    42120 => -49,
    42121 => -49,
    42122 => -49,
    42123 => -49,
    42124 => -49,
    42125 => -49,
    42126 => -49,
    42127 => -49,
    42128 => -49,
    42129 => -49,
    42130 => -49,
    42131 => -49,
    42132 => -49,
    42133 => -49,
    42134 => -49,
    42135 => -49,
    42136 => -49,
    42137 => -49,
    42138 => -49,
    42139 => -49,
    42140 => -49,
    42141 => -49,
    42142 => -49,
    42143 => -49,
    42144 => -49,
    42145 => -49,
    42146 => -49,
    42147 => -49,
    42148 => -49,
    42149 => -49,
    42150 => -49,
    42151 => -49,
    42152 => -49,
    42153 => -49,
    42154 => -49,
    42155 => -49,
    42156 => -49,
    42157 => -49,
    42158 => -49,
    42159 => -49,
    42160 => -49,
    42161 => -49,
    42162 => -49,
    42163 => -49,
    42164 => -49,
    42165 => -49,
    42166 => -49,
    42167 => -49,
    42168 => -49,
    42169 => -49,
    42170 => -49,
    42171 => -49,
    42172 => -49,
    42173 => -49,
    42174 => -49,
    42175 => -49,
    42176 => -49,
    42177 => -49,
    42178 => -49,
    42179 => -49,
    42180 => -49,
    42181 => -49,
    42182 => -49,
    42183 => -49,
    42184 => -49,
    42185 => -49,
    42186 => -49,
    42187 => -49,
    42188 => -49,
    42189 => -49,
    42190 => -49,
    42191 => -49,
    42192 => -49,
    42193 => -49,
    42194 => -49,
    42195 => -49,
    42196 => -50,
    42197 => -50,
    42198 => -50,
    42199 => -50,
    42200 => -50,
    42201 => -50,
    42202 => -50,
    42203 => -50,
    42204 => -50,
    42205 => -50,
    42206 => -50,
    42207 => -50,
    42208 => -50,
    42209 => -50,
    42210 => -50,
    42211 => -50,
    42212 => -50,
    42213 => -50,
    42214 => -50,
    42215 => -50,
    42216 => -50,
    42217 => -50,
    42218 => -50,
    42219 => -50,
    42220 => -50,
    42221 => -50,
    42222 => -50,
    42223 => -50,
    42224 => -50,
    42225 => -50,
    42226 => -50,
    42227 => -50,
    42228 => -50,
    42229 => -50,
    42230 => -50,
    42231 => -50,
    42232 => -50,
    42233 => -50,
    42234 => -50,
    42235 => -50,
    42236 => -50,
    42237 => -50,
    42238 => -50,
    42239 => -50,
    42240 => -50,
    42241 => -50,
    42242 => -50,
    42243 => -50,
    42244 => -50,
    42245 => -50,
    42246 => -50,
    42247 => -50,
    42248 => -50,
    42249 => -50,
    42250 => -50,
    42251 => -50,
    42252 => -50,
    42253 => -50,
    42254 => -50,
    42255 => -50,
    42256 => -50,
    42257 => -50,
    42258 => -50,
    42259 => -50,
    42260 => -50,
    42261 => -50,
    42262 => -50,
    42263 => -50,
    42264 => -50,
    42265 => -50,
    42266 => -50,
    42267 => -50,
    42268 => -50,
    42269 => -50,
    42270 => -50,
    42271 => -50,
    42272 => -50,
    42273 => -50,
    42274 => -50,
    42275 => -50,
    42276 => -50,
    42277 => -50,
    42278 => -50,
    42279 => -50,
    42280 => -50,
    42281 => -50,
    42282 => -50,
    42283 => -50,
    42284 => -50,
    42285 => -50,
    42286 => -50,
    42287 => -50,
    42288 => -50,
    42289 => -50,
    42290 => -50,
    42291 => -50,
    42292 => -50,
    42293 => -50,
    42294 => -50,
    42295 => -50,
    42296 => -50,
    42297 => -50,
    42298 => -50,
    42299 => -50,
    42300 => -50,
    42301 => -50,
    42302 => -50,
    42303 => -50,
    42304 => -50,
    42305 => -50,
    42306 => -50,
    42307 => -50,
    42308 => -50,
    42309 => -50,
    42310 => -50,
    42311 => -50,
    42312 => -50,
    42313 => -50,
    42314 => -50,
    42315 => -50,
    42316 => -50,
    42317 => -50,
    42318 => -50,
    42319 => -50,
    42320 => -50,
    42321 => -50,
    42322 => -50,
    42323 => -50,
    42324 => -50,
    42325 => -50,
    42326 => -50,
    42327 => -50,
    42328 => -50,
    42329 => -50,
    42330 => -50,
    42331 => -50,
    42332 => -50,
    42333 => -50,
    42334 => -50,
    42335 => -50,
    42336 => -50,
    42337 => -50,
    42338 => -50,
    42339 => -50,
    42340 => -50,
    42341 => -50,
    42342 => -50,
    42343 => -50,
    42344 => -50,
    42345 => -50,
    42346 => -50,
    42347 => -50,
    42348 => -50,
    42349 => -50,
    42350 => -50,
    42351 => -50,
    42352 => -50,
    42353 => -50,
    42354 => -50,
    42355 => -50,
    42356 => -50,
    42357 => -50,
    42358 => -50,
    42359 => -50,
    42360 => -50,
    42361 => -50,
    42362 => -50,
    42363 => -50,
    42364 => -50,
    42365 => -50,
    42366 => -50,
    42367 => -50,
    42368 => -50,
    42369 => -50,
    42370 => -50,
    42371 => -50,
    42372 => -50,
    42373 => -50,
    42374 => -50,
    42375 => -50,
    42376 => -50,
    42377 => -50,
    42378 => -50,
    42379 => -50,
    42380 => -50,
    42381 => -50,
    42382 => -50,
    42383 => -50,
    42384 => -50,
    42385 => -50,
    42386 => -50,
    42387 => -50,
    42388 => -50,
    42389 => -50,
    42390 => -50,
    42391 => -50,
    42392 => -50,
    42393 => -50,
    42394 => -50,
    42395 => -50,
    42396 => -50,
    42397 => -50,
    42398 => -50,
    42399 => -50,
    42400 => -50,
    42401 => -50,
    42402 => -50,
    42403 => -50,
    42404 => -50,
    42405 => -50,
    42406 => -50,
    42407 => -50,
    42408 => -50,
    42409 => -50,
    42410 => -50,
    42411 => -50,
    42412 => -50,
    42413 => -50,
    42414 => -50,
    42415 => -50,
    42416 => -50,
    42417 => -50,
    42418 => -50,
    42419 => -50,
    42420 => -50,
    42421 => -50,
    42422 => -50,
    42423 => -50,
    42424 => -50,
    42425 => -50,
    42426 => -50,
    42427 => -50,
    42428 => -50,
    42429 => -50,
    42430 => -50,
    42431 => -50,
    42432 => -50,
    42433 => -50,
    42434 => -50,
    42435 => -50,
    42436 => -50,
    42437 => -50,
    42438 => -50,
    42439 => -50,
    42440 => -50,
    42441 => -50,
    42442 => -50,
    42443 => -50,
    42444 => -50,
    42445 => -50,
    42446 => -50,
    42447 => -50,
    42448 => -50,
    42449 => -50,
    42450 => -50,
    42451 => -50,
    42452 => -50,
    42453 => -50,
    42454 => -50,
    42455 => -50,
    42456 => -50,
    42457 => -50,
    42458 => -50,
    42459 => -50,
    42460 => -50,
    42461 => -50,
    42462 => -50,
    42463 => -50,
    42464 => -50,
    42465 => -50,
    42466 => -50,
    42467 => -50,
    42468 => -51,
    42469 => -51,
    42470 => -51,
    42471 => -51,
    42472 => -51,
    42473 => -51,
    42474 => -51,
    42475 => -51,
    42476 => -51,
    42477 => -51,
    42478 => -51,
    42479 => -51,
    42480 => -51,
    42481 => -51,
    42482 => -51,
    42483 => -51,
    42484 => -51,
    42485 => -51,
    42486 => -51,
    42487 => -51,
    42488 => -51,
    42489 => -51,
    42490 => -51,
    42491 => -51,
    42492 => -51,
    42493 => -51,
    42494 => -51,
    42495 => -51,
    42496 => -51,
    42497 => -51,
    42498 => -51,
    42499 => -51,
    42500 => -51,
    42501 => -51,
    42502 => -51,
    42503 => -51,
    42504 => -51,
    42505 => -51,
    42506 => -51,
    42507 => -51,
    42508 => -51,
    42509 => -51,
    42510 => -51,
    42511 => -51,
    42512 => -51,
    42513 => -51,
    42514 => -51,
    42515 => -51,
    42516 => -51,
    42517 => -51,
    42518 => -51,
    42519 => -51,
    42520 => -51,
    42521 => -51,
    42522 => -51,
    42523 => -51,
    42524 => -51,
    42525 => -51,
    42526 => -51,
    42527 => -51,
    42528 => -51,
    42529 => -51,
    42530 => -51,
    42531 => -51,
    42532 => -51,
    42533 => -51,
    42534 => -51,
    42535 => -51,
    42536 => -51,
    42537 => -51,
    42538 => -51,
    42539 => -51,
    42540 => -51,
    42541 => -51,
    42542 => -51,
    42543 => -51,
    42544 => -51,
    42545 => -51,
    42546 => -51,
    42547 => -51,
    42548 => -51,
    42549 => -51,
    42550 => -51,
    42551 => -51,
    42552 => -51,
    42553 => -51,
    42554 => -51,
    42555 => -51,
    42556 => -51,
    42557 => -51,
    42558 => -51,
    42559 => -51,
    42560 => -51,
    42561 => -51,
    42562 => -51,
    42563 => -51,
    42564 => -51,
    42565 => -51,
    42566 => -51,
    42567 => -51,
    42568 => -51,
    42569 => -51,
    42570 => -51,
    42571 => -51,
    42572 => -51,
    42573 => -51,
    42574 => -51,
    42575 => -51,
    42576 => -51,
    42577 => -51,
    42578 => -51,
    42579 => -51,
    42580 => -51,
    42581 => -51,
    42582 => -51,
    42583 => -51,
    42584 => -51,
    42585 => -51,
    42586 => -51,
    42587 => -51,
    42588 => -51,
    42589 => -51,
    42590 => -51,
    42591 => -51,
    42592 => -51,
    42593 => -51,
    42594 => -51,
    42595 => -51,
    42596 => -51,
    42597 => -51,
    42598 => -51,
    42599 => -51,
    42600 => -51,
    42601 => -51,
    42602 => -51,
    42603 => -51,
    42604 => -51,
    42605 => -51,
    42606 => -51,
    42607 => -51,
    42608 => -51,
    42609 => -51,
    42610 => -51,
    42611 => -51,
    42612 => -51,
    42613 => -51,
    42614 => -51,
    42615 => -51,
    42616 => -51,
    42617 => -51,
    42618 => -51,
    42619 => -51,
    42620 => -51,
    42621 => -51,
    42622 => -51,
    42623 => -51,
    42624 => -51,
    42625 => -51,
    42626 => -51,
    42627 => -51,
    42628 => -51,
    42629 => -51,
    42630 => -51,
    42631 => -51,
    42632 => -51,
    42633 => -51,
    42634 => -51,
    42635 => -51,
    42636 => -51,
    42637 => -51,
    42638 => -51,
    42639 => -51,
    42640 => -51,
    42641 => -51,
    42642 => -51,
    42643 => -51,
    42644 => -51,
    42645 => -51,
    42646 => -51,
    42647 => -51,
    42648 => -51,
    42649 => -51,
    42650 => -51,
    42651 => -51,
    42652 => -51,
    42653 => -51,
    42654 => -51,
    42655 => -51,
    42656 => -51,
    42657 => -51,
    42658 => -51,
    42659 => -51,
    42660 => -51,
    42661 => -51,
    42662 => -51,
    42663 => -51,
    42664 => -51,
    42665 => -51,
    42666 => -51,
    42667 => -51,
    42668 => -51,
    42669 => -51,
    42670 => -51,
    42671 => -51,
    42672 => -51,
    42673 => -51,
    42674 => -51,
    42675 => -51,
    42676 => -51,
    42677 => -51,
    42678 => -51,
    42679 => -51,
    42680 => -51,
    42681 => -51,
    42682 => -51,
    42683 => -51,
    42684 => -51,
    42685 => -51,
    42686 => -51,
    42687 => -51,
    42688 => -51,
    42689 => -51,
    42690 => -51,
    42691 => -51,
    42692 => -51,
    42693 => -51,
    42694 => -51,
    42695 => -51,
    42696 => -51,
    42697 => -51,
    42698 => -51,
    42699 => -51,
    42700 => -51,
    42701 => -51,
    42702 => -51,
    42703 => -51,
    42704 => -51,
    42705 => -51,
    42706 => -51,
    42707 => -51,
    42708 => -51,
    42709 => -51,
    42710 => -51,
    42711 => -51,
    42712 => -51,
    42713 => -51,
    42714 => -51,
    42715 => -51,
    42716 => -51,
    42717 => -51,
    42718 => -51,
    42719 => -51,
    42720 => -51,
    42721 => -51,
    42722 => -51,
    42723 => -51,
    42724 => -51,
    42725 => -51,
    42726 => -51,
    42727 => -51,
    42728 => -51,
    42729 => -51,
    42730 => -51,
    42731 => -51,
    42732 => -51,
    42733 => -51,
    42734 => -51,
    42735 => -51,
    42736 => -51,
    42737 => -51,
    42738 => -51,
    42739 => -51,
    42740 => -51,
    42741 => -51,
    42742 => -51,
    42743 => -51,
    42744 => -51,
    42745 => -51,
    42746 => -51,
    42747 => -51,
    42748 => -51,
    42749 => -51,
    42750 => -52,
    42751 => -52,
    42752 => -52,
    42753 => -52,
    42754 => -52,
    42755 => -52,
    42756 => -52,
    42757 => -52,
    42758 => -52,
    42759 => -52,
    42760 => -52,
    42761 => -52,
    42762 => -52,
    42763 => -52,
    42764 => -52,
    42765 => -52,
    42766 => -52,
    42767 => -52,
    42768 => -52,
    42769 => -52,
    42770 => -52,
    42771 => -52,
    42772 => -52,
    42773 => -52,
    42774 => -52,
    42775 => -52,
    42776 => -52,
    42777 => -52,
    42778 => -52,
    42779 => -52,
    42780 => -52,
    42781 => -52,
    42782 => -52,
    42783 => -52,
    42784 => -52,
    42785 => -52,
    42786 => -52,
    42787 => -52,
    42788 => -52,
    42789 => -52,
    42790 => -52,
    42791 => -52,
    42792 => -52,
    42793 => -52,
    42794 => -52,
    42795 => -52,
    42796 => -52,
    42797 => -52,
    42798 => -52,
    42799 => -52,
    42800 => -52,
    42801 => -52,
    42802 => -52,
    42803 => -52,
    42804 => -52,
    42805 => -52,
    42806 => -52,
    42807 => -52,
    42808 => -52,
    42809 => -52,
    42810 => -52,
    42811 => -52,
    42812 => -52,
    42813 => -52,
    42814 => -52,
    42815 => -52,
    42816 => -52,
    42817 => -52,
    42818 => -52,
    42819 => -52,
    42820 => -52,
    42821 => -52,
    42822 => -52,
    42823 => -52,
    42824 => -52,
    42825 => -52,
    42826 => -52,
    42827 => -52,
    42828 => -52,
    42829 => -52,
    42830 => -52,
    42831 => -52,
    42832 => -52,
    42833 => -52,
    42834 => -52,
    42835 => -52,
    42836 => -52,
    42837 => -52,
    42838 => -52,
    42839 => -52,
    42840 => -52,
    42841 => -52,
    42842 => -52,
    42843 => -52,
    42844 => -52,
    42845 => -52,
    42846 => -52,
    42847 => -52,
    42848 => -52,
    42849 => -52,
    42850 => -52,
    42851 => -52,
    42852 => -52,
    42853 => -52,
    42854 => -52,
    42855 => -52,
    42856 => -52,
    42857 => -52,
    42858 => -52,
    42859 => -52,
    42860 => -52,
    42861 => -52,
    42862 => -52,
    42863 => -52,
    42864 => -52,
    42865 => -52,
    42866 => -52,
    42867 => -52,
    42868 => -52,
    42869 => -52,
    42870 => -52,
    42871 => -52,
    42872 => -52,
    42873 => -52,
    42874 => -52,
    42875 => -52,
    42876 => -52,
    42877 => -52,
    42878 => -52,
    42879 => -52,
    42880 => -52,
    42881 => -52,
    42882 => -52,
    42883 => -52,
    42884 => -52,
    42885 => -52,
    42886 => -52,
    42887 => -52,
    42888 => -52,
    42889 => -52,
    42890 => -52,
    42891 => -52,
    42892 => -52,
    42893 => -52,
    42894 => -52,
    42895 => -52,
    42896 => -52,
    42897 => -52,
    42898 => -52,
    42899 => -52,
    42900 => -52,
    42901 => -52,
    42902 => -52,
    42903 => -52,
    42904 => -52,
    42905 => -52,
    42906 => -52,
    42907 => -52,
    42908 => -52,
    42909 => -52,
    42910 => -52,
    42911 => -52,
    42912 => -52,
    42913 => -52,
    42914 => -52,
    42915 => -52,
    42916 => -52,
    42917 => -52,
    42918 => -52,
    42919 => -52,
    42920 => -52,
    42921 => -52,
    42922 => -52,
    42923 => -52,
    42924 => -52,
    42925 => -52,
    42926 => -52,
    42927 => -52,
    42928 => -52,
    42929 => -52,
    42930 => -52,
    42931 => -52,
    42932 => -52,
    42933 => -52,
    42934 => -52,
    42935 => -52,
    42936 => -52,
    42937 => -52,
    42938 => -52,
    42939 => -52,
    42940 => -52,
    42941 => -52,
    42942 => -52,
    42943 => -52,
    42944 => -52,
    42945 => -52,
    42946 => -52,
    42947 => -52,
    42948 => -52,
    42949 => -52,
    42950 => -52,
    42951 => -52,
    42952 => -52,
    42953 => -52,
    42954 => -52,
    42955 => -52,
    42956 => -52,
    42957 => -52,
    42958 => -52,
    42959 => -52,
    42960 => -52,
    42961 => -52,
    42962 => -52,
    42963 => -52,
    42964 => -52,
    42965 => -52,
    42966 => -52,
    42967 => -52,
    42968 => -52,
    42969 => -52,
    42970 => -52,
    42971 => -52,
    42972 => -52,
    42973 => -52,
    42974 => -52,
    42975 => -52,
    42976 => -52,
    42977 => -52,
    42978 => -52,
    42979 => -52,
    42980 => -52,
    42981 => -52,
    42982 => -52,
    42983 => -52,
    42984 => -52,
    42985 => -52,
    42986 => -52,
    42987 => -52,
    42988 => -52,
    42989 => -52,
    42990 => -52,
    42991 => -52,
    42992 => -52,
    42993 => -52,
    42994 => -52,
    42995 => -52,
    42996 => -52,
    42997 => -52,
    42998 => -52,
    42999 => -52,
    43000 => -52,
    43001 => -52,
    43002 => -52,
    43003 => -52,
    43004 => -52,
    43005 => -52,
    43006 => -52,
    43007 => -52,
    43008 => -52,
    43009 => -52,
    43010 => -52,
    43011 => -52,
    43012 => -52,
    43013 => -52,
    43014 => -52,
    43015 => -52,
    43016 => -52,
    43017 => -52,
    43018 => -52,
    43019 => -52,
    43020 => -52,
    43021 => -52,
    43022 => -52,
    43023 => -52,
    43024 => -52,
    43025 => -52,
    43026 => -52,
    43027 => -52,
    43028 => -52,
    43029 => -52,
    43030 => -52,
    43031 => -52,
    43032 => -52,
    43033 => -52,
    43034 => -52,
    43035 => -52,
    43036 => -52,
    43037 => -52,
    43038 => -52,
    43039 => -52,
    43040 => -52,
    43041 => -52,
    43042 => -52,
    43043 => -52,
    43044 => -53,
    43045 => -53,
    43046 => -53,
    43047 => -53,
    43048 => -53,
    43049 => -53,
    43050 => -53,
    43051 => -53,
    43052 => -53,
    43053 => -53,
    43054 => -53,
    43055 => -53,
    43056 => -53,
    43057 => -53,
    43058 => -53,
    43059 => -53,
    43060 => -53,
    43061 => -53,
    43062 => -53,
    43063 => -53,
    43064 => -53,
    43065 => -53,
    43066 => -53,
    43067 => -53,
    43068 => -53,
    43069 => -53,
    43070 => -53,
    43071 => -53,
    43072 => -53,
    43073 => -53,
    43074 => -53,
    43075 => -53,
    43076 => -53,
    43077 => -53,
    43078 => -53,
    43079 => -53,
    43080 => -53,
    43081 => -53,
    43082 => -53,
    43083 => -53,
    43084 => -53,
    43085 => -53,
    43086 => -53,
    43087 => -53,
    43088 => -53,
    43089 => -53,
    43090 => -53,
    43091 => -53,
    43092 => -53,
    43093 => -53,
    43094 => -53,
    43095 => -53,
    43096 => -53,
    43097 => -53,
    43098 => -53,
    43099 => -53,
    43100 => -53,
    43101 => -53,
    43102 => -53,
    43103 => -53,
    43104 => -53,
    43105 => -53,
    43106 => -53,
    43107 => -53,
    43108 => -53,
    43109 => -53,
    43110 => -53,
    43111 => -53,
    43112 => -53,
    43113 => -53,
    43114 => -53,
    43115 => -53,
    43116 => -53,
    43117 => -53,
    43118 => -53,
    43119 => -53,
    43120 => -53,
    43121 => -53,
    43122 => -53,
    43123 => -53,
    43124 => -53,
    43125 => -53,
    43126 => -53,
    43127 => -53,
    43128 => -53,
    43129 => -53,
    43130 => -53,
    43131 => -53,
    43132 => -53,
    43133 => -53,
    43134 => -53,
    43135 => -53,
    43136 => -53,
    43137 => -53,
    43138 => -53,
    43139 => -53,
    43140 => -53,
    43141 => -53,
    43142 => -53,
    43143 => -53,
    43144 => -53,
    43145 => -53,
    43146 => -53,
    43147 => -53,
    43148 => -53,
    43149 => -53,
    43150 => -53,
    43151 => -53,
    43152 => -53,
    43153 => -53,
    43154 => -53,
    43155 => -53,
    43156 => -53,
    43157 => -53,
    43158 => -53,
    43159 => -53,
    43160 => -53,
    43161 => -53,
    43162 => -53,
    43163 => -53,
    43164 => -53,
    43165 => -53,
    43166 => -53,
    43167 => -53,
    43168 => -53,
    43169 => -53,
    43170 => -53,
    43171 => -53,
    43172 => -53,
    43173 => -53,
    43174 => -53,
    43175 => -53,
    43176 => -53,
    43177 => -53,
    43178 => -53,
    43179 => -53,
    43180 => -53,
    43181 => -53,
    43182 => -53,
    43183 => -53,
    43184 => -53,
    43185 => -53,
    43186 => -53,
    43187 => -53,
    43188 => -53,
    43189 => -53,
    43190 => -53,
    43191 => -53,
    43192 => -53,
    43193 => -53,
    43194 => -53,
    43195 => -53,
    43196 => -53,
    43197 => -53,
    43198 => -53,
    43199 => -53,
    43200 => -53,
    43201 => -53,
    43202 => -53,
    43203 => -53,
    43204 => -53,
    43205 => -53,
    43206 => -53,
    43207 => -53,
    43208 => -53,
    43209 => -53,
    43210 => -53,
    43211 => -53,
    43212 => -53,
    43213 => -53,
    43214 => -53,
    43215 => -53,
    43216 => -53,
    43217 => -53,
    43218 => -53,
    43219 => -53,
    43220 => -53,
    43221 => -53,
    43222 => -53,
    43223 => -53,
    43224 => -53,
    43225 => -53,
    43226 => -53,
    43227 => -53,
    43228 => -53,
    43229 => -53,
    43230 => -53,
    43231 => -53,
    43232 => -53,
    43233 => -53,
    43234 => -53,
    43235 => -53,
    43236 => -53,
    43237 => -53,
    43238 => -53,
    43239 => -53,
    43240 => -53,
    43241 => -53,
    43242 => -53,
    43243 => -53,
    43244 => -53,
    43245 => -53,
    43246 => -53,
    43247 => -53,
    43248 => -53,
    43249 => -53,
    43250 => -53,
    43251 => -53,
    43252 => -53,
    43253 => -53,
    43254 => -53,
    43255 => -53,
    43256 => -53,
    43257 => -53,
    43258 => -53,
    43259 => -53,
    43260 => -53,
    43261 => -53,
    43262 => -53,
    43263 => -53,
    43264 => -53,
    43265 => -53,
    43266 => -53,
    43267 => -53,
    43268 => -53,
    43269 => -53,
    43270 => -53,
    43271 => -53,
    43272 => -53,
    43273 => -53,
    43274 => -53,
    43275 => -53,
    43276 => -53,
    43277 => -53,
    43278 => -53,
    43279 => -53,
    43280 => -53,
    43281 => -53,
    43282 => -53,
    43283 => -53,
    43284 => -53,
    43285 => -53,
    43286 => -53,
    43287 => -53,
    43288 => -53,
    43289 => -53,
    43290 => -53,
    43291 => -53,
    43292 => -53,
    43293 => -53,
    43294 => -53,
    43295 => -53,
    43296 => -53,
    43297 => -53,
    43298 => -53,
    43299 => -53,
    43300 => -53,
    43301 => -53,
    43302 => -53,
    43303 => -53,
    43304 => -53,
    43305 => -53,
    43306 => -53,
    43307 => -53,
    43308 => -53,
    43309 => -53,
    43310 => -53,
    43311 => -53,
    43312 => -53,
    43313 => -53,
    43314 => -53,
    43315 => -53,
    43316 => -53,
    43317 => -53,
    43318 => -53,
    43319 => -53,
    43320 => -53,
    43321 => -53,
    43322 => -53,
    43323 => -53,
    43324 => -53,
    43325 => -53,
    43326 => -53,
    43327 => -53,
    43328 => -53,
    43329 => -53,
    43330 => -53,
    43331 => -53,
    43332 => -53,
    43333 => -53,
    43334 => -53,
    43335 => -53,
    43336 => -53,
    43337 => -53,
    43338 => -53,
    43339 => -53,
    43340 => -53,
    43341 => -53,
    43342 => -53,
    43343 => -53,
    43344 => -53,
    43345 => -53,
    43346 => -53,
    43347 => -53,
    43348 => -53,
    43349 => -53,
    43350 => -54,
    43351 => -54,
    43352 => -54,
    43353 => -54,
    43354 => -54,
    43355 => -54,
    43356 => -54,
    43357 => -54,
    43358 => -54,
    43359 => -54,
    43360 => -54,
    43361 => -54,
    43362 => -54,
    43363 => -54,
    43364 => -54,
    43365 => -54,
    43366 => -54,
    43367 => -54,
    43368 => -54,
    43369 => -54,
    43370 => -54,
    43371 => -54,
    43372 => -54,
    43373 => -54,
    43374 => -54,
    43375 => -54,
    43376 => -54,
    43377 => -54,
    43378 => -54,
    43379 => -54,
    43380 => -54,
    43381 => -54,
    43382 => -54,
    43383 => -54,
    43384 => -54,
    43385 => -54,
    43386 => -54,
    43387 => -54,
    43388 => -54,
    43389 => -54,
    43390 => -54,
    43391 => -54,
    43392 => -54,
    43393 => -54,
    43394 => -54,
    43395 => -54,
    43396 => -54,
    43397 => -54,
    43398 => -54,
    43399 => -54,
    43400 => -54,
    43401 => -54,
    43402 => -54,
    43403 => -54,
    43404 => -54,
    43405 => -54,
    43406 => -54,
    43407 => -54,
    43408 => -54,
    43409 => -54,
    43410 => -54,
    43411 => -54,
    43412 => -54,
    43413 => -54,
    43414 => -54,
    43415 => -54,
    43416 => -54,
    43417 => -54,
    43418 => -54,
    43419 => -54,
    43420 => -54,
    43421 => -54,
    43422 => -54,
    43423 => -54,
    43424 => -54,
    43425 => -54,
    43426 => -54,
    43427 => -54,
    43428 => -54,
    43429 => -54,
    43430 => -54,
    43431 => -54,
    43432 => -54,
    43433 => -54,
    43434 => -54,
    43435 => -54,
    43436 => -54,
    43437 => -54,
    43438 => -54,
    43439 => -54,
    43440 => -54,
    43441 => -54,
    43442 => -54,
    43443 => -54,
    43444 => -54,
    43445 => -54,
    43446 => -54,
    43447 => -54,
    43448 => -54,
    43449 => -54,
    43450 => -54,
    43451 => -54,
    43452 => -54,
    43453 => -54,
    43454 => -54,
    43455 => -54,
    43456 => -54,
    43457 => -54,
    43458 => -54,
    43459 => -54,
    43460 => -54,
    43461 => -54,
    43462 => -54,
    43463 => -54,
    43464 => -54,
    43465 => -54,
    43466 => -54,
    43467 => -54,
    43468 => -54,
    43469 => -54,
    43470 => -54,
    43471 => -54,
    43472 => -54,
    43473 => -54,
    43474 => -54,
    43475 => -54,
    43476 => -54,
    43477 => -54,
    43478 => -54,
    43479 => -54,
    43480 => -54,
    43481 => -54,
    43482 => -54,
    43483 => -54,
    43484 => -54,
    43485 => -54,
    43486 => -54,
    43487 => -54,
    43488 => -54,
    43489 => -54,
    43490 => -54,
    43491 => -54,
    43492 => -54,
    43493 => -54,
    43494 => -54,
    43495 => -54,
    43496 => -54,
    43497 => -54,
    43498 => -54,
    43499 => -54,
    43500 => -54,
    43501 => -54,
    43502 => -54,
    43503 => -54,
    43504 => -54,
    43505 => -54,
    43506 => -54,
    43507 => -54,
    43508 => -54,
    43509 => -54,
    43510 => -54,
    43511 => -54,
    43512 => -54,
    43513 => -54,
    43514 => -54,
    43515 => -54,
    43516 => -54,
    43517 => -54,
    43518 => -54,
    43519 => -54,
    43520 => -54,
    43521 => -54,
    43522 => -54,
    43523 => -54,
    43524 => -54,
    43525 => -54,
    43526 => -54,
    43527 => -54,
    43528 => -54,
    43529 => -54,
    43530 => -54,
    43531 => -54,
    43532 => -54,
    43533 => -54,
    43534 => -54,
    43535 => -54,
    43536 => -54,
    43537 => -54,
    43538 => -54,
    43539 => -54,
    43540 => -54,
    43541 => -54,
    43542 => -54,
    43543 => -54,
    43544 => -54,
    43545 => -54,
    43546 => -54,
    43547 => -54,
    43548 => -54,
    43549 => -54,
    43550 => -54,
    43551 => -54,
    43552 => -54,
    43553 => -54,
    43554 => -54,
    43555 => -54,
    43556 => -54,
    43557 => -54,
    43558 => -54,
    43559 => -54,
    43560 => -54,
    43561 => -54,
    43562 => -54,
    43563 => -54,
    43564 => -54,
    43565 => -54,
    43566 => -54,
    43567 => -54,
    43568 => -54,
    43569 => -54,
    43570 => -54,
    43571 => -54,
    43572 => -54,
    43573 => -54,
    43574 => -54,
    43575 => -54,
    43576 => -54,
    43577 => -54,
    43578 => -54,
    43579 => -54,
    43580 => -54,
    43581 => -54,
    43582 => -54,
    43583 => -54,
    43584 => -54,
    43585 => -54,
    43586 => -54,
    43587 => -54,
    43588 => -54,
    43589 => -54,
    43590 => -54,
    43591 => -54,
    43592 => -54,
    43593 => -54,
    43594 => -54,
    43595 => -54,
    43596 => -54,
    43597 => -54,
    43598 => -54,
    43599 => -54,
    43600 => -54,
    43601 => -54,
    43602 => -54,
    43603 => -54,
    43604 => -54,
    43605 => -54,
    43606 => -54,
    43607 => -54,
    43608 => -54,
    43609 => -54,
    43610 => -54,
    43611 => -54,
    43612 => -54,
    43613 => -54,
    43614 => -54,
    43615 => -54,
    43616 => -54,
    43617 => -54,
    43618 => -54,
    43619 => -54,
    43620 => -54,
    43621 => -54,
    43622 => -54,
    43623 => -54,
    43624 => -54,
    43625 => -54,
    43626 => -54,
    43627 => -54,
    43628 => -54,
    43629 => -54,
    43630 => -54,
    43631 => -54,
    43632 => -54,
    43633 => -54,
    43634 => -54,
    43635 => -54,
    43636 => -54,
    43637 => -54,
    43638 => -54,
    43639 => -54,
    43640 => -54,
    43641 => -54,
    43642 => -54,
    43643 => -54,
    43644 => -54,
    43645 => -54,
    43646 => -54,
    43647 => -54,
    43648 => -54,
    43649 => -54,
    43650 => -54,
    43651 => -54,
    43652 => -54,
    43653 => -54,
    43654 => -54,
    43655 => -54,
    43656 => -54,
    43657 => -54,
    43658 => -54,
    43659 => -54,
    43660 => -54,
    43661 => -54,
    43662 => -54,
    43663 => -54,
    43664 => -54,
    43665 => -54,
    43666 => -54,
    43667 => -54,
    43668 => -54,
    43669 => -54,
    43670 => -54,
    43671 => -55,
    43672 => -55,
    43673 => -55,
    43674 => -55,
    43675 => -55,
    43676 => -55,
    43677 => -55,
    43678 => -55,
    43679 => -55,
    43680 => -55,
    43681 => -55,
    43682 => -55,
    43683 => -55,
    43684 => -55,
    43685 => -55,
    43686 => -55,
    43687 => -55,
    43688 => -55,
    43689 => -55,
    43690 => -55,
    43691 => -55,
    43692 => -55,
    43693 => -55,
    43694 => -55,
    43695 => -55,
    43696 => -55,
    43697 => -55,
    43698 => -55,
    43699 => -55,
    43700 => -55,
    43701 => -55,
    43702 => -55,
    43703 => -55,
    43704 => -55,
    43705 => -55,
    43706 => -55,
    43707 => -55,
    43708 => -55,
    43709 => -55,
    43710 => -55,
    43711 => -55,
    43712 => -55,
    43713 => -55,
    43714 => -55,
    43715 => -55,
    43716 => -55,
    43717 => -55,
    43718 => -55,
    43719 => -55,
    43720 => -55,
    43721 => -55,
    43722 => -55,
    43723 => -55,
    43724 => -55,
    43725 => -55,
    43726 => -55,
    43727 => -55,
    43728 => -55,
    43729 => -55,
    43730 => -55,
    43731 => -55,
    43732 => -55,
    43733 => -55,
    43734 => -55,
    43735 => -55,
    43736 => -55,
    43737 => -55,
    43738 => -55,
    43739 => -55,
    43740 => -55,
    43741 => -55,
    43742 => -55,
    43743 => -55,
    43744 => -55,
    43745 => -55,
    43746 => -55,
    43747 => -55,
    43748 => -55,
    43749 => -55,
    43750 => -55,
    43751 => -55,
    43752 => -55,
    43753 => -55,
    43754 => -55,
    43755 => -55,
    43756 => -55,
    43757 => -55,
    43758 => -55,
    43759 => -55,
    43760 => -55,
    43761 => -55,
    43762 => -55,
    43763 => -55,
    43764 => -55,
    43765 => -55,
    43766 => -55,
    43767 => -55,
    43768 => -55,
    43769 => -55,
    43770 => -55,
    43771 => -55,
    43772 => -55,
    43773 => -55,
    43774 => -55,
    43775 => -55,
    43776 => -55,
    43777 => -55,
    43778 => -55,
    43779 => -55,
    43780 => -55,
    43781 => -55,
    43782 => -55,
    43783 => -55,
    43784 => -55,
    43785 => -55,
    43786 => -55,
    43787 => -55,
    43788 => -55,
    43789 => -55,
    43790 => -55,
    43791 => -55,
    43792 => -55,
    43793 => -55,
    43794 => -55,
    43795 => -55,
    43796 => -55,
    43797 => -55,
    43798 => -55,
    43799 => -55,
    43800 => -55,
    43801 => -55,
    43802 => -55,
    43803 => -55,
    43804 => -55,
    43805 => -55,
    43806 => -55,
    43807 => -55,
    43808 => -55,
    43809 => -55,
    43810 => -55,
    43811 => -55,
    43812 => -55,
    43813 => -55,
    43814 => -55,
    43815 => -55,
    43816 => -55,
    43817 => -55,
    43818 => -55,
    43819 => -55,
    43820 => -55,
    43821 => -55,
    43822 => -55,
    43823 => -55,
    43824 => -55,
    43825 => -55,
    43826 => -55,
    43827 => -55,
    43828 => -55,
    43829 => -55,
    43830 => -55,
    43831 => -55,
    43832 => -55,
    43833 => -55,
    43834 => -55,
    43835 => -55,
    43836 => -55,
    43837 => -55,
    43838 => -55,
    43839 => -55,
    43840 => -55,
    43841 => -55,
    43842 => -55,
    43843 => -55,
    43844 => -55,
    43845 => -55,
    43846 => -55,
    43847 => -55,
    43848 => -55,
    43849 => -55,
    43850 => -55,
    43851 => -55,
    43852 => -55,
    43853 => -55,
    43854 => -55,
    43855 => -55,
    43856 => -55,
    43857 => -55,
    43858 => -55,
    43859 => -55,
    43860 => -55,
    43861 => -55,
    43862 => -55,
    43863 => -55,
    43864 => -55,
    43865 => -55,
    43866 => -55,
    43867 => -55,
    43868 => -55,
    43869 => -55,
    43870 => -55,
    43871 => -55,
    43872 => -55,
    43873 => -55,
    43874 => -55,
    43875 => -55,
    43876 => -55,
    43877 => -55,
    43878 => -55,
    43879 => -55,
    43880 => -55,
    43881 => -55,
    43882 => -55,
    43883 => -55,
    43884 => -55,
    43885 => -55,
    43886 => -55,
    43887 => -55,
    43888 => -55,
    43889 => -55,
    43890 => -55,
    43891 => -55,
    43892 => -55,
    43893 => -55,
    43894 => -55,
    43895 => -55,
    43896 => -55,
    43897 => -55,
    43898 => -55,
    43899 => -55,
    43900 => -55,
    43901 => -55,
    43902 => -55,
    43903 => -55,
    43904 => -55,
    43905 => -55,
    43906 => -55,
    43907 => -55,
    43908 => -55,
    43909 => -55,
    43910 => -55,
    43911 => -55,
    43912 => -55,
    43913 => -55,
    43914 => -55,
    43915 => -55,
    43916 => -55,
    43917 => -55,
    43918 => -55,
    43919 => -55,
    43920 => -55,
    43921 => -55,
    43922 => -55,
    43923 => -55,
    43924 => -55,
    43925 => -55,
    43926 => -55,
    43927 => -55,
    43928 => -55,
    43929 => -55,
    43930 => -55,
    43931 => -55,
    43932 => -55,
    43933 => -55,
    43934 => -55,
    43935 => -55,
    43936 => -55,
    43937 => -55,
    43938 => -55,
    43939 => -55,
    43940 => -55,
    43941 => -55,
    43942 => -55,
    43943 => -55,
    43944 => -55,
    43945 => -55,
    43946 => -55,
    43947 => -55,
    43948 => -55,
    43949 => -55,
    43950 => -55,
    43951 => -55,
    43952 => -55,
    43953 => -55,
    43954 => -55,
    43955 => -55,
    43956 => -55,
    43957 => -55,
    43958 => -55,
    43959 => -55,
    43960 => -55,
    43961 => -55,
    43962 => -55,
    43963 => -55,
    43964 => -55,
    43965 => -55,
    43966 => -55,
    43967 => -55,
    43968 => -55,
    43969 => -55,
    43970 => -55,
    43971 => -55,
    43972 => -55,
    43973 => -55,
    43974 => -55,
    43975 => -55,
    43976 => -55,
    43977 => -55,
    43978 => -55,
    43979 => -55,
    43980 => -55,
    43981 => -55,
    43982 => -55,
    43983 => -55,
    43984 => -55,
    43985 => -55,
    43986 => -55,
    43987 => -55,
    43988 => -55,
    43989 => -55,
    43990 => -55,
    43991 => -55,
    43992 => -55,
    43993 => -55,
    43994 => -55,
    43995 => -55,
    43996 => -55,
    43997 => -55,
    43998 => -55,
    43999 => -55,
    44000 => -55,
    44001 => -55,
    44002 => -55,
    44003 => -55,
    44004 => -55,
    44005 => -55,
    44006 => -55,
    44007 => -55,
    44008 => -55,
    44009 => -55,
    44010 => -55,
    44011 => -56,
    44012 => -56,
    44013 => -56,
    44014 => -56,
    44015 => -56,
    44016 => -56,
    44017 => -56,
    44018 => -56,
    44019 => -56,
    44020 => -56,
    44021 => -56,
    44022 => -56,
    44023 => -56,
    44024 => -56,
    44025 => -56,
    44026 => -56,
    44027 => -56,
    44028 => -56,
    44029 => -56,
    44030 => -56,
    44031 => -56,
    44032 => -56,
    44033 => -56,
    44034 => -56,
    44035 => -56,
    44036 => -56,
    44037 => -56,
    44038 => -56,
    44039 => -56,
    44040 => -56,
    44041 => -56,
    44042 => -56,
    44043 => -56,
    44044 => -56,
    44045 => -56,
    44046 => -56,
    44047 => -56,
    44048 => -56,
    44049 => -56,
    44050 => -56,
    44051 => -56,
    44052 => -56,
    44053 => -56,
    44054 => -56,
    44055 => -56,
    44056 => -56,
    44057 => -56,
    44058 => -56,
    44059 => -56,
    44060 => -56,
    44061 => -56,
    44062 => -56,
    44063 => -56,
    44064 => -56,
    44065 => -56,
    44066 => -56,
    44067 => -56,
    44068 => -56,
    44069 => -56,
    44070 => -56,
    44071 => -56,
    44072 => -56,
    44073 => -56,
    44074 => -56,
    44075 => -56,
    44076 => -56,
    44077 => -56,
    44078 => -56,
    44079 => -56,
    44080 => -56,
    44081 => -56,
    44082 => -56,
    44083 => -56,
    44084 => -56,
    44085 => -56,
    44086 => -56,
    44087 => -56,
    44088 => -56,
    44089 => -56,
    44090 => -56,
    44091 => -56,
    44092 => -56,
    44093 => -56,
    44094 => -56,
    44095 => -56,
    44096 => -56,
    44097 => -56,
    44098 => -56,
    44099 => -56,
    44100 => -56,
    44101 => -56,
    44102 => -56,
    44103 => -56,
    44104 => -56,
    44105 => -56,
    44106 => -56,
    44107 => -56,
    44108 => -56,
    44109 => -56,
    44110 => -56,
    44111 => -56,
    44112 => -56,
    44113 => -56,
    44114 => -56,
    44115 => -56,
    44116 => -56,
    44117 => -56,
    44118 => -56,
    44119 => -56,
    44120 => -56,
    44121 => -56,
    44122 => -56,
    44123 => -56,
    44124 => -56,
    44125 => -56,
    44126 => -56,
    44127 => -56,
    44128 => -56,
    44129 => -56,
    44130 => -56,
    44131 => -56,
    44132 => -56,
    44133 => -56,
    44134 => -56,
    44135 => -56,
    44136 => -56,
    44137 => -56,
    44138 => -56,
    44139 => -56,
    44140 => -56,
    44141 => -56,
    44142 => -56,
    44143 => -56,
    44144 => -56,
    44145 => -56,
    44146 => -56,
    44147 => -56,
    44148 => -56,
    44149 => -56,
    44150 => -56,
    44151 => -56,
    44152 => -56,
    44153 => -56,
    44154 => -56,
    44155 => -56,
    44156 => -56,
    44157 => -56,
    44158 => -56,
    44159 => -56,
    44160 => -56,
    44161 => -56,
    44162 => -56,
    44163 => -56,
    44164 => -56,
    44165 => -56,
    44166 => -56,
    44167 => -56,
    44168 => -56,
    44169 => -56,
    44170 => -56,
    44171 => -56,
    44172 => -56,
    44173 => -56,
    44174 => -56,
    44175 => -56,
    44176 => -56,
    44177 => -56,
    44178 => -56,
    44179 => -56,
    44180 => -56,
    44181 => -56,
    44182 => -56,
    44183 => -56,
    44184 => -56,
    44185 => -56,
    44186 => -56,
    44187 => -56,
    44188 => -56,
    44189 => -56,
    44190 => -56,
    44191 => -56,
    44192 => -56,
    44193 => -56,
    44194 => -56,
    44195 => -56,
    44196 => -56,
    44197 => -56,
    44198 => -56,
    44199 => -56,
    44200 => -56,
    44201 => -56,
    44202 => -56,
    44203 => -56,
    44204 => -56,
    44205 => -56,
    44206 => -56,
    44207 => -56,
    44208 => -56,
    44209 => -56,
    44210 => -56,
    44211 => -56,
    44212 => -56,
    44213 => -56,
    44214 => -56,
    44215 => -56,
    44216 => -56,
    44217 => -56,
    44218 => -56,
    44219 => -56,
    44220 => -56,
    44221 => -56,
    44222 => -56,
    44223 => -56,
    44224 => -56,
    44225 => -56,
    44226 => -56,
    44227 => -56,
    44228 => -56,
    44229 => -56,
    44230 => -56,
    44231 => -56,
    44232 => -56,
    44233 => -56,
    44234 => -56,
    44235 => -56,
    44236 => -56,
    44237 => -56,
    44238 => -56,
    44239 => -56,
    44240 => -56,
    44241 => -56,
    44242 => -56,
    44243 => -56,
    44244 => -56,
    44245 => -56,
    44246 => -56,
    44247 => -56,
    44248 => -56,
    44249 => -56,
    44250 => -56,
    44251 => -56,
    44252 => -56,
    44253 => -56,
    44254 => -56,
    44255 => -56,
    44256 => -56,
    44257 => -56,
    44258 => -56,
    44259 => -56,
    44260 => -56,
    44261 => -56,
    44262 => -56,
    44263 => -56,
    44264 => -56,
    44265 => -56,
    44266 => -56,
    44267 => -56,
    44268 => -56,
    44269 => -56,
    44270 => -56,
    44271 => -56,
    44272 => -56,
    44273 => -56,
    44274 => -56,
    44275 => -56,
    44276 => -56,
    44277 => -56,
    44278 => -56,
    44279 => -56,
    44280 => -56,
    44281 => -56,
    44282 => -56,
    44283 => -56,
    44284 => -56,
    44285 => -56,
    44286 => -56,
    44287 => -56,
    44288 => -56,
    44289 => -56,
    44290 => -56,
    44291 => -56,
    44292 => -56,
    44293 => -56,
    44294 => -56,
    44295 => -56,
    44296 => -56,
    44297 => -56,
    44298 => -56,
    44299 => -56,
    44300 => -56,
    44301 => -56,
    44302 => -56,
    44303 => -56,
    44304 => -56,
    44305 => -56,
    44306 => -56,
    44307 => -56,
    44308 => -56,
    44309 => -56,
    44310 => -56,
    44311 => -56,
    44312 => -56,
    44313 => -56,
    44314 => -56,
    44315 => -56,
    44316 => -56,
    44317 => -56,
    44318 => -56,
    44319 => -56,
    44320 => -56,
    44321 => -56,
    44322 => -56,
    44323 => -56,
    44324 => -56,
    44325 => -56,
    44326 => -56,
    44327 => -56,
    44328 => -56,
    44329 => -56,
    44330 => -56,
    44331 => -56,
    44332 => -56,
    44333 => -56,
    44334 => -56,
    44335 => -56,
    44336 => -56,
    44337 => -56,
    44338 => -56,
    44339 => -56,
    44340 => -56,
    44341 => -56,
    44342 => -56,
    44343 => -56,
    44344 => -56,
    44345 => -56,
    44346 => -56,
    44347 => -56,
    44348 => -56,
    44349 => -56,
    44350 => -56,
    44351 => -56,
    44352 => -56,
    44353 => -56,
    44354 => -56,
    44355 => -56,
    44356 => -56,
    44357 => -56,
    44358 => -56,
    44359 => -56,
    44360 => -56,
    44361 => -56,
    44362 => -56,
    44363 => -56,
    44364 => -56,
    44365 => -56,
    44366 => -56,
    44367 => -56,
    44368 => -56,
    44369 => -56,
    44370 => -56,
    44371 => -56,
    44372 => -56,
    44373 => -57,
    44374 => -57,
    44375 => -57,
    44376 => -57,
    44377 => -57,
    44378 => -57,
    44379 => -57,
    44380 => -57,
    44381 => -57,
    44382 => -57,
    44383 => -57,
    44384 => -57,
    44385 => -57,
    44386 => -57,
    44387 => -57,
    44388 => -57,
    44389 => -57,
    44390 => -57,
    44391 => -57,
    44392 => -57,
    44393 => -57,
    44394 => -57,
    44395 => -57,
    44396 => -57,
    44397 => -57,
    44398 => -57,
    44399 => -57,
    44400 => -57,
    44401 => -57,
    44402 => -57,
    44403 => -57,
    44404 => -57,
    44405 => -57,
    44406 => -57,
    44407 => -57,
    44408 => -57,
    44409 => -57,
    44410 => -57,
    44411 => -57,
    44412 => -57,
    44413 => -57,
    44414 => -57,
    44415 => -57,
    44416 => -57,
    44417 => -57,
    44418 => -57,
    44419 => -57,
    44420 => -57,
    44421 => -57,
    44422 => -57,
    44423 => -57,
    44424 => -57,
    44425 => -57,
    44426 => -57,
    44427 => -57,
    44428 => -57,
    44429 => -57,
    44430 => -57,
    44431 => -57,
    44432 => -57,
    44433 => -57,
    44434 => -57,
    44435 => -57,
    44436 => -57,
    44437 => -57,
    44438 => -57,
    44439 => -57,
    44440 => -57,
    44441 => -57,
    44442 => -57,
    44443 => -57,
    44444 => -57,
    44445 => -57,
    44446 => -57,
    44447 => -57,
    44448 => -57,
    44449 => -57,
    44450 => -57,
    44451 => -57,
    44452 => -57,
    44453 => -57,
    44454 => -57,
    44455 => -57,
    44456 => -57,
    44457 => -57,
    44458 => -57,
    44459 => -57,
    44460 => -57,
    44461 => -57,
    44462 => -57,
    44463 => -57,
    44464 => -57,
    44465 => -57,
    44466 => -57,
    44467 => -57,
    44468 => -57,
    44469 => -57,
    44470 => -57,
    44471 => -57,
    44472 => -57,
    44473 => -57,
    44474 => -57,
    44475 => -57,
    44476 => -57,
    44477 => -57,
    44478 => -57,
    44479 => -57,
    44480 => -57,
    44481 => -57,
    44482 => -57,
    44483 => -57,
    44484 => -57,
    44485 => -57,
    44486 => -57,
    44487 => -57,
    44488 => -57,
    44489 => -57,
    44490 => -57,
    44491 => -57,
    44492 => -57,
    44493 => -57,
    44494 => -57,
    44495 => -57,
    44496 => -57,
    44497 => -57,
    44498 => -57,
    44499 => -57,
    44500 => -57,
    44501 => -57,
    44502 => -57,
    44503 => -57,
    44504 => -57,
    44505 => -57,
    44506 => -57,
    44507 => -57,
    44508 => -57,
    44509 => -57,
    44510 => -57,
    44511 => -57,
    44512 => -57,
    44513 => -57,
    44514 => -57,
    44515 => -57,
    44516 => -57,
    44517 => -57,
    44518 => -57,
    44519 => -57,
    44520 => -57,
    44521 => -57,
    44522 => -57,
    44523 => -57,
    44524 => -57,
    44525 => -57,
    44526 => -57,
    44527 => -57,
    44528 => -57,
    44529 => -57,
    44530 => -57,
    44531 => -57,
    44532 => -57,
    44533 => -57,
    44534 => -57,
    44535 => -57,
    44536 => -57,
    44537 => -57,
    44538 => -57,
    44539 => -57,
    44540 => -57,
    44541 => -57,
    44542 => -57,
    44543 => -57,
    44544 => -57,
    44545 => -57,
    44546 => -57,
    44547 => -57,
    44548 => -57,
    44549 => -57,
    44550 => -57,
    44551 => -57,
    44552 => -57,
    44553 => -57,
    44554 => -57,
    44555 => -57,
    44556 => -57,
    44557 => -57,
    44558 => -57,
    44559 => -57,
    44560 => -57,
    44561 => -57,
    44562 => -57,
    44563 => -57,
    44564 => -57,
    44565 => -57,
    44566 => -57,
    44567 => -57,
    44568 => -57,
    44569 => -57,
    44570 => -57,
    44571 => -57,
    44572 => -57,
    44573 => -57,
    44574 => -57,
    44575 => -57,
    44576 => -57,
    44577 => -57,
    44578 => -57,
    44579 => -57,
    44580 => -57,
    44581 => -57,
    44582 => -57,
    44583 => -57,
    44584 => -57,
    44585 => -57,
    44586 => -57,
    44587 => -57,
    44588 => -57,
    44589 => -57,
    44590 => -57,
    44591 => -57,
    44592 => -57,
    44593 => -57,
    44594 => -57,
    44595 => -57,
    44596 => -57,
    44597 => -57,
    44598 => -57,
    44599 => -57,
    44600 => -57,
    44601 => -57,
    44602 => -57,
    44603 => -57,
    44604 => -57,
    44605 => -57,
    44606 => -57,
    44607 => -57,
    44608 => -57,
    44609 => -57,
    44610 => -57,
    44611 => -57,
    44612 => -57,
    44613 => -57,
    44614 => -57,
    44615 => -57,
    44616 => -57,
    44617 => -57,
    44618 => -57,
    44619 => -57,
    44620 => -57,
    44621 => -57,
    44622 => -57,
    44623 => -57,
    44624 => -57,
    44625 => -57,
    44626 => -57,
    44627 => -57,
    44628 => -57,
    44629 => -57,
    44630 => -57,
    44631 => -57,
    44632 => -57,
    44633 => -57,
    44634 => -57,
    44635 => -57,
    44636 => -57,
    44637 => -57,
    44638 => -57,
    44639 => -57,
    44640 => -57,
    44641 => -57,
    44642 => -57,
    44643 => -57,
    44644 => -57,
    44645 => -57,
    44646 => -57,
    44647 => -57,
    44648 => -57,
    44649 => -57,
    44650 => -57,
    44651 => -57,
    44652 => -57,
    44653 => -57,
    44654 => -57,
    44655 => -57,
    44656 => -57,
    44657 => -57,
    44658 => -57,
    44659 => -57,
    44660 => -57,
    44661 => -57,
    44662 => -57,
    44663 => -57,
    44664 => -57,
    44665 => -57,
    44666 => -57,
    44667 => -57,
    44668 => -57,
    44669 => -57,
    44670 => -57,
    44671 => -57,
    44672 => -57,
    44673 => -57,
    44674 => -57,
    44675 => -57,
    44676 => -57,
    44677 => -57,
    44678 => -57,
    44679 => -57,
    44680 => -57,
    44681 => -57,
    44682 => -57,
    44683 => -57,
    44684 => -57,
    44685 => -57,
    44686 => -57,
    44687 => -57,
    44688 => -57,
    44689 => -57,
    44690 => -57,
    44691 => -57,
    44692 => -57,
    44693 => -57,
    44694 => -57,
    44695 => -57,
    44696 => -57,
    44697 => -57,
    44698 => -57,
    44699 => -57,
    44700 => -57,
    44701 => -57,
    44702 => -57,
    44703 => -57,
    44704 => -57,
    44705 => -57,
    44706 => -57,
    44707 => -57,
    44708 => -57,
    44709 => -57,
    44710 => -57,
    44711 => -57,
    44712 => -57,
    44713 => -57,
    44714 => -57,
    44715 => -57,
    44716 => -57,
    44717 => -57,
    44718 => -57,
    44719 => -57,
    44720 => -57,
    44721 => -57,
    44722 => -57,
    44723 => -57,
    44724 => -57,
    44725 => -57,
    44726 => -57,
    44727 => -57,
    44728 => -57,
    44729 => -57,
    44730 => -57,
    44731 => -57,
    44732 => -57,
    44733 => -57,
    44734 => -57,
    44735 => -57,
    44736 => -57,
    44737 => -57,
    44738 => -57,
    44739 => -57,
    44740 => -57,
    44741 => -57,
    44742 => -57,
    44743 => -57,
    44744 => -57,
    44745 => -57,
    44746 => -57,
    44747 => -57,
    44748 => -57,
    44749 => -57,
    44750 => -57,
    44751 => -57,
    44752 => -57,
    44753 => -57,
    44754 => -57,
    44755 => -57,
    44756 => -57,
    44757 => -57,
    44758 => -57,
    44759 => -57,
    44760 => -57,
    44761 => -57,
    44762 => -58,
    44763 => -58,
    44764 => -58,
    44765 => -58,
    44766 => -58,
    44767 => -58,
    44768 => -58,
    44769 => -58,
    44770 => -58,
    44771 => -58,
    44772 => -58,
    44773 => -58,
    44774 => -58,
    44775 => -58,
    44776 => -58,
    44777 => -58,
    44778 => -58,
    44779 => -58,
    44780 => -58,
    44781 => -58,
    44782 => -58,
    44783 => -58,
    44784 => -58,
    44785 => -58,
    44786 => -58,
    44787 => -58,
    44788 => -58,
    44789 => -58,
    44790 => -58,
    44791 => -58,
    44792 => -58,
    44793 => -58,
    44794 => -58,
    44795 => -58,
    44796 => -58,
    44797 => -58,
    44798 => -58,
    44799 => -58,
    44800 => -58,
    44801 => -58,
    44802 => -58,
    44803 => -58,
    44804 => -58,
    44805 => -58,
    44806 => -58,
    44807 => -58,
    44808 => -58,
    44809 => -58,
    44810 => -58,
    44811 => -58,
    44812 => -58,
    44813 => -58,
    44814 => -58,
    44815 => -58,
    44816 => -58,
    44817 => -58,
    44818 => -58,
    44819 => -58,
    44820 => -58,
    44821 => -58,
    44822 => -58,
    44823 => -58,
    44824 => -58,
    44825 => -58,
    44826 => -58,
    44827 => -58,
    44828 => -58,
    44829 => -58,
    44830 => -58,
    44831 => -58,
    44832 => -58,
    44833 => -58,
    44834 => -58,
    44835 => -58,
    44836 => -58,
    44837 => -58,
    44838 => -58,
    44839 => -58,
    44840 => -58,
    44841 => -58,
    44842 => -58,
    44843 => -58,
    44844 => -58,
    44845 => -58,
    44846 => -58,
    44847 => -58,
    44848 => -58,
    44849 => -58,
    44850 => -58,
    44851 => -58,
    44852 => -58,
    44853 => -58,
    44854 => -58,
    44855 => -58,
    44856 => -58,
    44857 => -58,
    44858 => -58,
    44859 => -58,
    44860 => -58,
    44861 => -58,
    44862 => -58,
    44863 => -58,
    44864 => -58,
    44865 => -58,
    44866 => -58,
    44867 => -58,
    44868 => -58,
    44869 => -58,
    44870 => -58,
    44871 => -58,
    44872 => -58,
    44873 => -58,
    44874 => -58,
    44875 => -58,
    44876 => -58,
    44877 => -58,
    44878 => -58,
    44879 => -58,
    44880 => -58,
    44881 => -58,
    44882 => -58,
    44883 => -58,
    44884 => -58,
    44885 => -58,
    44886 => -58,
    44887 => -58,
    44888 => -58,
    44889 => -58,
    44890 => -58,
    44891 => -58,
    44892 => -58,
    44893 => -58,
    44894 => -58,
    44895 => -58,
    44896 => -58,
    44897 => -58,
    44898 => -58,
    44899 => -58,
    44900 => -58,
    44901 => -58,
    44902 => -58,
    44903 => -58,
    44904 => -58,
    44905 => -58,
    44906 => -58,
    44907 => -58,
    44908 => -58,
    44909 => -58,
    44910 => -58,
    44911 => -58,
    44912 => -58,
    44913 => -58,
    44914 => -58,
    44915 => -58,
    44916 => -58,
    44917 => -58,
    44918 => -58,
    44919 => -58,
    44920 => -58,
    44921 => -58,
    44922 => -58,
    44923 => -58,
    44924 => -58,
    44925 => -58,
    44926 => -58,
    44927 => -58,
    44928 => -58,
    44929 => -58,
    44930 => -58,
    44931 => -58,
    44932 => -58,
    44933 => -58,
    44934 => -58,
    44935 => -58,
    44936 => -58,
    44937 => -58,
    44938 => -58,
    44939 => -58,
    44940 => -58,
    44941 => -58,
    44942 => -58,
    44943 => -58,
    44944 => -58,
    44945 => -58,
    44946 => -58,
    44947 => -58,
    44948 => -58,
    44949 => -58,
    44950 => -58,
    44951 => -58,
    44952 => -58,
    44953 => -58,
    44954 => -58,
    44955 => -58,
    44956 => -58,
    44957 => -58,
    44958 => -58,
    44959 => -58,
    44960 => -58,
    44961 => -58,
    44962 => -58,
    44963 => -58,
    44964 => -58,
    44965 => -58,
    44966 => -58,
    44967 => -58,
    44968 => -58,
    44969 => -58,
    44970 => -58,
    44971 => -58,
    44972 => -58,
    44973 => -58,
    44974 => -58,
    44975 => -58,
    44976 => -58,
    44977 => -58,
    44978 => -58,
    44979 => -58,
    44980 => -58,
    44981 => -58,
    44982 => -58,
    44983 => -58,
    44984 => -58,
    44985 => -58,
    44986 => -58,
    44987 => -58,
    44988 => -58,
    44989 => -58,
    44990 => -58,
    44991 => -58,
    44992 => -58,
    44993 => -58,
    44994 => -58,
    44995 => -58,
    44996 => -58,
    44997 => -58,
    44998 => -58,
    44999 => -58,
    45000 => -58,
    45001 => -58,
    45002 => -58,
    45003 => -58,
    45004 => -58,
    45005 => -58,
    45006 => -58,
    45007 => -58,
    45008 => -58,
    45009 => -58,
    45010 => -58,
    45011 => -58,
    45012 => -58,
    45013 => -58,
    45014 => -58,
    45015 => -58,
    45016 => -58,
    45017 => -58,
    45018 => -58,
    45019 => -58,
    45020 => -58,
    45021 => -58,
    45022 => -58,
    45023 => -58,
    45024 => -58,
    45025 => -58,
    45026 => -58,
    45027 => -58,
    45028 => -58,
    45029 => -58,
    45030 => -58,
    45031 => -58,
    45032 => -58,
    45033 => -58,
    45034 => -58,
    45035 => -58,
    45036 => -58,
    45037 => -58,
    45038 => -58,
    45039 => -58,
    45040 => -58,
    45041 => -58,
    45042 => -58,
    45043 => -58,
    45044 => -58,
    45045 => -58,
    45046 => -58,
    45047 => -58,
    45048 => -58,
    45049 => -58,
    45050 => -58,
    45051 => -58,
    45052 => -58,
    45053 => -58,
    45054 => -58,
    45055 => -58,
    45056 => -58,
    45057 => -58,
    45058 => -58,
    45059 => -58,
    45060 => -58,
    45061 => -58,
    45062 => -58,
    45063 => -58,
    45064 => -58,
    45065 => -58,
    45066 => -58,
    45067 => -58,
    45068 => -58,
    45069 => -58,
    45070 => -58,
    45071 => -58,
    45072 => -58,
    45073 => -58,
    45074 => -58,
    45075 => -58,
    45076 => -58,
    45077 => -58,
    45078 => -58,
    45079 => -58,
    45080 => -58,
    45081 => -58,
    45082 => -58,
    45083 => -58,
    45084 => -58,
    45085 => -58,
    45086 => -58,
    45087 => -58,
    45088 => -58,
    45089 => -58,
    45090 => -58,
    45091 => -58,
    45092 => -58,
    45093 => -58,
    45094 => -58,
    45095 => -58,
    45096 => -58,
    45097 => -58,
    45098 => -58,
    45099 => -58,
    45100 => -58,
    45101 => -58,
    45102 => -58,
    45103 => -58,
    45104 => -58,
    45105 => -58,
    45106 => -58,
    45107 => -58,
    45108 => -58,
    45109 => -58,
    45110 => -58,
    45111 => -58,
    45112 => -58,
    45113 => -58,
    45114 => -58,
    45115 => -58,
    45116 => -58,
    45117 => -58,
    45118 => -58,
    45119 => -58,
    45120 => -58,
    45121 => -58,
    45122 => -58,
    45123 => -58,
    45124 => -58,
    45125 => -58,
    45126 => -58,
    45127 => -58,
    45128 => -58,
    45129 => -58,
    45130 => -58,
    45131 => -58,
    45132 => -58,
    45133 => -58,
    45134 => -58,
    45135 => -58,
    45136 => -58,
    45137 => -58,
    45138 => -58,
    45139 => -58,
    45140 => -58,
    45141 => -58,
    45142 => -58,
    45143 => -58,
    45144 => -58,
    45145 => -58,
    45146 => -58,
    45147 => -58,
    45148 => -58,
    45149 => -58,
    45150 => -58,
    45151 => -58,
    45152 => -58,
    45153 => -58,
    45154 => -58,
    45155 => -58,
    45156 => -58,
    45157 => -58,
    45158 => -58,
    45159 => -58,
    45160 => -58,
    45161 => -58,
    45162 => -58,
    45163 => -58,
    45164 => -58,
    45165 => -58,
    45166 => -58,
    45167 => -58,
    45168 => -58,
    45169 => -58,
    45170 => -58,
    45171 => -58,
    45172 => -58,
    45173 => -58,
    45174 => -58,
    45175 => -58,
    45176 => -58,
    45177 => -58,
    45178 => -58,
    45179 => -58,
    45180 => -58,
    45181 => -58,
    45182 => -58,
    45183 => -58,
    45184 => -58,
    45185 => -58,
    45186 => -59,
    45187 => -59,
    45188 => -59,
    45189 => -59,
    45190 => -59,
    45191 => -59,
    45192 => -59,
    45193 => -59,
    45194 => -59,
    45195 => -59,
    45196 => -59,
    45197 => -59,
    45198 => -59,
    45199 => -59,
    45200 => -59,
    45201 => -59,
    45202 => -59,
    45203 => -59,
    45204 => -59,
    45205 => -59,
    45206 => -59,
    45207 => -59,
    45208 => -59,
    45209 => -59,
    45210 => -59,
    45211 => -59,
    45212 => -59,
    45213 => -59,
    45214 => -59,
    45215 => -59,
    45216 => -59,
    45217 => -59,
    45218 => -59,
    45219 => -59,
    45220 => -59,
    45221 => -59,
    45222 => -59,
    45223 => -59,
    45224 => -59,
    45225 => -59,
    45226 => -59,
    45227 => -59,
    45228 => -59,
    45229 => -59,
    45230 => -59,
    45231 => -59,
    45232 => -59,
    45233 => -59,
    45234 => -59,
    45235 => -59,
    45236 => -59,
    45237 => -59,
    45238 => -59,
    45239 => -59,
    45240 => -59,
    45241 => -59,
    45242 => -59,
    45243 => -59,
    45244 => -59,
    45245 => -59,
    45246 => -59,
    45247 => -59,
    45248 => -59,
    45249 => -59,
    45250 => -59,
    45251 => -59,
    45252 => -59,
    45253 => -59,
    45254 => -59,
    45255 => -59,
    45256 => -59,
    45257 => -59,
    45258 => -59,
    45259 => -59,
    45260 => -59,
    45261 => -59,
    45262 => -59,
    45263 => -59,
    45264 => -59,
    45265 => -59,
    45266 => -59,
    45267 => -59,
    45268 => -59,
    45269 => -59,
    45270 => -59,
    45271 => -59,
    45272 => -59,
    45273 => -59,
    45274 => -59,
    45275 => -59,
    45276 => -59,
    45277 => -59,
    45278 => -59,
    45279 => -59,
    45280 => -59,
    45281 => -59,
    45282 => -59,
    45283 => -59,
    45284 => -59,
    45285 => -59,
    45286 => -59,
    45287 => -59,
    45288 => -59,
    45289 => -59,
    45290 => -59,
    45291 => -59,
    45292 => -59,
    45293 => -59,
    45294 => -59,
    45295 => -59,
    45296 => -59,
    45297 => -59,
    45298 => -59,
    45299 => -59,
    45300 => -59,
    45301 => -59,
    45302 => -59,
    45303 => -59,
    45304 => -59,
    45305 => -59,
    45306 => -59,
    45307 => -59,
    45308 => -59,
    45309 => -59,
    45310 => -59,
    45311 => -59,
    45312 => -59,
    45313 => -59,
    45314 => -59,
    45315 => -59,
    45316 => -59,
    45317 => -59,
    45318 => -59,
    45319 => -59,
    45320 => -59,
    45321 => -59,
    45322 => -59,
    45323 => -59,
    45324 => -59,
    45325 => -59,
    45326 => -59,
    45327 => -59,
    45328 => -59,
    45329 => -59,
    45330 => -59,
    45331 => -59,
    45332 => -59,
    45333 => -59,
    45334 => -59,
    45335 => -59,
    45336 => -59,
    45337 => -59,
    45338 => -59,
    45339 => -59,
    45340 => -59,
    45341 => -59,
    45342 => -59,
    45343 => -59,
    45344 => -59,
    45345 => -59,
    45346 => -59,
    45347 => -59,
    45348 => -59,
    45349 => -59,
    45350 => -59,
    45351 => -59,
    45352 => -59,
    45353 => -59,
    45354 => -59,
    45355 => -59,
    45356 => -59,
    45357 => -59,
    45358 => -59,
    45359 => -59,
    45360 => -59,
    45361 => -59,
    45362 => -59,
    45363 => -59,
    45364 => -59,
    45365 => -59,
    45366 => -59,
    45367 => -59,
    45368 => -59,
    45369 => -59,
    45370 => -59,
    45371 => -59,
    45372 => -59,
    45373 => -59,
    45374 => -59,
    45375 => -59,
    45376 => -59,
    45377 => -59,
    45378 => -59,
    45379 => -59,
    45380 => -59,
    45381 => -59,
    45382 => -59,
    45383 => -59,
    45384 => -59,
    45385 => -59,
    45386 => -59,
    45387 => -59,
    45388 => -59,
    45389 => -59,
    45390 => -59,
    45391 => -59,
    45392 => -59,
    45393 => -59,
    45394 => -59,
    45395 => -59,
    45396 => -59,
    45397 => -59,
    45398 => -59,
    45399 => -59,
    45400 => -59,
    45401 => -59,
    45402 => -59,
    45403 => -59,
    45404 => -59,
    45405 => -59,
    45406 => -59,
    45407 => -59,
    45408 => -59,
    45409 => -59,
    45410 => -59,
    45411 => -59,
    45412 => -59,
    45413 => -59,
    45414 => -59,
    45415 => -59,
    45416 => -59,
    45417 => -59,
    45418 => -59,
    45419 => -59,
    45420 => -59,
    45421 => -59,
    45422 => -59,
    45423 => -59,
    45424 => -59,
    45425 => -59,
    45426 => -59,
    45427 => -59,
    45428 => -59,
    45429 => -59,
    45430 => -59,
    45431 => -59,
    45432 => -59,
    45433 => -59,
    45434 => -59,
    45435 => -59,
    45436 => -59,
    45437 => -59,
    45438 => -59,
    45439 => -59,
    45440 => -59,
    45441 => -59,
    45442 => -59,
    45443 => -59,
    45444 => -59,
    45445 => -59,
    45446 => -59,
    45447 => -59,
    45448 => -59,
    45449 => -59,
    45450 => -59,
    45451 => -59,
    45452 => -59,
    45453 => -59,
    45454 => -59,
    45455 => -59,
    45456 => -59,
    45457 => -59,
    45458 => -59,
    45459 => -59,
    45460 => -59,
    45461 => -59,
    45462 => -59,
    45463 => -59,
    45464 => -59,
    45465 => -59,
    45466 => -59,
    45467 => -59,
    45468 => -59,
    45469 => -59,
    45470 => -59,
    45471 => -59,
    45472 => -59,
    45473 => -59,
    45474 => -59,
    45475 => -59,
    45476 => -59,
    45477 => -59,
    45478 => -59,
    45479 => -59,
    45480 => -59,
    45481 => -59,
    45482 => -59,
    45483 => -59,
    45484 => -59,
    45485 => -59,
    45486 => -59,
    45487 => -59,
    45488 => -59,
    45489 => -59,
    45490 => -59,
    45491 => -59,
    45492 => -59,
    45493 => -59,
    45494 => -59,
    45495 => -59,
    45496 => -59,
    45497 => -59,
    45498 => -59,
    45499 => -59,
    45500 => -59,
    45501 => -59,
    45502 => -59,
    45503 => -59,
    45504 => -59,
    45505 => -59,
    45506 => -59,
    45507 => -59,
    45508 => -59,
    45509 => -59,
    45510 => -59,
    45511 => -59,
    45512 => -59,
    45513 => -59,
    45514 => -59,
    45515 => -59,
    45516 => -59,
    45517 => -59,
    45518 => -59,
    45519 => -59,
    45520 => -59,
    45521 => -59,
    45522 => -59,
    45523 => -59,
    45524 => -59,
    45525 => -59,
    45526 => -59,
    45527 => -59,
    45528 => -59,
    45529 => -59,
    45530 => -59,
    45531 => -59,
    45532 => -59,
    45533 => -59,
    45534 => -59,
    45535 => -59,
    45536 => -59,
    45537 => -59,
    45538 => -59,
    45539 => -59,
    45540 => -59,
    45541 => -59,
    45542 => -59,
    45543 => -59,
    45544 => -59,
    45545 => -59,
    45546 => -59,
    45547 => -59,
    45548 => -59,
    45549 => -59,
    45550 => -59,
    45551 => -59,
    45552 => -59,
    45553 => -59,
    45554 => -59,
    45555 => -59,
    45556 => -59,
    45557 => -59,
    45558 => -59,
    45559 => -59,
    45560 => -59,
    45561 => -59,
    45562 => -59,
    45563 => -59,
    45564 => -59,
    45565 => -59,
    45566 => -59,
    45567 => -59,
    45568 => -59,
    45569 => -59,
    45570 => -59,
    45571 => -59,
    45572 => -59,
    45573 => -59,
    45574 => -59,
    45575 => -59,
    45576 => -59,
    45577 => -59,
    45578 => -59,
    45579 => -59,
    45580 => -59,
    45581 => -59,
    45582 => -59,
    45583 => -59,
    45584 => -59,
    45585 => -59,
    45586 => -59,
    45587 => -59,
    45588 => -59,
    45589 => -59,
    45590 => -59,
    45591 => -59,
    45592 => -59,
    45593 => -59,
    45594 => -59,
    45595 => -59,
    45596 => -59,
    45597 => -59,
    45598 => -59,
    45599 => -59,
    45600 => -59,
    45601 => -59,
    45602 => -59,
    45603 => -59,
    45604 => -59,
    45605 => -59,
    45606 => -59,
    45607 => -59,
    45608 => -59,
    45609 => -59,
    45610 => -59,
    45611 => -59,
    45612 => -59,
    45613 => -59,
    45614 => -59,
    45615 => -59,
    45616 => -59,
    45617 => -59,
    45618 => -59,
    45619 => -59,
    45620 => -59,
    45621 => -59,
    45622 => -59,
    45623 => -59,
    45624 => -59,
    45625 => -59,
    45626 => -59,
    45627 => -59,
    45628 => -59,
    45629 => -59,
    45630 => -59,
    45631 => -59,
    45632 => -59,
    45633 => -59,
    45634 => -59,
    45635 => -59,
    45636 => -59,
    45637 => -59,
    45638 => -59,
    45639 => -59,
    45640 => -59,
    45641 => -59,
    45642 => -59,
    45643 => -59,
    45644 => -59,
    45645 => -59,
    45646 => -59,
    45647 => -59,
    45648 => -59,
    45649 => -59,
    45650 => -59,
    45651 => -59,
    45652 => -59,
    45653 => -59,
    45654 => -59,
    45655 => -59,
    45656 => -59,
    45657 => -59,
    45658 => -59,
    45659 => -60,
    45660 => -60,
    45661 => -60,
    45662 => -60,
    45663 => -60,
    45664 => -60,
    45665 => -60,
    45666 => -60,
    45667 => -60,
    45668 => -60,
    45669 => -60,
    45670 => -60,
    45671 => -60,
    45672 => -60,
    45673 => -60,
    45674 => -60,
    45675 => -60,
    45676 => -60,
    45677 => -60,
    45678 => -60,
    45679 => -60,
    45680 => -60,
    45681 => -60,
    45682 => -60,
    45683 => -60,
    45684 => -60,
    45685 => -60,
    45686 => -60,
    45687 => -60,
    45688 => -60,
    45689 => -60,
    45690 => -60,
    45691 => -60,
    45692 => -60,
    45693 => -60,
    45694 => -60,
    45695 => -60,
    45696 => -60,
    45697 => -60,
    45698 => -60,
    45699 => -60,
    45700 => -60,
    45701 => -60,
    45702 => -60,
    45703 => -60,
    45704 => -60,
    45705 => -60,
    45706 => -60,
    45707 => -60,
    45708 => -60,
    45709 => -60,
    45710 => -60,
    45711 => -60,
    45712 => -60,
    45713 => -60,
    45714 => -60,
    45715 => -60,
    45716 => -60,
    45717 => -60,
    45718 => -60,
    45719 => -60,
    45720 => -60,
    45721 => -60,
    45722 => -60,
    45723 => -60,
    45724 => -60,
    45725 => -60,
    45726 => -60,
    45727 => -60,
    45728 => -60,
    45729 => -60,
    45730 => -60,
    45731 => -60,
    45732 => -60,
    45733 => -60,
    45734 => -60,
    45735 => -60,
    45736 => -60,
    45737 => -60,
    45738 => -60,
    45739 => -60,
    45740 => -60,
    45741 => -60,
    45742 => -60,
    45743 => -60,
    45744 => -60,
    45745 => -60,
    45746 => -60,
    45747 => -60,
    45748 => -60,
    45749 => -60,
    45750 => -60,
    45751 => -60,
    45752 => -60,
    45753 => -60,
    45754 => -60,
    45755 => -60,
    45756 => -60,
    45757 => -60,
    45758 => -60,
    45759 => -60,
    45760 => -60,
    45761 => -60,
    45762 => -60,
    45763 => -60,
    45764 => -60,
    45765 => -60,
    45766 => -60,
    45767 => -60,
    45768 => -60,
    45769 => -60,
    45770 => -60,
    45771 => -60,
    45772 => -60,
    45773 => -60,
    45774 => -60,
    45775 => -60,
    45776 => -60,
    45777 => -60,
    45778 => -60,
    45779 => -60,
    45780 => -60,
    45781 => -60,
    45782 => -60,
    45783 => -60,
    45784 => -60,
    45785 => -60,
    45786 => -60,
    45787 => -60,
    45788 => -60,
    45789 => -60,
    45790 => -60,
    45791 => -60,
    45792 => -60,
    45793 => -60,
    45794 => -60,
    45795 => -60,
    45796 => -60,
    45797 => -60,
    45798 => -60,
    45799 => -60,
    45800 => -60,
    45801 => -60,
    45802 => -60,
    45803 => -60,
    45804 => -60,
    45805 => -60,
    45806 => -60,
    45807 => -60,
    45808 => -60,
    45809 => -60,
    45810 => -60,
    45811 => -60,
    45812 => -60,
    45813 => -60,
    45814 => -60,
    45815 => -60,
    45816 => -60,
    45817 => -60,
    45818 => -60,
    45819 => -60,
    45820 => -60,
    45821 => -60,
    45822 => -60,
    45823 => -60,
    45824 => -60,
    45825 => -60,
    45826 => -60,
    45827 => -60,
    45828 => -60,
    45829 => -60,
    45830 => -60,
    45831 => -60,
    45832 => -60,
    45833 => -60,
    45834 => -60,
    45835 => -60,
    45836 => -60,
    45837 => -60,
    45838 => -60,
    45839 => -60,
    45840 => -60,
    45841 => -60,
    45842 => -60,
    45843 => -60,
    45844 => -60,
    45845 => -60,
    45846 => -60,
    45847 => -60,
    45848 => -60,
    45849 => -60,
    45850 => -60,
    45851 => -60,
    45852 => -60,
    45853 => -60,
    45854 => -60,
    45855 => -60,
    45856 => -60,
    45857 => -60,
    45858 => -60,
    45859 => -60,
    45860 => -60,
    45861 => -60,
    45862 => -60,
    45863 => -60,
    45864 => -60,
    45865 => -60,
    45866 => -60,
    45867 => -60,
    45868 => -60,
    45869 => -60,
    45870 => -60,
    45871 => -60,
    45872 => -60,
    45873 => -60,
    45874 => -60,
    45875 => -60,
    45876 => -60,
    45877 => -60,
    45878 => -60,
    45879 => -60,
    45880 => -60,
    45881 => -60,
    45882 => -60,
    45883 => -60,
    45884 => -60,
    45885 => -60,
    45886 => -60,
    45887 => -60,
    45888 => -60,
    45889 => -60,
    45890 => -60,
    45891 => -60,
    45892 => -60,
    45893 => -60,
    45894 => -60,
    45895 => -60,
    45896 => -60,
    45897 => -60,
    45898 => -60,
    45899 => -60,
    45900 => -60,
    45901 => -60,
    45902 => -60,
    45903 => -60,
    45904 => -60,
    45905 => -60,
    45906 => -60,
    45907 => -60,
    45908 => -60,
    45909 => -60,
    45910 => -60,
    45911 => -60,
    45912 => -60,
    45913 => -60,
    45914 => -60,
    45915 => -60,
    45916 => -60,
    45917 => -60,
    45918 => -60,
    45919 => -60,
    45920 => -60,
    45921 => -60,
    45922 => -60,
    45923 => -60,
    45924 => -60,
    45925 => -60,
    45926 => -60,
    45927 => -60,
    45928 => -60,
    45929 => -60,
    45930 => -60,
    45931 => -60,
    45932 => -60,
    45933 => -60,
    45934 => -60,
    45935 => -60,
    45936 => -60,
    45937 => -60,
    45938 => -60,
    45939 => -60,
    45940 => -60,
    45941 => -60,
    45942 => -60,
    45943 => -60,
    45944 => -60,
    45945 => -60,
    45946 => -60,
    45947 => -60,
    45948 => -60,
    45949 => -60,
    45950 => -60,
    45951 => -60,
    45952 => -60,
    45953 => -60,
    45954 => -60,
    45955 => -60,
    45956 => -60,
    45957 => -60,
    45958 => -60,
    45959 => -60,
    45960 => -60,
    45961 => -60,
    45962 => -60,
    45963 => -60,
    45964 => -60,
    45965 => -60,
    45966 => -60,
    45967 => -60,
    45968 => -60,
    45969 => -60,
    45970 => -60,
    45971 => -60,
    45972 => -60,
    45973 => -60,
    45974 => -60,
    45975 => -60,
    45976 => -60,
    45977 => -60,
    45978 => -60,
    45979 => -60,
    45980 => -60,
    45981 => -60,
    45982 => -60,
    45983 => -60,
    45984 => -60,
    45985 => -60,
    45986 => -60,
    45987 => -60,
    45988 => -60,
    45989 => -60,
    45990 => -60,
    45991 => -60,
    45992 => -60,
    45993 => -60,
    45994 => -60,
    45995 => -60,
    45996 => -60,
    45997 => -60,
    45998 => -60,
    45999 => -60,
    46000 => -60,
    46001 => -60,
    46002 => -60,
    46003 => -60,
    46004 => -60,
    46005 => -60,
    46006 => -60,
    46007 => -60,
    46008 => -60,
    46009 => -60,
    46010 => -60,
    46011 => -60,
    46012 => -60,
    46013 => -60,
    46014 => -60,
    46015 => -60,
    46016 => -60,
    46017 => -60,
    46018 => -60,
    46019 => -60,
    46020 => -60,
    46021 => -60,
    46022 => -60,
    46023 => -60,
    46024 => -60,
    46025 => -60,
    46026 => -60,
    46027 => -60,
    46028 => -60,
    46029 => -60,
    46030 => -60,
    46031 => -60,
    46032 => -60,
    46033 => -60,
    46034 => -60,
    46035 => -60,
    46036 => -60,
    46037 => -60,
    46038 => -60,
    46039 => -60,
    46040 => -60,
    46041 => -60,
    46042 => -60,
    46043 => -60,
    46044 => -60,
    46045 => -60,
    46046 => -60,
    46047 => -60,
    46048 => -60,
    46049 => -60,
    46050 => -60,
    46051 => -60,
    46052 => -60,
    46053 => -60,
    46054 => -60,
    46055 => -60,
    46056 => -60,
    46057 => -60,
    46058 => -60,
    46059 => -60,
    46060 => -60,
    46061 => -60,
    46062 => -60,
    46063 => -60,
    46064 => -60,
    46065 => -60,
    46066 => -60,
    46067 => -60,
    46068 => -60,
    46069 => -60,
    46070 => -60,
    46071 => -60,
    46072 => -60,
    46073 => -60,
    46074 => -60,
    46075 => -60,
    46076 => -60,
    46077 => -60,
    46078 => -60,
    46079 => -60,
    46080 => -60,
    46081 => -60,
    46082 => -60,
    46083 => -60,
    46084 => -60,
    46085 => -60,
    46086 => -60,
    46087 => -60,
    46088 => -60,
    46089 => -60,
    46090 => -60,
    46091 => -60,
    46092 => -60,
    46093 => -60,
    46094 => -60,
    46095 => -60,
    46096 => -60,
    46097 => -60,
    46098 => -60,
    46099 => -60,
    46100 => -60,
    46101 => -60,
    46102 => -60,
    46103 => -60,
    46104 => -60,
    46105 => -60,
    46106 => -60,
    46107 => -60,
    46108 => -60,
    46109 => -60,
    46110 => -60,
    46111 => -60,
    46112 => -60,
    46113 => -60,
    46114 => -60,
    46115 => -60,
    46116 => -60,
    46117 => -60,
    46118 => -60,
    46119 => -60,
    46120 => -60,
    46121 => -60,
    46122 => -60,
    46123 => -60,
    46124 => -60,
    46125 => -60,
    46126 => -60,
    46127 => -60,
    46128 => -60,
    46129 => -60,
    46130 => -60,
    46131 => -60,
    46132 => -60,
    46133 => -60,
    46134 => -60,
    46135 => -60,
    46136 => -60,
    46137 => -60,
    46138 => -60,
    46139 => -60,
    46140 => -60,
    46141 => -60,
    46142 => -60,
    46143 => -60,
    46144 => -60,
    46145 => -60,
    46146 => -60,
    46147 => -60,
    46148 => -60,
    46149 => -60,
    46150 => -60,
    46151 => -60,
    46152 => -60,
    46153 => -60,
    46154 => -60,
    46155 => -60,
    46156 => -60,
    46157 => -60,
    46158 => -60,
    46159 => -60,
    46160 => -60,
    46161 => -60,
    46162 => -60,
    46163 => -60,
    46164 => -60,
    46165 => -60,
    46166 => -60,
    46167 => -60,
    46168 => -60,
    46169 => -60,
    46170 => -60,
    46171 => -60,
    46172 => -60,
    46173 => -60,
    46174 => -60,
    46175 => -60,
    46176 => -60,
    46177 => -60,
    46178 => -60,
    46179 => -60,
    46180 => -60,
    46181 => -60,
    46182 => -60,
    46183 => -60,
    46184 => -60,
    46185 => -60,
    46186 => -60,
    46187 => -60,
    46188 => -60,
    46189 => -60,
    46190 => -60,
    46191 => -60,
    46192 => -60,
    46193 => -60,
    46194 => -60,
    46195 => -60,
    46196 => -60,
    46197 => -60,
    46198 => -60,
    46199 => -60,
    46200 => -60,
    46201 => -60,
    46202 => -60,
    46203 => -60,
    46204 => -61,
    46205 => -61,
    46206 => -61,
    46207 => -61,
    46208 => -61,
    46209 => -61,
    46210 => -61,
    46211 => -61,
    46212 => -61,
    46213 => -61,
    46214 => -61,
    46215 => -61,
    46216 => -61,
    46217 => -61,
    46218 => -61,
    46219 => -61,
    46220 => -61,
    46221 => -61,
    46222 => -61,
    46223 => -61,
    46224 => -61,
    46225 => -61,
    46226 => -61,
    46227 => -61,
    46228 => -61,
    46229 => -61,
    46230 => -61,
    46231 => -61,
    46232 => -61,
    46233 => -61,
    46234 => -61,
    46235 => -61,
    46236 => -61,
    46237 => -61,
    46238 => -61,
    46239 => -61,
    46240 => -61,
    46241 => -61,
    46242 => -61,
    46243 => -61,
    46244 => -61,
    46245 => -61,
    46246 => -61,
    46247 => -61,
    46248 => -61,
    46249 => -61,
    46250 => -61,
    46251 => -61,
    46252 => -61,
    46253 => -61,
    46254 => -61,
    46255 => -61,
    46256 => -61,
    46257 => -61,
    46258 => -61,
    46259 => -61,
    46260 => -61,
    46261 => -61,
    46262 => -61,
    46263 => -61,
    46264 => -61,
    46265 => -61,
    46266 => -61,
    46267 => -61,
    46268 => -61,
    46269 => -61,
    46270 => -61,
    46271 => -61,
    46272 => -61,
    46273 => -61,
    46274 => -61,
    46275 => -61,
    46276 => -61,
    46277 => -61,
    46278 => -61,
    46279 => -61,
    46280 => -61,
    46281 => -61,
    46282 => -61,
    46283 => -61,
    46284 => -61,
    46285 => -61,
    46286 => -61,
    46287 => -61,
    46288 => -61,
    46289 => -61,
    46290 => -61,
    46291 => -61,
    46292 => -61,
    46293 => -61,
    46294 => -61,
    46295 => -61,
    46296 => -61,
    46297 => -61,
    46298 => -61,
    46299 => -61,
    46300 => -61,
    46301 => -61,
    46302 => -61,
    46303 => -61,
    46304 => -61,
    46305 => -61,
    46306 => -61,
    46307 => -61,
    46308 => -61,
    46309 => -61,
    46310 => -61,
    46311 => -61,
    46312 => -61,
    46313 => -61,
    46314 => -61,
    46315 => -61,
    46316 => -61,
    46317 => -61,
    46318 => -61,
    46319 => -61,
    46320 => -61,
    46321 => -61,
    46322 => -61,
    46323 => -61,
    46324 => -61,
    46325 => -61,
    46326 => -61,
    46327 => -61,
    46328 => -61,
    46329 => -61,
    46330 => -61,
    46331 => -61,
    46332 => -61,
    46333 => -61,
    46334 => -61,
    46335 => -61,
    46336 => -61,
    46337 => -61,
    46338 => -61,
    46339 => -61,
    46340 => -61,
    46341 => -61,
    46342 => -61,
    46343 => -61,
    46344 => -61,
    46345 => -61,
    46346 => -61,
    46347 => -61,
    46348 => -61,
    46349 => -61,
    46350 => -61,
    46351 => -61,
    46352 => -61,
    46353 => -61,
    46354 => -61,
    46355 => -61,
    46356 => -61,
    46357 => -61,
    46358 => -61,
    46359 => -61,
    46360 => -61,
    46361 => -61,
    46362 => -61,
    46363 => -61,
    46364 => -61,
    46365 => -61,
    46366 => -61,
    46367 => -61,
    46368 => -61,
    46369 => -61,
    46370 => -61,
    46371 => -61,
    46372 => -61,
    46373 => -61,
    46374 => -61,
    46375 => -61,
    46376 => -61,
    46377 => -61,
    46378 => -61,
    46379 => -61,
    46380 => -61,
    46381 => -61,
    46382 => -61,
    46383 => -61,
    46384 => -61,
    46385 => -61,
    46386 => -61,
    46387 => -61,
    46388 => -61,
    46389 => -61,
    46390 => -61,
    46391 => -61,
    46392 => -61,
    46393 => -61,
    46394 => -61,
    46395 => -61,
    46396 => -61,
    46397 => -61,
    46398 => -61,
    46399 => -61,
    46400 => -61,
    46401 => -61,
    46402 => -61,
    46403 => -61,
    46404 => -61,
    46405 => -61,
    46406 => -61,
    46407 => -61,
    46408 => -61,
    46409 => -61,
    46410 => -61,
    46411 => -61,
    46412 => -61,
    46413 => -61,
    46414 => -61,
    46415 => -61,
    46416 => -61,
    46417 => -61,
    46418 => -61,
    46419 => -61,
    46420 => -61,
    46421 => -61,
    46422 => -61,
    46423 => -61,
    46424 => -61,
    46425 => -61,
    46426 => -61,
    46427 => -61,
    46428 => -61,
    46429 => -61,
    46430 => -61,
    46431 => -61,
    46432 => -61,
    46433 => -61,
    46434 => -61,
    46435 => -61,
    46436 => -61,
    46437 => -61,
    46438 => -61,
    46439 => -61,
    46440 => -61,
    46441 => -61,
    46442 => -61,
    46443 => -61,
    46444 => -61,
    46445 => -61,
    46446 => -61,
    46447 => -61,
    46448 => -61,
    46449 => -61,
    46450 => -61,
    46451 => -61,
    46452 => -61,
    46453 => -61,
    46454 => -61,
    46455 => -61,
    46456 => -61,
    46457 => -61,
    46458 => -61,
    46459 => -61,
    46460 => -61,
    46461 => -61,
    46462 => -61,
    46463 => -61,
    46464 => -61,
    46465 => -61,
    46466 => -61,
    46467 => -61,
    46468 => -61,
    46469 => -61,
    46470 => -61,
    46471 => -61,
    46472 => -61,
    46473 => -61,
    46474 => -61,
    46475 => -61,
    46476 => -61,
    46477 => -61,
    46478 => -61,
    46479 => -61,
    46480 => -61,
    46481 => -61,
    46482 => -61,
    46483 => -61,
    46484 => -61,
    46485 => -61,
    46486 => -61,
    46487 => -61,
    46488 => -61,
    46489 => -61,
    46490 => -61,
    46491 => -61,
    46492 => -61,
    46493 => -61,
    46494 => -61,
    46495 => -61,
    46496 => -61,
    46497 => -61,
    46498 => -61,
    46499 => -61,
    46500 => -61,
    46501 => -61,
    46502 => -61,
    46503 => -61,
    46504 => -61,
    46505 => -61,
    46506 => -61,
    46507 => -61,
    46508 => -61,
    46509 => -61,
    46510 => -61,
    46511 => -61,
    46512 => -61,
    46513 => -61,
    46514 => -61,
    46515 => -61,
    46516 => -61,
    46517 => -61,
    46518 => -61,
    46519 => -61,
    46520 => -61,
    46521 => -61,
    46522 => -61,
    46523 => -61,
    46524 => -61,
    46525 => -61,
    46526 => -61,
    46527 => -61,
    46528 => -61,
    46529 => -61,
    46530 => -61,
    46531 => -61,
    46532 => -61,
    46533 => -61,
    46534 => -61,
    46535 => -61,
    46536 => -61,
    46537 => -61,
    46538 => -61,
    46539 => -61,
    46540 => -61,
    46541 => -61,
    46542 => -61,
    46543 => -61,
    46544 => -61,
    46545 => -61,
    46546 => -61,
    46547 => -61,
    46548 => -61,
    46549 => -61,
    46550 => -61,
    46551 => -61,
    46552 => -61,
    46553 => -61,
    46554 => -61,
    46555 => -61,
    46556 => -61,
    46557 => -61,
    46558 => -61,
    46559 => -61,
    46560 => -61,
    46561 => -61,
    46562 => -61,
    46563 => -61,
    46564 => -61,
    46565 => -61,
    46566 => -61,
    46567 => -61,
    46568 => -61,
    46569 => -61,
    46570 => -61,
    46571 => -61,
    46572 => -61,
    46573 => -61,
    46574 => -61,
    46575 => -61,
    46576 => -61,
    46577 => -61,
    46578 => -61,
    46579 => -61,
    46580 => -61,
    46581 => -61,
    46582 => -61,
    46583 => -61,
    46584 => -61,
    46585 => -61,
    46586 => -61,
    46587 => -61,
    46588 => -61,
    46589 => -61,
    46590 => -61,
    46591 => -61,
    46592 => -61,
    46593 => -61,
    46594 => -61,
    46595 => -61,
    46596 => -61,
    46597 => -61,
    46598 => -61,
    46599 => -61,
    46600 => -61,
    46601 => -61,
    46602 => -61,
    46603 => -61,
    46604 => -61,
    46605 => -61,
    46606 => -61,
    46607 => -61,
    46608 => -61,
    46609 => -61,
    46610 => -61,
    46611 => -61,
    46612 => -61,
    46613 => -61,
    46614 => -61,
    46615 => -61,
    46616 => -61,
    46617 => -61,
    46618 => -61,
    46619 => -61,
    46620 => -61,
    46621 => -61,
    46622 => -61,
    46623 => -61,
    46624 => -61,
    46625 => -61,
    46626 => -61,
    46627 => -61,
    46628 => -61,
    46629 => -61,
    46630 => -61,
    46631 => -61,
    46632 => -61,
    46633 => -61,
    46634 => -61,
    46635 => -61,
    46636 => -61,
    46637 => -61,
    46638 => -61,
    46639 => -61,
    46640 => -61,
    46641 => -61,
    46642 => -61,
    46643 => -61,
    46644 => -61,
    46645 => -61,
    46646 => -61,
    46647 => -61,
    46648 => -61,
    46649 => -61,
    46650 => -61,
    46651 => -61,
    46652 => -61,
    46653 => -61,
    46654 => -61,
    46655 => -61,
    46656 => -61,
    46657 => -61,
    46658 => -61,
    46659 => -61,
    46660 => -61,
    46661 => -61,
    46662 => -61,
    46663 => -61,
    46664 => -61,
    46665 => -61,
    46666 => -61,
    46667 => -61,
    46668 => -61,
    46669 => -61,
    46670 => -61,
    46671 => -61,
    46672 => -61,
    46673 => -61,
    46674 => -61,
    46675 => -61,
    46676 => -61,
    46677 => -61,
    46678 => -61,
    46679 => -61,
    46680 => -61,
    46681 => -61,
    46682 => -61,
    46683 => -61,
    46684 => -61,
    46685 => -61,
    46686 => -61,
    46687 => -61,
    46688 => -61,
    46689 => -61,
    46690 => -61,
    46691 => -61,
    46692 => -61,
    46693 => -61,
    46694 => -61,
    46695 => -61,
    46696 => -61,
    46697 => -61,
    46698 => -61,
    46699 => -61,
    46700 => -61,
    46701 => -61,
    46702 => -61,
    46703 => -61,
    46704 => -61,
    46705 => -61,
    46706 => -61,
    46707 => -61,
    46708 => -61,
    46709 => -61,
    46710 => -61,
    46711 => -61,
    46712 => -61,
    46713 => -61,
    46714 => -61,
    46715 => -61,
    46716 => -61,
    46717 => -61,
    46718 => -61,
    46719 => -61,
    46720 => -61,
    46721 => -61,
    46722 => -61,
    46723 => -61,
    46724 => -61,
    46725 => -61,
    46726 => -61,
    46727 => -61,
    46728 => -61,
    46729 => -61,
    46730 => -61,
    46731 => -61,
    46732 => -61,
    46733 => -61,
    46734 => -61,
    46735 => -61,
    46736 => -61,
    46737 => -61,
    46738 => -61,
    46739 => -61,
    46740 => -61,
    46741 => -61,
    46742 => -61,
    46743 => -61,
    46744 => -61,
    46745 => -61,
    46746 => -61,
    46747 => -61,
    46748 => -61,
    46749 => -61,
    46750 => -61,
    46751 => -61,
    46752 => -61,
    46753 => -61,
    46754 => -61,
    46755 => -61,
    46756 => -61,
    46757 => -61,
    46758 => -61,
    46759 => -61,
    46760 => -61,
    46761 => -61,
    46762 => -61,
    46763 => -61,
    46764 => -61,
    46765 => -61,
    46766 => -61,
    46767 => -61,
    46768 => -61,
    46769 => -61,
    46770 => -61,
    46771 => -61,
    46772 => -61,
    46773 => -61,
    46774 => -61,
    46775 => -61,
    46776 => -61,
    46777 => -61,
    46778 => -61,
    46779 => -61,
    46780 => -61,
    46781 => -61,
    46782 => -61,
    46783 => -61,
    46784 => -61,
    46785 => -61,
    46786 => -61,
    46787 => -61,
    46788 => -61,
    46789 => -61,
    46790 => -61,
    46791 => -61,
    46792 => -61,
    46793 => -61,
    46794 => -61,
    46795 => -61,
    46796 => -61,
    46797 => -61,
    46798 => -61,
    46799 => -61,
    46800 => -61,
    46801 => -61,
    46802 => -61,
    46803 => -61,
    46804 => -61,
    46805 => -61,
    46806 => -61,
    46807 => -61,
    46808 => -61,
    46809 => -61,
    46810 => -61,
    46811 => -61,
    46812 => -61,
    46813 => -61,
    46814 => -61,
    46815 => -61,
    46816 => -61,
    46817 => -61,
    46818 => -61,
    46819 => -61,
    46820 => -61,
    46821 => -61,
    46822 => -61,
    46823 => -61,
    46824 => -61,
    46825 => -61,
    46826 => -61,
    46827 => -61,
    46828 => -61,
    46829 => -61,
    46830 => -61,
    46831 => -61,
    46832 => -61,
    46833 => -61,
    46834 => -61,
    46835 => -61,
    46836 => -61,
    46837 => -61,
    46838 => -61,
    46839 => -61,
    46840 => -61,
    46841 => -61,
    46842 => -61,
    46843 => -61,
    46844 => -61,
    46845 => -61,
    46846 => -61,
    46847 => -61,
    46848 => -61,
    46849 => -61,
    46850 => -61,
    46851 => -61,
    46852 => -61,
    46853 => -61,
    46854 => -61,
    46855 => -61,
    46856 => -61,
    46857 => -61,
    46858 => -61,
    46859 => -61,
    46860 => -61,
    46861 => -61,
    46862 => -61,
    46863 => -61,
    46864 => -61,
    46865 => -61,
    46866 => -61,
    46867 => -61,
    46868 => -61,
    46869 => -61,
    46870 => -61,
    46871 => -61,
    46872 => -62,
    46873 => -62,
    46874 => -62,
    46875 => -62,
    46876 => -62,
    46877 => -62,
    46878 => -62,
    46879 => -62,
    46880 => -62,
    46881 => -62,
    46882 => -62,
    46883 => -62,
    46884 => -62,
    46885 => -62,
    46886 => -62,
    46887 => -62,
    46888 => -62,
    46889 => -62,
    46890 => -62,
    46891 => -62,
    46892 => -62,
    46893 => -62,
    46894 => -62,
    46895 => -62,
    46896 => -62,
    46897 => -62,
    46898 => -62,
    46899 => -62,
    46900 => -62,
    46901 => -62,
    46902 => -62,
    46903 => -62,
    46904 => -62,
    46905 => -62,
    46906 => -62,
    46907 => -62,
    46908 => -62,
    46909 => -62,
    46910 => -62,
    46911 => -62,
    46912 => -62,
    46913 => -62,
    46914 => -62,
    46915 => -62,
    46916 => -62,
    46917 => -62,
    46918 => -62,
    46919 => -62,
    46920 => -62,
    46921 => -62,
    46922 => -62,
    46923 => -62,
    46924 => -62,
    46925 => -62,
    46926 => -62,
    46927 => -62,
    46928 => -62,
    46929 => -62,
    46930 => -62,
    46931 => -62,
    46932 => -62,
    46933 => -62,
    46934 => -62,
    46935 => -62,
    46936 => -62,
    46937 => -62,
    46938 => -62,
    46939 => -62,
    46940 => -62,
    46941 => -62,
    46942 => -62,
    46943 => -62,
    46944 => -62,
    46945 => -62,
    46946 => -62,
    46947 => -62,
    46948 => -62,
    46949 => -62,
    46950 => -62,
    46951 => -62,
    46952 => -62,
    46953 => -62,
    46954 => -62,
    46955 => -62,
    46956 => -62,
    46957 => -62,
    46958 => -62,
    46959 => -62,
    46960 => -62,
    46961 => -62,
    46962 => -62,
    46963 => -62,
    46964 => -62,
    46965 => -62,
    46966 => -62,
    46967 => -62,
    46968 => -62,
    46969 => -62,
    46970 => -62,
    46971 => -62,
    46972 => -62,
    46973 => -62,
    46974 => -62,
    46975 => -62,
    46976 => -62,
    46977 => -62,
    46978 => -62,
    46979 => -62,
    46980 => -62,
    46981 => -62,
    46982 => -62,
    46983 => -62,
    46984 => -62,
    46985 => -62,
    46986 => -62,
    46987 => -62,
    46988 => -62,
    46989 => -62,
    46990 => -62,
    46991 => -62,
    46992 => -62,
    46993 => -62,
    46994 => -62,
    46995 => -62,
    46996 => -62,
    46997 => -62,
    46998 => -62,
    46999 => -62,
    47000 => -62,
    47001 => -62,
    47002 => -62,
    47003 => -62,
    47004 => -62,
    47005 => -62,
    47006 => -62,
    47007 => -62,
    47008 => -62,
    47009 => -62,
    47010 => -62,
    47011 => -62,
    47012 => -62,
    47013 => -62,
    47014 => -62,
    47015 => -62,
    47016 => -62,
    47017 => -62,
    47018 => -62,
    47019 => -62,
    47020 => -62,
    47021 => -62,
    47022 => -62,
    47023 => -62,
    47024 => -62,
    47025 => -62,
    47026 => -62,
    47027 => -62,
    47028 => -62,
    47029 => -62,
    47030 => -62,
    47031 => -62,
    47032 => -62,
    47033 => -62,
    47034 => -62,
    47035 => -62,
    47036 => -62,
    47037 => -62,
    47038 => -62,
    47039 => -62,
    47040 => -62,
    47041 => -62,
    47042 => -62,
    47043 => -62,
    47044 => -62,
    47045 => -62,
    47046 => -62,
    47047 => -62,
    47048 => -62,
    47049 => -62,
    47050 => -62,
    47051 => -62,
    47052 => -62,
    47053 => -62,
    47054 => -62,
    47055 => -62,
    47056 => -62,
    47057 => -62,
    47058 => -62,
    47059 => -62,
    47060 => -62,
    47061 => -62,
    47062 => -62,
    47063 => -62,
    47064 => -62,
    47065 => -62,
    47066 => -62,
    47067 => -62,
    47068 => -62,
    47069 => -62,
    47070 => -62,
    47071 => -62,
    47072 => -62,
    47073 => -62,
    47074 => -62,
    47075 => -62,
    47076 => -62,
    47077 => -62,
    47078 => -62,
    47079 => -62,
    47080 => -62,
    47081 => -62,
    47082 => -62,
    47083 => -62,
    47084 => -62,
    47085 => -62,
    47086 => -62,
    47087 => -62,
    47088 => -62,
    47089 => -62,
    47090 => -62,
    47091 => -62,
    47092 => -62,
    47093 => -62,
    47094 => -62,
    47095 => -62,
    47096 => -62,
    47097 => -62,
    47098 => -62,
    47099 => -62,
    47100 => -62,
    47101 => -62,
    47102 => -62,
    47103 => -62,
    47104 => -62,
    47105 => -62,
    47106 => -62,
    47107 => -62,
    47108 => -62,
    47109 => -62,
    47110 => -62,
    47111 => -62,
    47112 => -62,
    47113 => -62,
    47114 => -62,
    47115 => -62,
    47116 => -62,
    47117 => -62,
    47118 => -62,
    47119 => -62,
    47120 => -62,
    47121 => -62,
    47122 => -62,
    47123 => -62,
    47124 => -62,
    47125 => -62,
    47126 => -62,
    47127 => -62,
    47128 => -62,
    47129 => -62,
    47130 => -62,
    47131 => -62,
    47132 => -62,
    47133 => -62,
    47134 => -62,
    47135 => -62,
    47136 => -62,
    47137 => -62,
    47138 => -62,
    47139 => -62,
    47140 => -62,
    47141 => -62,
    47142 => -62,
    47143 => -62,
    47144 => -62,
    47145 => -62,
    47146 => -62,
    47147 => -62,
    47148 => -62,
    47149 => -62,
    47150 => -62,
    47151 => -62,
    47152 => -62,
    47153 => -62,
    47154 => -62,
    47155 => -62,
    47156 => -62,
    47157 => -62,
    47158 => -62,
    47159 => -62,
    47160 => -62,
    47161 => -62,
    47162 => -62,
    47163 => -62,
    47164 => -62,
    47165 => -62,
    47166 => -62,
    47167 => -62,
    47168 => -62,
    47169 => -62,
    47170 => -62,
    47171 => -62,
    47172 => -62,
    47173 => -62,
    47174 => -62,
    47175 => -62,
    47176 => -62,
    47177 => -62,
    47178 => -62,
    47179 => -62,
    47180 => -62,
    47181 => -62,
    47182 => -62,
    47183 => -62,
    47184 => -62,
    47185 => -62,
    47186 => -62,
    47187 => -62,
    47188 => -62,
    47189 => -62,
    47190 => -62,
    47191 => -62,
    47192 => -62,
    47193 => -62,
    47194 => -62,
    47195 => -62,
    47196 => -62,
    47197 => -62,
    47198 => -62,
    47199 => -62,
    47200 => -62,
    47201 => -62,
    47202 => -62,
    47203 => -62,
    47204 => -62,
    47205 => -62,
    47206 => -62,
    47207 => -62,
    47208 => -62,
    47209 => -62,
    47210 => -62,
    47211 => -62,
    47212 => -62,
    47213 => -62,
    47214 => -62,
    47215 => -62,
    47216 => -62,
    47217 => -62,
    47218 => -62,
    47219 => -62,
    47220 => -62,
    47221 => -62,
    47222 => -62,
    47223 => -62,
    47224 => -62,
    47225 => -62,
    47226 => -62,
    47227 => -62,
    47228 => -62,
    47229 => -62,
    47230 => -62,
    47231 => -62,
    47232 => -62,
    47233 => -62,
    47234 => -62,
    47235 => -62,
    47236 => -62,
    47237 => -62,
    47238 => -62,
    47239 => -62,
    47240 => -62,
    47241 => -62,
    47242 => -62,
    47243 => -62,
    47244 => -62,
    47245 => -62,
    47246 => -62,
    47247 => -62,
    47248 => -62,
    47249 => -62,
    47250 => -62,
    47251 => -62,
    47252 => -62,
    47253 => -62,
    47254 => -62,
    47255 => -62,
    47256 => -62,
    47257 => -62,
    47258 => -62,
    47259 => -62,
    47260 => -62,
    47261 => -62,
    47262 => -62,
    47263 => -62,
    47264 => -62,
    47265 => -62,
    47266 => -62,
    47267 => -62,
    47268 => -62,
    47269 => -62,
    47270 => -62,
    47271 => -62,
    47272 => -62,
    47273 => -62,
    47274 => -62,
    47275 => -62,
    47276 => -62,
    47277 => -62,
    47278 => -62,
    47279 => -62,
    47280 => -62,
    47281 => -62,
    47282 => -62,
    47283 => -62,
    47284 => -62,
    47285 => -62,
    47286 => -62,
    47287 => -62,
    47288 => -62,
    47289 => -62,
    47290 => -62,
    47291 => -62,
    47292 => -62,
    47293 => -62,
    47294 => -62,
    47295 => -62,
    47296 => -62,
    47297 => -62,
    47298 => -62,
    47299 => -62,
    47300 => -62,
    47301 => -62,
    47302 => -62,
    47303 => -62,
    47304 => -62,
    47305 => -62,
    47306 => -62,
    47307 => -62,
    47308 => -62,
    47309 => -62,
    47310 => -62,
    47311 => -62,
    47312 => -62,
    47313 => -62,
    47314 => -62,
    47315 => -62,
    47316 => -62,
    47317 => -62,
    47318 => -62,
    47319 => -62,
    47320 => -62,
    47321 => -62,
    47322 => -62,
    47323 => -62,
    47324 => -62,
    47325 => -62,
    47326 => -62,
    47327 => -62,
    47328 => -62,
    47329 => -62,
    47330 => -62,
    47331 => -62,
    47332 => -62,
    47333 => -62,
    47334 => -62,
    47335 => -62,
    47336 => -62,
    47337 => -62,
    47338 => -62,
    47339 => -62,
    47340 => -62,
    47341 => -62,
    47342 => -62,
    47343 => -62,
    47344 => -62,
    47345 => -62,
    47346 => -62,
    47347 => -62,
    47348 => -62,
    47349 => -62,
    47350 => -62,
    47351 => -62,
    47352 => -62,
    47353 => -62,
    47354 => -62,
    47355 => -62,
    47356 => -62,
    47357 => -62,
    47358 => -62,
    47359 => -62,
    47360 => -62,
    47361 => -62,
    47362 => -62,
    47363 => -62,
    47364 => -62,
    47365 => -62,
    47366 => -62,
    47367 => -62,
    47368 => -62,
    47369 => -62,
    47370 => -62,
    47371 => -62,
    47372 => -62,
    47373 => -62,
    47374 => -62,
    47375 => -62,
    47376 => -62,
    47377 => -62,
    47378 => -62,
    47379 => -62,
    47380 => -62,
    47381 => -62,
    47382 => -62,
    47383 => -62,
    47384 => -62,
    47385 => -62,
    47386 => -62,
    47387 => -62,
    47388 => -62,
    47389 => -62,
    47390 => -62,
    47391 => -62,
    47392 => -62,
    47393 => -62,
    47394 => -62,
    47395 => -62,
    47396 => -62,
    47397 => -62,
    47398 => -62,
    47399 => -62,
    47400 => -62,
    47401 => -62,
    47402 => -62,
    47403 => -62,
    47404 => -62,
    47405 => -62,
    47406 => -62,
    47407 => -62,
    47408 => -62,
    47409 => -62,
    47410 => -62,
    47411 => -62,
    47412 => -62,
    47413 => -62,
    47414 => -62,
    47415 => -62,
    47416 => -62,
    47417 => -62,
    47418 => -62,
    47419 => -62,
    47420 => -62,
    47421 => -62,
    47422 => -62,
    47423 => -62,
    47424 => -62,
    47425 => -62,
    47426 => -62,
    47427 => -62,
    47428 => -62,
    47429 => -62,
    47430 => -62,
    47431 => -62,
    47432 => -62,
    47433 => -62,
    47434 => -62,
    47435 => -62,
    47436 => -62,
    47437 => -62,
    47438 => -62,
    47439 => -62,
    47440 => -62,
    47441 => -62,
    47442 => -62,
    47443 => -62,
    47444 => -62,
    47445 => -62,
    47446 => -62,
    47447 => -62,
    47448 => -62,
    47449 => -62,
    47450 => -62,
    47451 => -62,
    47452 => -62,
    47453 => -62,
    47454 => -62,
    47455 => -62,
    47456 => -62,
    47457 => -62,
    47458 => -62,
    47459 => -62,
    47460 => -62,
    47461 => -62,
    47462 => -62,
    47463 => -62,
    47464 => -62,
    47465 => -62,
    47466 => -62,
    47467 => -62,
    47468 => -62,
    47469 => -62,
    47470 => -62,
    47471 => -62,
    47472 => -62,
    47473 => -62,
    47474 => -62,
    47475 => -62,
    47476 => -62,
    47477 => -62,
    47478 => -62,
    47479 => -62,
    47480 => -62,
    47481 => -62,
    47482 => -62,
    47483 => -62,
    47484 => -62,
    47485 => -62,
    47486 => -62,
    47487 => -62,
    47488 => -62,
    47489 => -62,
    47490 => -62,
    47491 => -62,
    47492 => -62,
    47493 => -62,
    47494 => -62,
    47495 => -62,
    47496 => -62,
    47497 => -62,
    47498 => -62,
    47499 => -62,
    47500 => -62,
    47501 => -62,
    47502 => -62,
    47503 => -62,
    47504 => -62,
    47505 => -62,
    47506 => -62,
    47507 => -62,
    47508 => -62,
    47509 => -62,
    47510 => -62,
    47511 => -62,
    47512 => -62,
    47513 => -62,
    47514 => -62,
    47515 => -62,
    47516 => -62,
    47517 => -62,
    47518 => -62,
    47519 => -62,
    47520 => -62,
    47521 => -62,
    47522 => -62,
    47523 => -62,
    47524 => -62,
    47525 => -62,
    47526 => -62,
    47527 => -62,
    47528 => -62,
    47529 => -62,
    47530 => -62,
    47531 => -62,
    47532 => -62,
    47533 => -62,
    47534 => -62,
    47535 => -62,
    47536 => -62,
    47537 => -62,
    47538 => -62,
    47539 => -62,
    47540 => -62,
    47541 => -62,
    47542 => -62,
    47543 => -62,
    47544 => -62,
    47545 => -62,
    47546 => -62,
    47547 => -62,
    47548 => -62,
    47549 => -62,
    47550 => -62,
    47551 => -62,
    47552 => -62,
    47553 => -62,
    47554 => -62,
    47555 => -62,
    47556 => -62,
    47557 => -62,
    47558 => -62,
    47559 => -62,
    47560 => -62,
    47561 => -62,
    47562 => -62,
    47563 => -62,
    47564 => -62,
    47565 => -62,
    47566 => -62,
    47567 => -62,
    47568 => -62,
    47569 => -62,
    47570 => -62,
    47571 => -62,
    47572 => -62,
    47573 => -62,
    47574 => -62,
    47575 => -62,
    47576 => -62,
    47577 => -62,
    47578 => -62,
    47579 => -62,
    47580 => -62,
    47581 => -62,
    47582 => -62,
    47583 => -62,
    47584 => -62,
    47585 => -62,
    47586 => -62,
    47587 => -62,
    47588 => -62,
    47589 => -62,
    47590 => -62,
    47591 => -62,
    47592 => -62,
    47593 => -62,
    47594 => -62,
    47595 => -62,
    47596 => -62,
    47597 => -62,
    47598 => -62,
    47599 => -62,
    47600 => -62,
    47601 => -62,
    47602 => -62,
    47603 => -62,
    47604 => -62,
    47605 => -62,
    47606 => -62,
    47607 => -62,
    47608 => -62,
    47609 => -62,
    47610 => -62,
    47611 => -62,
    47612 => -62,
    47613 => -62,
    47614 => -62,
    47615 => -62,
    47616 => -62,
    47617 => -62,
    47618 => -62,
    47619 => -62,
    47620 => -62,
    47621 => -62,
    47622 => -62,
    47623 => -62,
    47624 => -62,
    47625 => -62,
    47626 => -62,
    47627 => -62,
    47628 => -62,
    47629 => -62,
    47630 => -62,
    47631 => -62,
    47632 => -62,
    47633 => -62,
    47634 => -62,
    47635 => -62,
    47636 => -62,
    47637 => -62,
    47638 => -62,
    47639 => -62,
    47640 => -62,
    47641 => -62,
    47642 => -62,
    47643 => -62,
    47644 => -62,
    47645 => -62,
    47646 => -62,
    47647 => -62,
    47648 => -62,
    47649 => -62,
    47650 => -62,
    47651 => -62,
    47652 => -62,
    47653 => -62,
    47654 => -62,
    47655 => -62,
    47656 => -62,
    47657 => -62,
    47658 => -62,
    47659 => -62,
    47660 => -62,
    47661 => -62,
    47662 => -62,
    47663 => -62,
    47664 => -62,
    47665 => -62,
    47666 => -62,
    47667 => -62,
    47668 => -62,
    47669 => -62,
    47670 => -62,
    47671 => -62,
    47672 => -62,
    47673 => -62,
    47674 => -62,
    47675 => -62,
    47676 => -62,
    47677 => -62,
    47678 => -62,
    47679 => -62,
    47680 => -62,
    47681 => -62,
    47682 => -62,
    47683 => -62,
    47684 => -62,
    47685 => -62,
    47686 => -62,
    47687 => -62,
    47688 => -62,
    47689 => -62,
    47690 => -62,
    47691 => -62,
    47692 => -62,
    47693 => -62,
    47694 => -62,
    47695 => -62,
    47696 => -62,
    47697 => -62,
    47698 => -62,
    47699 => -62,
    47700 => -62,
    47701 => -62,
    47702 => -62,
    47703 => -62,
    47704 => -62,
    47705 => -62,
    47706 => -62,
    47707 => -62,
    47708 => -62,
    47709 => -62,
    47710 => -62,
    47711 => -62,
    47712 => -62,
    47713 => -62,
    47714 => -62,
    47715 => -62,
    47716 => -62,
    47717 => -62,
    47718 => -62,
    47719 => -62,
    47720 => -62,
    47721 => -62,
    47722 => -62,
    47723 => -62,
    47724 => -62,
    47725 => -62,
    47726 => -62,
    47727 => -62,
    47728 => -62,
    47729 => -62,
    47730 => -62,
    47731 => -62,
    47732 => -62,
    47733 => -62,
    47734 => -62,
    47735 => -62,
    47736 => -62,
    47737 => -62,
    47738 => -62,
    47739 => -62,
    47740 => -62,
    47741 => -62,
    47742 => -62,
    47743 => -62,
    47744 => -62,
    47745 => -62,
    47746 => -62,
    47747 => -62,
    47748 => -62,
    47749 => -62,
    47750 => -62,
    47751 => -62,
    47752 => -62,
    47753 => -62,
    47754 => -62,
    47755 => -62,
    47756 => -62,
    47757 => -62,
    47758 => -62,
    47759 => -62,
    47760 => -62,
    47761 => -62,
    47762 => -62,
    47763 => -62,
    47764 => -62,
    47765 => -62,
    47766 => -62,
    47767 => -62,
    47768 => -62,
    47769 => -62,
    47770 => -62,
    47771 => -62,
    47772 => -62,
    47773 => -62,
    47774 => -62,
    47775 => -62,
    47776 => -62,
    47777 => -62,
    47778 => -62,
    47779 => -62,
    47780 => -62,
    47781 => -62,
    47782 => -62,
    47783 => -62,
    47784 => -62,
    47785 => -62,
    47786 => -62,
    47787 => -62,
    47788 => -62,
    47789 => -62,
    47790 => -62,
    47791 => -62,
    47792 => -62,
    47793 => -62,
    47794 => -62,
    47795 => -62,
    47796 => -62,
    47797 => -62,
    47798 => -62,
    47799 => -62,
    47800 => -62,
    47801 => -62,
    47802 => -62,
    47803 => -62,
    47804 => -62,
    47805 => -62,
    47806 => -62,
    47807 => -62,
    47808 => -62,
    47809 => -62,
    47810 => -62,
    47811 => -62,
    47812 => -62,
    47813 => -62,
    47814 => -62,
    47815 => -62,
    47816 => -62,
    47817 => -62,
    47818 => -62,
    47819 => -62,
    47820 => -62,
    47821 => -62,
    47822 => -62,
    47823 => -62,
    47824 => -62,
    47825 => -62,
    47826 => -62,
    47827 => -62,
    47828 => -62,
    47829 => -62,
    47830 => -62,
    47831 => -62,
    47832 => -62,
    47833 => -62,
    47834 => -62,
    47835 => -62,
    47836 => -62,
    47837 => -62,
    47838 => -63,
    47839 => -63,
    47840 => -63,
    47841 => -63,
    47842 => -63,
    47843 => -63,
    47844 => -63,
    47845 => -63,
    47846 => -63,
    47847 => -63,
    47848 => -63,
    47849 => -63,
    47850 => -63,
    47851 => -63,
    47852 => -63,
    47853 => -63,
    47854 => -63,
    47855 => -63,
    47856 => -63,
    47857 => -63,
    47858 => -63,
    47859 => -63,
    47860 => -63,
    47861 => -63,
    47862 => -63,
    47863 => -63,
    47864 => -63,
    47865 => -63,
    47866 => -63,
    47867 => -63,
    47868 => -63,
    47869 => -63,
    47870 => -63,
    47871 => -63,
    47872 => -63,
    47873 => -63,
    47874 => -63,
    47875 => -63,
    47876 => -63,
    47877 => -63,
    47878 => -63,
    47879 => -63,
    47880 => -63,
    47881 => -63,
    47882 => -63,
    47883 => -63,
    47884 => -63,
    47885 => -63,
    47886 => -63,
    47887 => -63,
    47888 => -63,
    47889 => -63,
    47890 => -63,
    47891 => -63,
    47892 => -63,
    47893 => -63,
    47894 => -63,
    47895 => -63,
    47896 => -63,
    47897 => -63,
    47898 => -63,
    47899 => -63,
    47900 => -63,
    47901 => -63,
    47902 => -63,
    47903 => -63,
    47904 => -63,
    47905 => -63,
    47906 => -63,
    47907 => -63,
    47908 => -63,
    47909 => -63,
    47910 => -63,
    47911 => -63,
    47912 => -63,
    47913 => -63,
    47914 => -63,
    47915 => -63,
    47916 => -63,
    47917 => -63,
    47918 => -63,
    47919 => -63,
    47920 => -63,
    47921 => -63,
    47922 => -63,
    47923 => -63,
    47924 => -63,
    47925 => -63,
    47926 => -63,
    47927 => -63,
    47928 => -63,
    47929 => -63,
    47930 => -63,
    47931 => -63,
    47932 => -63,
    47933 => -63,
    47934 => -63,
    47935 => -63,
    47936 => -63,
    47937 => -63,
    47938 => -63,
    47939 => -63,
    47940 => -63,
    47941 => -63,
    47942 => -63,
    47943 => -63,
    47944 => -63,
    47945 => -63,
    47946 => -63,
    47947 => -63,
    47948 => -63,
    47949 => -63,
    47950 => -63,
    47951 => -63,
    47952 => -63,
    47953 => -63,
    47954 => -63,
    47955 => -63,
    47956 => -63,
    47957 => -63,
    47958 => -63,
    47959 => -63,
    47960 => -63,
    47961 => -63,
    47962 => -63,
    47963 => -63,
    47964 => -63,
    47965 => -63,
    47966 => -63,
    47967 => -63,
    47968 => -63,
    47969 => -63,
    47970 => -63,
    47971 => -63,
    47972 => -63,
    47973 => -63,
    47974 => -63,
    47975 => -63,
    47976 => -63,
    47977 => -63,
    47978 => -63,
    47979 => -63,
    47980 => -63,
    47981 => -63,
    47982 => -63,
    47983 => -63,
    47984 => -63,
    47985 => -63,
    47986 => -63,
    47987 => -63,
    47988 => -63,
    47989 => -63,
    47990 => -63,
    47991 => -63,
    47992 => -63,
    47993 => -63,
    47994 => -63,
    47995 => -63,
    47996 => -63,
    47997 => -63,
    47998 => -63,
    47999 => -63,
    48000 => -63,
    48001 => -63,
    48002 => -63,
    48003 => -63,
    48004 => -63,
    48005 => -63,
    48006 => -63,
    48007 => -63,
    48008 => -63,
    48009 => -63,
    48010 => -63,
    48011 => -63,
    48012 => -63,
    48013 => -63,
    48014 => -63,
    48015 => -63,
    48016 => -63,
    48017 => -63,
    48018 => -63,
    48019 => -63,
    48020 => -63,
    48021 => -63,
    48022 => -63,
    48023 => -63,
    48024 => -63,
    48025 => -63,
    48026 => -63,
    48027 => -63,
    48028 => -63,
    48029 => -63,
    48030 => -63,
    48031 => -63,
    48032 => -63,
    48033 => -63,
    48034 => -63,
    48035 => -63,
    48036 => -63,
    48037 => -63,
    48038 => -63,
    48039 => -63,
    48040 => -63,
    48041 => -63,
    48042 => -63,
    48043 => -63,
    48044 => -63,
    48045 => -63,
    48046 => -63,
    48047 => -63,
    48048 => -63,
    48049 => -63,
    48050 => -63,
    48051 => -63,
    48052 => -63,
    48053 => -63,
    48054 => -63,
    48055 => -63,
    48056 => -63,
    48057 => -63,
    48058 => -63,
    48059 => -63,
    48060 => -63,
    48061 => -63,
    48062 => -63,
    48063 => -63,
    48064 => -63,
    48065 => -63,
    48066 => -63,
    48067 => -63,
    48068 => -63,
    48069 => -63,
    48070 => -63,
    48071 => -63,
    48072 => -63,
    48073 => -63,
    48074 => -63,
    48075 => -63,
    48076 => -63,
    48077 => -63,
    48078 => -63,
    48079 => -63,
    48080 => -63,
    48081 => -63,
    48082 => -63,
    48083 => -63,
    48084 => -63,
    48085 => -63,
    48086 => -63,
    48087 => -63,
    48088 => -63,
    48089 => -63,
    48090 => -63,
    48091 => -63,
    48092 => -63,
    48093 => -63,
    48094 => -63,
    48095 => -63,
    48096 => -63,
    48097 => -63,
    48098 => -63,
    48099 => -63,
    48100 => -63,
    48101 => -63,
    48102 => -63,
    48103 => -63,
    48104 => -63,
    48105 => -63,
    48106 => -63,
    48107 => -63,
    48108 => -63,
    48109 => -63,
    48110 => -63,
    48111 => -63,
    48112 => -63,
    48113 => -63,
    48114 => -63,
    48115 => -63,
    48116 => -63,
    48117 => -63,
    48118 => -63,
    48119 => -63,
    48120 => -63,
    48121 => -63,
    48122 => -63,
    48123 => -63,
    48124 => -63,
    48125 => -63,
    48126 => -63,
    48127 => -63,
    48128 => -63,
    48129 => -63,
    48130 => -63,
    48131 => -63,
    48132 => -63,
    48133 => -63,
    48134 => -63,
    48135 => -63,
    48136 => -63,
    48137 => -63,
    48138 => -63,
    48139 => -63,
    48140 => -63,
    48141 => -63,
    48142 => -63,
    48143 => -63,
    48144 => -63,
    48145 => -63,
    48146 => -63,
    48147 => -63,
    48148 => -63,
    48149 => -63,
    48150 => -63,
    48151 => -63,
    48152 => -63,
    48153 => -63,
    48154 => -63,
    48155 => -63,
    48156 => -63,
    48157 => -63,
    48158 => -63,
    48159 => -63,
    48160 => -63,
    48161 => -63,
    48162 => -63,
    48163 => -63,
    48164 => -63,
    48165 => -63,
    48166 => -63,
    48167 => -63,
    48168 => -63,
    48169 => -63,
    48170 => -63,
    48171 => -63,
    48172 => -63,
    48173 => -63,
    48174 => -63,
    48175 => -63,
    48176 => -63,
    48177 => -63,
    48178 => -63,
    48179 => -63,
    48180 => -63,
    48181 => -63,
    48182 => -63,
    48183 => -63,
    48184 => -63,
    48185 => -63,
    48186 => -63,
    48187 => -63,
    48188 => -63,
    48189 => -63,
    48190 => -63,
    48191 => -63,
    48192 => -63,
    48193 => -63,
    48194 => -63,
    48195 => -63,
    48196 => -63,
    48197 => -63,
    48198 => -63,
    48199 => -63,
    48200 => -63,
    48201 => -63,
    48202 => -63,
    48203 => -63,
    48204 => -63,
    48205 => -63,
    48206 => -63,
    48207 => -63,
    48208 => -63,
    48209 => -63,
    48210 => -63,
    48211 => -63,
    48212 => -63,
    48213 => -63,
    48214 => -63,
    48215 => -63,
    48216 => -63,
    48217 => -63,
    48218 => -63,
    48219 => -63,
    48220 => -63,
    48221 => -63,
    48222 => -63,
    48223 => -63,
    48224 => -63,
    48225 => -63,
    48226 => -63,
    48227 => -63,
    48228 => -63,
    48229 => -63,
    48230 => -63,
    48231 => -63,
    48232 => -63,
    48233 => -63,
    48234 => -63,
    48235 => -63,
    48236 => -63,
    48237 => -63,
    48238 => -63,
    48239 => -63,
    48240 => -63,
    48241 => -63,
    48242 => -63,
    48243 => -63,
    48244 => -63,
    48245 => -63,
    48246 => -63,
    48247 => -63,
    48248 => -63,
    48249 => -63,
    48250 => -63,
    48251 => -63,
    48252 => -63,
    48253 => -63,
    48254 => -63,
    48255 => -63,
    48256 => -63,
    48257 => -63,
    48258 => -63,
    48259 => -63,
    48260 => -63,
    48261 => -63,
    48262 => -63,
    48263 => -63,
    48264 => -63,
    48265 => -63,
    48266 => -63,
    48267 => -63,
    48268 => -63,
    48269 => -63,
    48270 => -63,
    48271 => -63,
    48272 => -63,
    48273 => -63,
    48274 => -63,
    48275 => -63,
    48276 => -63,
    48277 => -63,
    48278 => -63,
    48279 => -63,
    48280 => -63,
    48281 => -63,
    48282 => -63,
    48283 => -63,
    48284 => -63,
    48285 => -63,
    48286 => -63,
    48287 => -63,
    48288 => -63,
    48289 => -63,
    48290 => -63,
    48291 => -63,
    48292 => -63,
    48293 => -63,
    48294 => -63,
    48295 => -63,
    48296 => -63,
    48297 => -63,
    48298 => -63,
    48299 => -63,
    48300 => -63,
    48301 => -63,
    48302 => -63,
    48303 => -63,
    48304 => -63,
    48305 => -63,
    48306 => -63,
    48307 => -63,
    48308 => -63,
    48309 => -63,
    48310 => -63,
    48311 => -63,
    48312 => -63,
    48313 => -63,
    48314 => -63,
    48315 => -63,
    48316 => -63,
    48317 => -63,
    48318 => -63,
    48319 => -63,
    48320 => -63,
    48321 => -63,
    48322 => -63,
    48323 => -63,
    48324 => -63,
    48325 => -63,
    48326 => -63,
    48327 => -63,
    48328 => -63,
    48329 => -63,
    48330 => -63,
    48331 => -63,
    48332 => -63,
    48333 => -63,
    48334 => -63,
    48335 => -63,
    48336 => -63,
    48337 => -63,
    48338 => -63,
    48339 => -63,
    48340 => -63,
    48341 => -63,
    48342 => -63,
    48343 => -63,
    48344 => -63,
    48345 => -63,
    48346 => -63,
    48347 => -63,
    48348 => -63,
    48349 => -63,
    48350 => -63,
    48351 => -63,
    48352 => -63,
    48353 => -63,
    48354 => -63,
    48355 => -63,
    48356 => -63,
    48357 => -63,
    48358 => -63,
    48359 => -63,
    48360 => -63,
    48361 => -63,
    48362 => -63,
    48363 => -63,
    48364 => -63,
    48365 => -63,
    48366 => -63,
    48367 => -63,
    48368 => -63,
    48369 => -63,
    48370 => -63,
    48371 => -63,
    48372 => -63,
    48373 => -63,
    48374 => -63,
    48375 => -63,
    48376 => -63,
    48377 => -63,
    48378 => -63,
    48379 => -63,
    48380 => -63,
    48381 => -63,
    48382 => -63,
    48383 => -63,
    48384 => -63,
    48385 => -63,
    48386 => -63,
    48387 => -63,
    48388 => -63,
    48389 => -63,
    48390 => -63,
    48391 => -63,
    48392 => -63,
    48393 => -63,
    48394 => -63,
    48395 => -63,
    48396 => -63,
    48397 => -63,
    48398 => -63,
    48399 => -63,
    48400 => -63,
    48401 => -63,
    48402 => -63,
    48403 => -63,
    48404 => -63,
    48405 => -63,
    48406 => -63,
    48407 => -63,
    48408 => -63,
    48409 => -63,
    48410 => -63,
    48411 => -63,
    48412 => -63,
    48413 => -63,
    48414 => -63,
    48415 => -63,
    48416 => -63,
    48417 => -63,
    48418 => -63,
    48419 => -63,
    48420 => -63,
    48421 => -63,
    48422 => -63,
    48423 => -63,
    48424 => -63,
    48425 => -63,
    48426 => -63,
    48427 => -63,
    48428 => -63,
    48429 => -63,
    48430 => -63,
    48431 => -63,
    48432 => -63,
    48433 => -63,
    48434 => -63,
    48435 => -63,
    48436 => -63,
    48437 => -63,
    48438 => -63,
    48439 => -63,
    48440 => -63,
    48441 => -63,
    48442 => -63,
    48443 => -63,
    48444 => -63,
    48445 => -63,
    48446 => -63,
    48447 => -63,
    48448 => -63,
    48449 => -63,
    48450 => -63,
    48451 => -63,
    48452 => -63,
    48453 => -63,
    48454 => -63,
    48455 => -63,
    48456 => -63,
    48457 => -63,
    48458 => -63,
    48459 => -63,
    48460 => -63,
    48461 => -63,
    48462 => -63,
    48463 => -63,
    48464 => -63,
    48465 => -63,
    48466 => -63,
    48467 => -63,
    48468 => -63,
    48469 => -63,
    48470 => -63,
    48471 => -63,
    48472 => -63,
    48473 => -63,
    48474 => -63,
    48475 => -63,
    48476 => -63,
    48477 => -63,
    48478 => -63,
    48479 => -63,
    48480 => -63,
    48481 => -63,
    48482 => -63,
    48483 => -63,
    48484 => -63,
    48485 => -63,
    48486 => -63,
    48487 => -63,
    48488 => -63,
    48489 => -63,
    48490 => -63,
    48491 => -63,
    48492 => -63,
    48493 => -63,
    48494 => -63,
    48495 => -63,
    48496 => -63,
    48497 => -63,
    48498 => -63,
    48499 => -63,
    48500 => -63,
    48501 => -63,
    48502 => -63,
    48503 => -63,
    48504 => -63,
    48505 => -63,
    48506 => -63,
    48507 => -63,
    48508 => -63,
    48509 => -63,
    48510 => -63,
    48511 => -63,
    48512 => -63,
    48513 => -63,
    48514 => -63,
    48515 => -63,
    48516 => -63,
    48517 => -63,
    48518 => -63,
    48519 => -63,
    48520 => -63,
    48521 => -63,
    48522 => -63,
    48523 => -63,
    48524 => -63,
    48525 => -63,
    48526 => -63,
    48527 => -63,
    48528 => -63,
    48529 => -63,
    48530 => -63,
    48531 => -63,
    48532 => -63,
    48533 => -63,
    48534 => -63,
    48535 => -63,
    48536 => -63,
    48537 => -63,
    48538 => -63,
    48539 => -63,
    48540 => -63,
    48541 => -63,
    48542 => -63,
    48543 => -63,
    48544 => -63,
    48545 => -63,
    48546 => -63,
    48547 => -63,
    48548 => -63,
    48549 => -63,
    48550 => -63,
    48551 => -63,
    48552 => -63,
    48553 => -63,
    48554 => -63,
    48555 => -63,
    48556 => -63,
    48557 => -63,
    48558 => -63,
    48559 => -63,
    48560 => -63,
    48561 => -63,
    48562 => -63,
    48563 => -63,
    48564 => -63,
    48565 => -63,
    48566 => -63,
    48567 => -63,
    48568 => -63,
    48569 => -63,
    48570 => -63,
    48571 => -63,
    48572 => -63,
    48573 => -63,
    48574 => -63,
    48575 => -63,
    48576 => -63,
    48577 => -63,
    48578 => -63,
    48579 => -63,
    48580 => -63,
    48581 => -63,
    48582 => -63,
    48583 => -63,
    48584 => -63,
    48585 => -63,
    48586 => -63,
    48587 => -63,
    48588 => -63,
    48589 => -63,
    48590 => -63,
    48591 => -63,
    48592 => -63,
    48593 => -63,
    48594 => -63,
    48595 => -63,
    48596 => -63,
    48597 => -63,
    48598 => -63,
    48599 => -63,
    48600 => -63,
    48601 => -63,
    48602 => -63,
    48603 => -63,
    48604 => -63,
    48605 => -63,
    48606 => -63,
    48607 => -63,
    48608 => -63,
    48609 => -63,
    48610 => -63,
    48611 => -63,
    48612 => -63,
    48613 => -63,
    48614 => -63,
    48615 => -63,
    48616 => -63,
    48617 => -63,
    48618 => -63,
    48619 => -63,
    48620 => -63,
    48621 => -63,
    48622 => -63,
    48623 => -63,
    48624 => -63,
    48625 => -63,
    48626 => -63,
    48627 => -63,
    48628 => -63,
    48629 => -63,
    48630 => -63,
    48631 => -63,
    48632 => -63,
    48633 => -63,
    48634 => -63,
    48635 => -63,
    48636 => -63,
    48637 => -63,
    48638 => -63,
    48639 => -63,
    48640 => -63,
    48641 => -63,
    48642 => -63,
    48643 => -63,
    48644 => -63,
    48645 => -63,
    48646 => -63,
    48647 => -63,
    48648 => -63,
    48649 => -63,
    48650 => -63,
    48651 => -63,
    48652 => -63,
    48653 => -63,
    48654 => -63,
    48655 => -63,
    48656 => -63,
    48657 => -63,
    48658 => -63,
    48659 => -63,
    48660 => -63,
    48661 => -63,
    48662 => -63,
    48663 => -63,
    48664 => -63,
    48665 => -63,
    48666 => -63,
    48667 => -63,
    48668 => -63,
    48669 => -63,
    48670 => -63,
    48671 => -63,
    48672 => -63,
    48673 => -63,
    48674 => -63,
    48675 => -63,
    48676 => -63,
    48677 => -63,
    48678 => -63,
    48679 => -63,
    48680 => -63,
    48681 => -63,
    48682 => -63,
    48683 => -63,
    48684 => -63,
    48685 => -63,
    48686 => -63,
    48687 => -63,
    48688 => -63,
    48689 => -63,
    48690 => -63,
    48691 => -63,
    48692 => -63,
    48693 => -63,
    48694 => -63,
    48695 => -63,
    48696 => -63,
    48697 => -63,
    48698 => -63,
    48699 => -63,
    48700 => -63,
    48701 => -63,
    48702 => -63,
    48703 => -63,
    48704 => -63,
    48705 => -63,
    48706 => -63,
    48707 => -63,
    48708 => -63,
    48709 => -63,
    48710 => -63,
    48711 => -63,
    48712 => -63,
    48713 => -63,
    48714 => -63,
    48715 => -63,
    48716 => -63,
    48717 => -63,
    48718 => -63,
    48719 => -63,
    48720 => -63,
    48721 => -63,
    48722 => -63,
    48723 => -63,
    48724 => -63,
    48725 => -63,
    48726 => -63,
    48727 => -63,
    48728 => -63,
    48729 => -63,
    48730 => -63,
    48731 => -63,
    48732 => -63,
    48733 => -63,
    48734 => -63,
    48735 => -63,
    48736 => -63,
    48737 => -63,
    48738 => -63,
    48739 => -63,
    48740 => -63,
    48741 => -63,
    48742 => -63,
    48743 => -63,
    48744 => -63,
    48745 => -63,
    48746 => -63,
    48747 => -63,
    48748 => -63,
    48749 => -63,
    48750 => -63,
    48751 => -63,
    48752 => -63,
    48753 => -63,
    48754 => -63,
    48755 => -63,
    48756 => -63,
    48757 => -63,
    48758 => -63,
    48759 => -63,
    48760 => -63,
    48761 => -63,
    48762 => -63,
    48763 => -63,
    48764 => -63,
    48765 => -63,
    48766 => -63,
    48767 => -63,
    48768 => -63,
    48769 => -63,
    48770 => -63,
    48771 => -63,
    48772 => -63,
    48773 => -63,
    48774 => -63,
    48775 => -63,
    48776 => -63,
    48777 => -63,
    48778 => -63,
    48779 => -63,
    48780 => -63,
    48781 => -63,
    48782 => -63,
    48783 => -63,
    48784 => -63,
    48785 => -63,
    48786 => -63,
    48787 => -63,
    48788 => -63,
    48789 => -63,
    48790 => -63,
    48791 => -63,
    48792 => -63,
    48793 => -63,
    48794 => -63,
    48795 => -63,
    48796 => -63,
    48797 => -63,
    48798 => -63,
    48799 => -63,
    48800 => -63,
    48801 => -63,
    48802 => -63,
    48803 => -63,
    48804 => -63,
    48805 => -63,
    48806 => -63,
    48807 => -63,
    48808 => -63,
    48809 => -63,
    48810 => -63,
    48811 => -63,
    48812 => -63,
    48813 => -63,
    48814 => -63,
    48815 => -63,
    48816 => -63,
    48817 => -63,
    48818 => -63,
    48819 => -63,
    48820 => -63,
    48821 => -63,
    48822 => -63,
    48823 => -63,
    48824 => -63,
    48825 => -63,
    48826 => -63,
    48827 => -63,
    48828 => -63,
    48829 => -63,
    48830 => -63,
    48831 => -63,
    48832 => -63,
    48833 => -63,
    48834 => -63,
    48835 => -63,
    48836 => -63,
    48837 => -63,
    48838 => -63,
    48839 => -63,
    48840 => -63,
    48841 => -63,
    48842 => -63,
    48843 => -63,
    48844 => -63,
    48845 => -63,
    48846 => -63,
    48847 => -63,
    48848 => -63,
    48849 => -63,
    48850 => -63,
    48851 => -63,
    48852 => -63,
    48853 => -63,
    48854 => -63,
    48855 => -63,
    48856 => -63,
    48857 => -63,
    48858 => -63,
    48859 => -63,
    48860 => -63,
    48861 => -63,
    48862 => -63,
    48863 => -63,
    48864 => -63,
    48865 => -63,
    48866 => -63,
    48867 => -63,
    48868 => -63,
    48869 => -63,
    48870 => -63,
    48871 => -63,
    48872 => -63,
    48873 => -63,
    48874 => -63,
    48875 => -63,
    48876 => -63,
    48877 => -63,
    48878 => -63,
    48879 => -63,
    48880 => -63,
    48881 => -63,
    48882 => -63,
    48883 => -63,
    48884 => -63,
    48885 => -63,
    48886 => -63,
    48887 => -63,
    48888 => -63,
    48889 => -63,
    48890 => -63,
    48891 => -63,
    48892 => -63,
    48893 => -63,
    48894 => -63,
    48895 => -63,
    48896 => -63,
    48897 => -63,
    48898 => -63,
    48899 => -63,
    48900 => -63,
    48901 => -63,
    48902 => -63,
    48903 => -63,
    48904 => -63,
    48905 => -63,
    48906 => -63,
    48907 => -63,
    48908 => -63,
    48909 => -63,
    48910 => -63,
    48911 => -63,
    48912 => -63,
    48913 => -63,
    48914 => -63,
    48915 => -63,
    48916 => -63,
    48917 => -63,
    48918 => -63,
    48919 => -63,
    48920 => -63,
    48921 => -63,
    48922 => -63,
    48923 => -63,
    48924 => -63,
    48925 => -63,
    48926 => -63,
    48927 => -63,
    48928 => -63,
    48929 => -63,
    48930 => -63,
    48931 => -63,
    48932 => -63,
    48933 => -63,
    48934 => -63,
    48935 => -63,
    48936 => -63,
    48937 => -63,
    48938 => -63,
    48939 => -63,
    48940 => -63,
    48941 => -63,
    48942 => -63,
    48943 => -63,
    48944 => -63,
    48945 => -63,
    48946 => -63,
    48947 => -63,
    48948 => -63,
    48949 => -63,
    48950 => -63,
    48951 => -63,
    48952 => -63,
    48953 => -63,
    48954 => -63,
    48955 => -63,
    48956 => -63,
    48957 => -63,
    48958 => -63,
    48959 => -63,
    48960 => -63,
    48961 => -63,
    48962 => -63,
    48963 => -63,
    48964 => -63,
    48965 => -63,
    48966 => -63,
    48967 => -63,
    48968 => -63,
    48969 => -63,
    48970 => -63,
    48971 => -63,
    48972 => -63,
    48973 => -63,
    48974 => -63,
    48975 => -63,
    48976 => -63,
    48977 => -63,
    48978 => -63,
    48979 => -63,
    48980 => -63,
    48981 => -63,
    48982 => -63,
    48983 => -63,
    48984 => -63,
    48985 => -63,
    48986 => -63,
    48987 => -63,
    48988 => -63,
    48989 => -63,
    48990 => -63,
    48991 => -63,
    48992 => -63,
    48993 => -63,
    48994 => -63,
    48995 => -63,
    48996 => -63,
    48997 => -63,
    48998 => -63,
    48999 => -63,
    49000 => -63,
    49001 => -63,
    49002 => -63,
    49003 => -63,
    49004 => -63,
    49005 => -63,
    49006 => -63,
    49007 => -63,
    49008 => -63,
    49009 => -63,
    49010 => -63,
    49011 => -63,
    49012 => -63,
    49013 => -63,
    49014 => -63,
    49015 => -63,
    49016 => -63,
    49017 => -63,
    49018 => -63,
    49019 => -63,
    49020 => -63,
    49021 => -63,
    49022 => -63,
    49023 => -63,
    49024 => -63,
    49025 => -63,
    49026 => -63,
    49027 => -63,
    49028 => -63,
    49029 => -63,
    49030 => -63,
    49031 => -63,
    49032 => -63,
    49033 => -63,
    49034 => -63,
    49035 => -63,
    49036 => -63,
    49037 => -63,
    49038 => -63,
    49039 => -63,
    49040 => -63,
    49041 => -63,
    49042 => -63,
    49043 => -63,
    49044 => -63,
    49045 => -63,
    49046 => -63,
    49047 => -63,
    49048 => -63,
    49049 => -63,
    49050 => -63,
    49051 => -63,
    49052 => -63,
    49053 => -63,
    49054 => -63,
    49055 => -63,
    49056 => -63,
    49057 => -63,
    49058 => -63,
    49059 => -63,
    49060 => -63,
    49061 => -63,
    49062 => -63,
    49063 => -63,
    49064 => -63,
    49065 => -63,
    49066 => -63,
    49067 => -63,
    49068 => -63,
    49069 => -63,
    49070 => -63,
    49071 => -63,
    49072 => -63,
    49073 => -63,
    49074 => -63,
    49075 => -63,
    49076 => -63,
    49077 => -63,
    49078 => -63,
    49079 => -63,
    49080 => -63,
    49081 => -63,
    49082 => -63,
    49083 => -63,
    49084 => -63,
    49085 => -63,
    49086 => -63,
    49087 => -63,
    49088 => -63,
    49089 => -63,
    49090 => -63,
    49091 => -63,
    49092 => -63,
    49093 => -63,
    49094 => -63,
    49095 => -63,
    49096 => -63,
    49097 => -63,
    49098 => -63,
    49099 => -63,
    49100 => -63,
    49101 => -63,
    49102 => -63,
    49103 => -63,
    49104 => -63,
    49105 => -63,
    49106 => -63,
    49107 => -63,
    49108 => -63,
    49109 => -63,
    49110 => -63,
    49111 => -63,
    49112 => -63,
    49113 => -63,
    49114 => -63,
    49115 => -63,
    49116 => -63,
    49117 => -63,
    49118 => -63,
    49119 => -63,
    49120 => -63,
    49121 => -63,
    49122 => -63,
    49123 => -63,
    49124 => -63,
    49125 => -63,
    49126 => -63,
    49127 => -63,
    49128 => -63,
    49129 => -63,
    49130 => -63,
    49131 => -63,
    49132 => -63,
    49133 => -63,
    49134 => -63,
    49135 => -63,
    49136 => -63,
    49137 => -63,
    49138 => -63,
    49139 => -63,
    49140 => -63,
    49141 => -63,
    49142 => -63,
    49143 => -63,
    49144 => -63,
    49145 => -63,
    49146 => -63,
    49147 => -63,
    49148 => -63,
    49149 => -63,
    49150 => -63,
    49151 => -63,
    49152 => -63,
    49153 => -63,
    49154 => -63,
    49155 => -63,
    49156 => -63,
    49157 => -63,
    49158 => -63,
    49159 => -63,
    49160 => -63,
    49161 => -63,
    49162 => -63,
    49163 => -63,
    49164 => -63,
    49165 => -63,
    49166 => -63,
    49167 => -63,
    49168 => -63,
    49169 => -63,
    49170 => -63,
    49171 => -63,
    49172 => -63,
    49173 => -63,
    49174 => -63,
    49175 => -63,
    49176 => -63,
    49177 => -63,
    49178 => -63,
    49179 => -63,
    49180 => -63,
    49181 => -63,
    49182 => -63,
    49183 => -63,
    49184 => -63,
    49185 => -63,
    49186 => -63,
    49187 => -63,
    49188 => -63,
    49189 => -63,
    49190 => -63,
    49191 => -63,
    49192 => -63,
    49193 => -63,
    49194 => -63,
    49195 => -63,
    49196 => -63,
    49197 => -63,
    49198 => -63,
    49199 => -63,
    49200 => -63,
    49201 => -63,
    49202 => -63,
    49203 => -63,
    49204 => -63,
    49205 => -63,
    49206 => -63,
    49207 => -63,
    49208 => -63,
    49209 => -63,
    49210 => -63,
    49211 => -63,
    49212 => -63,
    49213 => -63,
    49214 => -63,
    49215 => -63,
    49216 => -63,
    49217 => -63,
    49218 => -63,
    49219 => -63,
    49220 => -63,
    49221 => -63,
    49222 => -63,
    49223 => -63,
    49224 => -63,
    49225 => -63,
    49226 => -63,
    49227 => -63,
    49228 => -63,
    49229 => -63,
    49230 => -63,
    49231 => -63,
    49232 => -63,
    49233 => -63,
    49234 => -63,
    49235 => -63,
    49236 => -63,
    49237 => -63,
    49238 => -63,
    49239 => -63,
    49240 => -63,
    49241 => -63,
    49242 => -63,
    49243 => -63,
    49244 => -63,
    49245 => -63,
    49246 => -63,
    49247 => -63,
    49248 => -63,
    49249 => -63,
    49250 => -63,
    49251 => -63,
    49252 => -63,
    49253 => -63,
    49254 => -63,
    49255 => -63,
    49256 => -63,
    49257 => -63,
    49258 => -63,
    49259 => -63,
    49260 => -63,
    49261 => -63,
    49262 => -63,
    49263 => -63,
    49264 => -63,
    49265 => -63,
    49266 => -63,
    49267 => -63,
    49268 => -63,
    49269 => -63,
    49270 => -63,
    49271 => -63,
    49272 => -63,
    49273 => -63,
    49274 => -63,
    49275 => -63,
    49276 => -63,
    49277 => -63,
    49278 => -63,
    49279 => -63,
    49280 => -63,
    49281 => -63,
    49282 => -63,
    49283 => -63,
    49284 => -63,
    49285 => -63,
    49286 => -63,
    49287 => -63,
    49288 => -63,
    49289 => -63,
    49290 => -63,
    49291 => -63,
    49292 => -63,
    49293 => -63,
    49294 => -63,
    49295 => -63,
    49296 => -63,
    49297 => -63,
    49298 => -63,
    49299 => -63,
    49300 => -63,
    49301 => -63,
    49302 => -63,
    49303 => -63,
    49304 => -63,
    49305 => -63,
    49306 => -63,
    49307 => -63,
    49308 => -63,
    49309 => -63,
    49310 => -63,
    49311 => -63,
    49312 => -63,
    49313 => -63,
    49314 => -63,
    49315 => -63,
    49316 => -63,
    49317 => -63,
    49318 => -63,
    49319 => -63,
    49320 => -63,
    49321 => -63,
    49322 => -63,
    49323 => -63,
    49324 => -63,
    49325 => -63,
    49326 => -63,
    49327 => -63,
    49328 => -63,
    49329 => -63,
    49330 => -63,
    49331 => -63,
    49332 => -63,
    49333 => -63,
    49334 => -63,
    49335 => -63,
    49336 => -63,
    49337 => -63,
    49338 => -63,
    49339 => -63,
    49340 => -63,
    49341 => -63,
    49342 => -63,
    49343 => -63,
    49344 => -63,
    49345 => -63,
    49346 => -63,
    49347 => -63,
    49348 => -63,
    49349 => -63,
    49350 => -63,
    49351 => -63,
    49352 => -63,
    49353 => -63,
    49354 => -63,
    49355 => -63,
    49356 => -63,
    49357 => -63,
    49358 => -63,
    49359 => -63,
    49360 => -63,
    49361 => -63,
    49362 => -63,
    49363 => -63,
    49364 => -63,
    49365 => -63,
    49366 => -63,
    49367 => -63,
    49368 => -63,
    49369 => -63,
    49370 => -63,
    49371 => -63,
    49372 => -63,
    49373 => -63,
    49374 => -63,
    49375 => -63,
    49376 => -63,
    49377 => -63,
    49378 => -63,
    49379 => -63,
    49380 => -63,
    49381 => -63,
    49382 => -63,
    49383 => -63,
    49384 => -63,
    49385 => -63,
    49386 => -63,
    49387 => -63,
    49388 => -63,
    49389 => -63,
    49390 => -63,
    49391 => -63,
    49392 => -63,
    49393 => -63,
    49394 => -63,
    49395 => -63,
    49396 => -63,
    49397 => -63,
    49398 => -63,
    49399 => -63,
    49400 => -63,
    49401 => -63,
    49402 => -63,
    49403 => -63,
    49404 => -63,
    49405 => -63,
    49406 => -63,
    49407 => -63,
    49408 => -63,
    49409 => -63,
    49410 => -63,
    49411 => -63,
    49412 => -63,
    49413 => -63,
    49414 => -63,
    49415 => -63,
    49416 => -63,
    49417 => -63,
    49418 => -63,
    49419 => -63,
    49420 => -63,
    49421 => -63,
    49422 => -63,
    49423 => -63,
    49424 => -63,
    49425 => -63,
    49426 => -63,
    49427 => -63,
    49428 => -63,
    49429 => -63,
    49430 => -63,
    49431 => -63,
    49432 => -63,
    49433 => -63,
    49434 => -63,
    49435 => -63,
    49436 => -63,
    49437 => -63,
    49438 => -63,
    49439 => -63,
    49440 => -63,
    49441 => -63,
    49442 => -63,
    49443 => -63,
    49444 => -63,
    49445 => -63,
    49446 => -63,
    49447 => -63,
    49448 => -63,
    49449 => -63,
    49450 => -63,
    49451 => -63,
    49452 => -63,
    49453 => -63,
    49454 => -63,
    49455 => -63,
    49456 => -63,
    49457 => -63,
    49458 => -63,
    49459 => -63,
    49460 => -63,
    49461 => -63,
    49462 => -63,
    49463 => -63,
    49464 => -63,
    49465 => -63,
    49466 => -63,
    49467 => -63,
    49468 => -63,
    49469 => -63,
    49470 => -63,
    49471 => -63,
    49472 => -63,
    49473 => -63,
    49474 => -63,
    49475 => -63,
    49476 => -63,
    49477 => -63,
    49478 => -63,
    49479 => -63,
    49480 => -63,
    49481 => -63,
    49482 => -63,
    49483 => -63,
    49484 => -63,
    49485 => -63,
    49486 => -63,
    49487 => -63,
    49488 => -63,
    49489 => -63,
    49490 => -63,
    49491 => -63,
    49492 => -63,
    49493 => -63,
    49494 => -63,
    49495 => -63,
    49496 => -63,
    49497 => -63,
    49498 => -63,
    49499 => -63,
    49500 => -63,
    49501 => -63,
    49502 => -63,
    49503 => -63,
    49504 => -63,
    49505 => -63,
    49506 => -63,
    49507 => -63,
    49508 => -63,
    49509 => -63,
    49510 => -63,
    49511 => -63,
    49512 => -63,
    49513 => -63,
    49514 => -63,
    49515 => -63,
    49516 => -63,
    49517 => -63,
    49518 => -63,
    49519 => -63,
    49520 => -63,
    49521 => -63,
    49522 => -63,
    49523 => -63,
    49524 => -63,
    49525 => -63,
    49526 => -63,
    49527 => -63,
    49528 => -63,
    49529 => -63,
    49530 => -63,
    49531 => -63,
    49532 => -63,
    49533 => -63,
    49534 => -63,
    49535 => -63,
    49536 => -63,
    49537 => -63,
    49538 => -63,
    49539 => -63,
    49540 => -63,
    49541 => -63,
    49542 => -63,
    49543 => -63,
    49544 => -63,
    49545 => -63,
    49546 => -63,
    49547 => -63,
    49548 => -63,
    49549 => -63,
    49550 => -63,
    49551 => -63,
    49552 => -63,
    49553 => -63,
    49554 => -63,
    49555 => -63,
    49556 => -63,
    49557 => -63,
    49558 => -63,
    49559 => -63,
    49560 => -63,
    49561 => -63,
    49562 => -63,
    49563 => -63,
    49564 => -63,
    49565 => -63,
    49566 => -63,
    49567 => -63,
    49568 => -63,
    49569 => -63,
    49570 => -63,
    49571 => -63,
    49572 => -63,
    49573 => -63,
    49574 => -63,
    49575 => -63,
    49576 => -63,
    49577 => -63,
    49578 => -63,
    49579 => -63,
    49580 => -63,
    49581 => -63,
    49582 => -63,
    49583 => -63,
    49584 => -63,
    49585 => -63,
    49586 => -63,
    49587 => -63,
    49588 => -63,
    49589 => -63,
    49590 => -63,
    49591 => -63,
    49592 => -63,
    49593 => -63,
    49594 => -63,
    49595 => -63,
    49596 => -63,
    49597 => -63,
    49598 => -63,
    49599 => -63,
    49600 => -63,
    49601 => -63,
    49602 => -63,
    49603 => -63,
    49604 => -63,
    49605 => -63,
    49606 => -63,
    49607 => -63,
    49608 => -63,
    49609 => -63,
    49610 => -63,
    49611 => -63,
    49612 => -63,
    49613 => -63,
    49614 => -63,
    49615 => -63,
    49616 => -63,
    49617 => -63,
    49618 => -63,
    49619 => -63,
    49620 => -63,
    49621 => -63,
    49622 => -63,
    49623 => -63,
    49624 => -63,
    49625 => -63,
    49626 => -63,
    49627 => -63,
    49628 => -63,
    49629 => -63,
    49630 => -63,
    49631 => -63,
    49632 => -63,
    49633 => -63,
    49634 => -63,
    49635 => -63,
    49636 => -63,
    49637 => -63,
    49638 => -63,
    49639 => -63,
    49640 => -63,
    49641 => -63,
    49642 => -63,
    49643 => -63,
    49644 => -63,
    49645 => -63,
    49646 => -63,
    49647 => -63,
    49648 => -63,
    49649 => -63,
    49650 => -63,
    49651 => -63,
    49652 => -63,
    49653 => -63,
    49654 => -63,
    49655 => -63,
    49656 => -63,
    49657 => -63,
    49658 => -63,
    49659 => -63,
    49660 => -63,
    49661 => -63,
    49662 => -63,
    49663 => -63,
    49664 => -63,
    49665 => -63,
    49666 => -63,
    49667 => -63,
    49668 => -63,
    49669 => -63,
    49670 => -63,
    49671 => -63,
    49672 => -63,
    49673 => -63,
    49674 => -63,
    49675 => -63,
    49676 => -63,
    49677 => -63,
    49678 => -63,
    49679 => -63,
    49680 => -63,
    49681 => -63,
    49682 => -63,
    49683 => -63,
    49684 => -63,
    49685 => -63,
    49686 => -63,
    49687 => -63,
    49688 => -63,
    49689 => -63,
    49690 => -63,
    49691 => -63,
    49692 => -63,
    49693 => -63,
    49694 => -63,
    49695 => -63,
    49696 => -63,
    49697 => -63,
    49698 => -63,
    49699 => -63,
    49700 => -63,
    49701 => -63,
    49702 => -63,
    49703 => -63,
    49704 => -63,
    49705 => -63,
    49706 => -63,
    49707 => -63,
    49708 => -63,
    49709 => -63,
    49710 => -63,
    49711 => -63,
    49712 => -63,
    49713 => -63,
    49714 => -63,
    49715 => -63,
    49716 => -63,
    49717 => -63,
    49718 => -63,
    49719 => -63,
    49720 => -63,
    49721 => -63,
    49722 => -63,
    49723 => -63,
    49724 => -63,
    49725 => -63,
    49726 => -63,
    49727 => -63,
    49728 => -63,
    49729 => -63,
    49730 => -63,
    49731 => -63,
    49732 => -63,
    49733 => -63,
    49734 => -63,
    49735 => -63,
    49736 => -63,
    49737 => -63,
    49738 => -63,
    49739 => -63,
    49740 => -63,
    49741 => -63,
    49742 => -63,
    49743 => -63,
    49744 => -63,
    49745 => -63,
    49746 => -63,
    49747 => -63,
    49748 => -63,
    49749 => -63,
    49750 => -63,
    49751 => -63,
    49752 => -63,
    49753 => -63,
    49754 => -63,
    49755 => -63,
    49756 => -63,
    49757 => -63,
    49758 => -63,
    49759 => -63,
    49760 => -63,
    49761 => -63,
    49762 => -63,
    49763 => -63,
    49764 => -63,
    49765 => -63,
    49766 => -63,
    49767 => -63,
    49768 => -63,
    49769 => -63,
    49770 => -63,
    49771 => -63,
    49772 => -63,
    49773 => -63,
    49774 => -63,
    49775 => -63,
    49776 => -63,
    49777 => -63,
    49778 => -63,
    49779 => -63,
    49780 => -63,
    49781 => -63,
    49782 => -63,
    49783 => -63,
    49784 => -63,
    49785 => -63,
    49786 => -63,
    49787 => -63,
    49788 => -63,
    49789 => -63,
    49790 => -63,
    49791 => -63,
    49792 => -63,
    49793 => -63,
    49794 => -63,
    49795 => -63,
    49796 => -63,
    49797 => -63,
    49798 => -63,
    49799 => -63,
    49800 => -63,
    49801 => -63,
    49802 => -63,
    49803 => -63,
    49804 => -63,
    49805 => -63,
    49806 => -63,
    49807 => -63,
    49808 => -63,
    49809 => -63,
    49810 => -63,
    49811 => -63,
    49812 => -63,
    49813 => -63,
    49814 => -63,
    49815 => -63,
    49816 => -63,
    49817 => -63,
    49818 => -63,
    49819 => -63,
    49820 => -63,
    49821 => -63,
    49822 => -63,
    49823 => -63,
    49824 => -63,
    49825 => -63,
    49826 => -63,
    49827 => -63,
    49828 => -63,
    49829 => -63,
    49830 => -63,
    49831 => -63,
    49832 => -63,
    49833 => -63,
    49834 => -63,
    49835 => -63,
    49836 => -63,
    49837 => -63,
    49838 => -63,
    49839 => -63,
    49840 => -63,
    49841 => -63,
    49842 => -63,
    49843 => -63,
    49844 => -63,
    49845 => -63,
    49846 => -63,
    49847 => -63,
    49848 => -63,
    49849 => -63,
    49850 => -63,
    49851 => -63,
    49852 => -63,
    49853 => -63,
    49854 => -63,
    49855 => -63,
    49856 => -63,
    49857 => -63,
    49858 => -63,
    49859 => -63,
    49860 => -63,
    49861 => -63,
    49862 => -63,
    49863 => -63,
    49864 => -63,
    49865 => -63,
    49866 => -63,
    49867 => -63,
    49868 => -63,
    49869 => -63,
    49870 => -63,
    49871 => -63,
    49872 => -63,
    49873 => -63,
    49874 => -63,
    49875 => -63,
    49876 => -63,
    49877 => -63,
    49878 => -63,
    49879 => -63,
    49880 => -63,
    49881 => -63,
    49882 => -63,
    49883 => -63,
    49884 => -63,
    49885 => -63,
    49886 => -63,
    49887 => -63,
    49888 => -63,
    49889 => -63,
    49890 => -63,
    49891 => -63,
    49892 => -63,
    49893 => -63,
    49894 => -63,
    49895 => -63,
    49896 => -63,
    49897 => -63,
    49898 => -63,
    49899 => -63,
    49900 => -63,
    49901 => -63,
    49902 => -63,
    49903 => -63,
    49904 => -63,
    49905 => -63,
    49906 => -63,
    49907 => -63,
    49908 => -63,
    49909 => -63,
    49910 => -63,
    49911 => -63,
    49912 => -63,
    49913 => -63,
    49914 => -63,
    49915 => -63,
    49916 => -63,
    49917 => -63,
    49918 => -63,
    49919 => -63,
    49920 => -63,
    49921 => -63,
    49922 => -63,
    49923 => -63,
    49924 => -63,
    49925 => -63,
    49926 => -63,
    49927 => -63,
    49928 => -63,
    49929 => -63,
    49930 => -63,
    49931 => -63,
    49932 => -63,
    49933 => -63,
    49934 => -63,
    49935 => -63,
    49936 => -63,
    49937 => -63,
    49938 => -63,
    49939 => -63,
    49940 => -63,
    49941 => -63,
    49942 => -63,
    49943 => -63,
    49944 => -63,
    49945 => -63,
    49946 => -63,
    49947 => -63,
    49948 => -63,
    49949 => -63,
    49950 => -63,
    49951 => -63,
    49952 => -63,
    49953 => -63,
    49954 => -63,
    49955 => -63,
    49956 => -63,
    49957 => -63,
    49958 => -63,
    49959 => -63,
    49960 => -63,
    49961 => -63,
    49962 => -63,
    49963 => -63,
    49964 => -63,
    49965 => -63,
    49966 => -63,
    49967 => -63,
    49968 => -63,
    49969 => -63,
    49970 => -63,
    49971 => -63,
    49972 => -63,
    49973 => -63,
    49974 => -63,
    49975 => -63,
    49976 => -63,
    49977 => -63,
    49978 => -63,
    49979 => -63,
    49980 => -63,
    49981 => -63,
    49982 => -63,
    49983 => -63,
    49984 => -63,
    49985 => -63,
    49986 => -63,
    49987 => -63,
    49988 => -63,
    49989 => -63,
    49990 => -63,
    49991 => -63,
    49992 => -63,
    49993 => -63,
    49994 => -63,
    49995 => -63,
    49996 => -63,
    49997 => -63,
    49998 => -63,
    49999 => -63,
    50000 => -63,
    50001 => -63,
    50002 => -63,
    50003 => -63,
    50004 => -63,
    50005 => -63,
    50006 => -63,
    50007 => -63,
    50008 => -63,
    50009 => -63,
    50010 => -63,
    50011 => -63,
    50012 => -63,
    50013 => -63,
    50014 => -63,
    50015 => -63,
    50016 => -63,
    50017 => -63,
    50018 => -63,
    50019 => -63,
    50020 => -63,
    50021 => -63,
    50022 => -63,
    50023 => -63,
    50024 => -63,
    50025 => -63,
    50026 => -63,
    50027 => -63,
    50028 => -63,
    50029 => -63,
    50030 => -63,
    50031 => -63,
    50032 => -63,
    50033 => -63,
    50034 => -63,
    50035 => -63,
    50036 => -63,
    50037 => -63,
    50038 => -63,
    50039 => -63,
    50040 => -63,
    50041 => -63,
    50042 => -63,
    50043 => -63,
    50044 => -63,
    50045 => -63,
    50046 => -63,
    50047 => -63,
    50048 => -63,
    50049 => -63,
    50050 => -63,
    50051 => -63,
    50052 => -63,
    50053 => -63,
    50054 => -63,
    50055 => -63,
    50056 => -63,
    50057 => -63,
    50058 => -63,
    50059 => -63,
    50060 => -63,
    50061 => -63,
    50062 => -63,
    50063 => -63,
    50064 => -63,
    50065 => -63,
    50066 => -63,
    50067 => -63,
    50068 => -63,
    50069 => -63,
    50070 => -63,
    50071 => -63,
    50072 => -63,
    50073 => -63,
    50074 => -63,
    50075 => -63,
    50076 => -63,
    50077 => -63,
    50078 => -63,
    50079 => -63,
    50080 => -63,
    50081 => -63,
    50082 => -63,
    50083 => -63,
    50084 => -63,
    50085 => -63,
    50086 => -63,
    50087 => -63,
    50088 => -63,
    50089 => -63,
    50090 => -63,
    50091 => -63,
    50092 => -63,
    50093 => -63,
    50094 => -63,
    50095 => -63,
    50096 => -63,
    50097 => -63,
    50098 => -63,
    50099 => -63,
    50100 => -63,
    50101 => -63,
    50102 => -63,
    50103 => -63,
    50104 => -63,
    50105 => -63,
    50106 => -63,
    50107 => -63,
    50108 => -63,
    50109 => -63,
    50110 => -63,
    50111 => -63,
    50112 => -63,
    50113 => -63,
    50114 => -63,
    50115 => -63,
    50116 => -63,
    50117 => -63,
    50118 => -63,
    50119 => -63,
    50120 => -63,
    50121 => -63,
    50122 => -63,
    50123 => -63,
    50124 => -63,
    50125 => -63,
    50126 => -63,
    50127 => -63,
    50128 => -63,
    50129 => -63,
    50130 => -63,
    50131 => -63,
    50132 => -63,
    50133 => -63,
    50134 => -63,
    50135 => -63,
    50136 => -63,
    50137 => -63,
    50138 => -63,
    50139 => -63,
    50140 => -63,
    50141 => -63,
    50142 => -63,
    50143 => -63,
    50144 => -63,
    50145 => -63,
    50146 => -63,
    50147 => -63,
    50148 => -63,
    50149 => -63,
    50150 => -63,
    50151 => -63,
    50152 => -63,
    50153 => -63,
    50154 => -63,
    50155 => -63,
    50156 => -63,
    50157 => -63,
    50158 => -63,
    50159 => -63,
    50160 => -63,
    50161 => -63,
    50162 => -63,
    50163 => -63,
    50164 => -63,
    50165 => -63,
    50166 => -63,
    50167 => -63,
    50168 => -63,
    50169 => -63,
    50170 => -63,
    50171 => -63,
    50172 => -63,
    50173 => -63,
    50174 => -63,
    50175 => -63,
    50176 => -63,
    50177 => -63,
    50178 => -63,
    50179 => -63,
    50180 => -63,
    50181 => -63,
    50182 => -63,
    50183 => -63,
    50184 => -63,
    50185 => -63,
    50186 => -63,
    50187 => -63,
    50188 => -63,
    50189 => -63,
    50190 => -63,
    50191 => -63,
    50192 => -63,
    50193 => -63,
    50194 => -63,
    50195 => -63,
    50196 => -63,
    50197 => -63,
    50198 => -63,
    50199 => -63,
    50200 => -63,
    50201 => -63,
    50202 => -63,
    50203 => -63,
    50204 => -63,
    50205 => -63,
    50206 => -63,
    50207 => -63,
    50208 => -63,
    50209 => -63,
    50210 => -63,
    50211 => -63,
    50212 => -63,
    50213 => -63,
    50214 => -63,
    50215 => -63,
    50216 => -63,
    50217 => -63,
    50218 => -63,
    50219 => -63,
    50220 => -63,
    50221 => -63,
    50222 => -63,
    50223 => -63,
    50224 => -63,
    50225 => -63,
    50226 => -63,
    50227 => -63,
    50228 => -63,
    50229 => -63,
    50230 => -63,
    50231 => -63,
    50232 => -63,
    50233 => -63,
    50234 => -63,
    50235 => -63,
    50236 => -63,
    50237 => -63,
    50238 => -63,
    50239 => -63,
    50240 => -63,
    50241 => -63,
    50242 => -63,
    50243 => -63,
    50244 => -63,
    50245 => -63,
    50246 => -63,
    50247 => -63,
    50248 => -63,
    50249 => -63,
    50250 => -63,
    50251 => -63,
    50252 => -63,
    50253 => -63,
    50254 => -63,
    50255 => -63,
    50256 => -63,
    50257 => -63,
    50258 => -63,
    50259 => -63,
    50260 => -63,
    50261 => -63,
    50262 => -63,
    50263 => -63,
    50264 => -63,
    50265 => -63,
    50266 => -63,
    50267 => -63,
    50268 => -63,
    50269 => -63,
    50270 => -63,
    50271 => -63,
    50272 => -63,
    50273 => -63,
    50274 => -63,
    50275 => -63,
    50276 => -63,
    50277 => -63,
    50278 => -63,
    50279 => -63,
    50280 => -63,
    50281 => -63,
    50282 => -63,
    50283 => -63,
    50284 => -63,
    50285 => -63,
    50286 => -63,
    50287 => -63,
    50288 => -63,
    50289 => -63,
    50290 => -63,
    50291 => -63,
    50292 => -63,
    50293 => -63,
    50294 => -63,
    50295 => -63,
    50296 => -63,
    50297 => -63,
    50298 => -63,
    50299 => -63,
    50300 => -63,
    50301 => -63,
    50302 => -63,
    50303 => -63,
    50304 => -63,
    50305 => -63,
    50306 => -63,
    50307 => -63,
    50308 => -63,
    50309 => -63,
    50310 => -63,
    50311 => -63,
    50312 => -63,
    50313 => -63,
    50314 => -63,
    50315 => -63,
    50316 => -63,
    50317 => -63,
    50318 => -63,
    50319 => -63,
    50320 => -63,
    50321 => -63,
    50322 => -63,
    50323 => -63,
    50324 => -63,
    50325 => -63,
    50326 => -63,
    50327 => -63,
    50328 => -63,
    50329 => -63,
    50330 => -63,
    50331 => -63,
    50332 => -63,
    50333 => -63,
    50334 => -63,
    50335 => -63,
    50336 => -63,
    50337 => -63,
    50338 => -63,
    50339 => -63,
    50340 => -63,
    50341 => -63,
    50342 => -63,
    50343 => -63,
    50344 => -63,
    50345 => -63,
    50346 => -63,
    50347 => -63,
    50348 => -63,
    50349 => -63,
    50350 => -63,
    50351 => -63,
    50352 => -63,
    50353 => -63,
    50354 => -63,
    50355 => -63,
    50356 => -63,
    50357 => -63,
    50358 => -63,
    50359 => -63,
    50360 => -63,
    50361 => -63,
    50362 => -63,
    50363 => -63,
    50364 => -63,
    50365 => -63,
    50366 => -63,
    50367 => -63,
    50368 => -63,
    50369 => -63,
    50370 => -63,
    50371 => -63,
    50372 => -63,
    50373 => -63,
    50374 => -63,
    50375 => -63,
    50376 => -63,
    50377 => -63,
    50378 => -63,
    50379 => -63,
    50380 => -63,
    50381 => -63,
    50382 => -63,
    50383 => -63,
    50384 => -63,
    50385 => -63,
    50386 => -63,
    50387 => -63,
    50388 => -63,
    50389 => -63,
    50390 => -63,
    50391 => -63,
    50392 => -63,
    50393 => -63,
    50394 => -63,
    50395 => -63,
    50396 => -63,
    50397 => -63,
    50398 => -63,
    50399 => -63,
    50400 => -63,
    50401 => -63,
    50402 => -63,
    50403 => -63,
    50404 => -63,
    50405 => -63,
    50406 => -63,
    50407 => -63,
    50408 => -63,
    50409 => -63,
    50410 => -63,
    50411 => -63,
    50412 => -63,
    50413 => -63,
    50414 => -63,
    50415 => -63,
    50416 => -63,
    50417 => -63,
    50418 => -63,
    50419 => -63,
    50420 => -63,
    50421 => -63,
    50422 => -63,
    50423 => -63,
    50424 => -63,
    50425 => -63,
    50426 => -63,
    50427 => -63,
    50428 => -63,
    50429 => -63,
    50430 => -63,
    50431 => -63,
    50432 => -63,
    50433 => -63,
    50434 => -63,
    50435 => -63,
    50436 => -63,
    50437 => -63,
    50438 => -63,
    50439 => -63,
    50440 => -63,
    50441 => -63,
    50442 => -63,
    50443 => -63,
    50444 => -63,
    50445 => -63,
    50446 => -63,
    50447 => -63,
    50448 => -63,
    50449 => -63,
    50450 => -63,
    50451 => -63,
    50452 => -63,
    50453 => -63,
    50454 => -63,
    50455 => -63,
    50456 => -63,
    50457 => -63,
    50458 => -63,
    50459 => -63,
    50460 => -63,
    50461 => -63,
    50462 => -63,
    50463 => -63,
    50464 => -63,
    50465 => -63,
    50466 => -63,
    50467 => -62,
    50468 => -62,
    50469 => -62,
    50470 => -62,
    50471 => -62,
    50472 => -62,
    50473 => -62,
    50474 => -62,
    50475 => -62,
    50476 => -62,
    50477 => -62,
    50478 => -62,
    50479 => -62,
    50480 => -62,
    50481 => -62,
    50482 => -62,
    50483 => -62,
    50484 => -62,
    50485 => -62,
    50486 => -62,
    50487 => -62,
    50488 => -62,
    50489 => -62,
    50490 => -62,
    50491 => -62,
    50492 => -62,
    50493 => -62,
    50494 => -62,
    50495 => -62,
    50496 => -62,
    50497 => -62,
    50498 => -62,
    50499 => -62,
    50500 => -62,
    50501 => -62,
    50502 => -62,
    50503 => -62,
    50504 => -62,
    50505 => -62,
    50506 => -62,
    50507 => -62,
    50508 => -62,
    50509 => -62,
    50510 => -62,
    50511 => -62,
    50512 => -62,
    50513 => -62,
    50514 => -62,
    50515 => -62,
    50516 => -62,
    50517 => -62,
    50518 => -62,
    50519 => -62,
    50520 => -62,
    50521 => -62,
    50522 => -62,
    50523 => -62,
    50524 => -62,
    50525 => -62,
    50526 => -62,
    50527 => -62,
    50528 => -62,
    50529 => -62,
    50530 => -62,
    50531 => -62,
    50532 => -62,
    50533 => -62,
    50534 => -62,
    50535 => -62,
    50536 => -62,
    50537 => -62,
    50538 => -62,
    50539 => -62,
    50540 => -62,
    50541 => -62,
    50542 => -62,
    50543 => -62,
    50544 => -62,
    50545 => -62,
    50546 => -62,
    50547 => -62,
    50548 => -62,
    50549 => -62,
    50550 => -62,
    50551 => -62,
    50552 => -62,
    50553 => -62,
    50554 => -62,
    50555 => -62,
    50556 => -62,
    50557 => -62,
    50558 => -62,
    50559 => -62,
    50560 => -62,
    50561 => -62,
    50562 => -62,
    50563 => -62,
    50564 => -62,
    50565 => -62,
    50566 => -62,
    50567 => -62,
    50568 => -62,
    50569 => -62,
    50570 => -62,
    50571 => -62,
    50572 => -62,
    50573 => -62,
    50574 => -62,
    50575 => -62,
    50576 => -62,
    50577 => -62,
    50578 => -62,
    50579 => -62,
    50580 => -62,
    50581 => -62,
    50582 => -62,
    50583 => -62,
    50584 => -62,
    50585 => -62,
    50586 => -62,
    50587 => -62,
    50588 => -62,
    50589 => -62,
    50590 => -62,
    50591 => -62,
    50592 => -62,
    50593 => -62,
    50594 => -62,
    50595 => -62,
    50596 => -62,
    50597 => -62,
    50598 => -62,
    50599 => -62,
    50600 => -62,
    50601 => -62,
    50602 => -62,
    50603 => -62,
    50604 => -62,
    50605 => -62,
    50606 => -62,
    50607 => -62,
    50608 => -62,
    50609 => -62,
    50610 => -62,
    50611 => -62,
    50612 => -62,
    50613 => -62,
    50614 => -62,
    50615 => -62,
    50616 => -62,
    50617 => -62,
    50618 => -62,
    50619 => -62,
    50620 => -62,
    50621 => -62,
    50622 => -62,
    50623 => -62,
    50624 => -62,
    50625 => -62,
    50626 => -62,
    50627 => -62,
    50628 => -62,
    50629 => -62,
    50630 => -62,
    50631 => -62,
    50632 => -62,
    50633 => -62,
    50634 => -62,
    50635 => -62,
    50636 => -62,
    50637 => -62,
    50638 => -62,
    50639 => -62,
    50640 => -62,
    50641 => -62,
    50642 => -62,
    50643 => -62,
    50644 => -62,
    50645 => -62,
    50646 => -62,
    50647 => -62,
    50648 => -62,
    50649 => -62,
    50650 => -62,
    50651 => -62,
    50652 => -62,
    50653 => -62,
    50654 => -62,
    50655 => -62,
    50656 => -62,
    50657 => -62,
    50658 => -62,
    50659 => -62,
    50660 => -62,
    50661 => -62,
    50662 => -62,
    50663 => -62,
    50664 => -62,
    50665 => -62,
    50666 => -62,
    50667 => -62,
    50668 => -62,
    50669 => -62,
    50670 => -62,
    50671 => -62,
    50672 => -62,
    50673 => -62,
    50674 => -62,
    50675 => -62,
    50676 => -62,
    50677 => -62,
    50678 => -62,
    50679 => -62,
    50680 => -62,
    50681 => -62,
    50682 => -62,
    50683 => -62,
    50684 => -62,
    50685 => -62,
    50686 => -62,
    50687 => -62,
    50688 => -62,
    50689 => -62,
    50690 => -62,
    50691 => -62,
    50692 => -62,
    50693 => -62,
    50694 => -62,
    50695 => -62,
    50696 => -62,
    50697 => -62,
    50698 => -62,
    50699 => -62,
    50700 => -62,
    50701 => -62,
    50702 => -62,
    50703 => -62,
    50704 => -62,
    50705 => -62,
    50706 => -62,
    50707 => -62,
    50708 => -62,
    50709 => -62,
    50710 => -62,
    50711 => -62,
    50712 => -62,
    50713 => -62,
    50714 => -62,
    50715 => -62,
    50716 => -62,
    50717 => -62,
    50718 => -62,
    50719 => -62,
    50720 => -62,
    50721 => -62,
    50722 => -62,
    50723 => -62,
    50724 => -62,
    50725 => -62,
    50726 => -62,
    50727 => -62,
    50728 => -62,
    50729 => -62,
    50730 => -62,
    50731 => -62,
    50732 => -62,
    50733 => -62,
    50734 => -62,
    50735 => -62,
    50736 => -62,
    50737 => -62,
    50738 => -62,
    50739 => -62,
    50740 => -62,
    50741 => -62,
    50742 => -62,
    50743 => -62,
    50744 => -62,
    50745 => -62,
    50746 => -62,
    50747 => -62,
    50748 => -62,
    50749 => -62,
    50750 => -62,
    50751 => -62,
    50752 => -62,
    50753 => -62,
    50754 => -62,
    50755 => -62,
    50756 => -62,
    50757 => -62,
    50758 => -62,
    50759 => -62,
    50760 => -62,
    50761 => -62,
    50762 => -62,
    50763 => -62,
    50764 => -62,
    50765 => -62,
    50766 => -62,
    50767 => -62,
    50768 => -62,
    50769 => -62,
    50770 => -62,
    50771 => -62,
    50772 => -62,
    50773 => -62,
    50774 => -62,
    50775 => -62,
    50776 => -62,
    50777 => -62,
    50778 => -62,
    50779 => -62,
    50780 => -62,
    50781 => -62,
    50782 => -62,
    50783 => -62,
    50784 => -62,
    50785 => -62,
    50786 => -62,
    50787 => -62,
    50788 => -62,
    50789 => -62,
    50790 => -62,
    50791 => -62,
    50792 => -62,
    50793 => -62,
    50794 => -62,
    50795 => -62,
    50796 => -62,
    50797 => -62,
    50798 => -62,
    50799 => -62,
    50800 => -62,
    50801 => -62,
    50802 => -62,
    50803 => -62,
    50804 => -62,
    50805 => -62,
    50806 => -62,
    50807 => -62,
    50808 => -62,
    50809 => -62,
    50810 => -62,
    50811 => -62,
    50812 => -62,
    50813 => -62,
    50814 => -62,
    50815 => -62,
    50816 => -62,
    50817 => -62,
    50818 => -62,
    50819 => -62,
    50820 => -62,
    50821 => -62,
    50822 => -62,
    50823 => -62,
    50824 => -62,
    50825 => -62,
    50826 => -62,
    50827 => -62,
    50828 => -62,
    50829 => -62,
    50830 => -62,
    50831 => -62,
    50832 => -62,
    50833 => -62,
    50834 => -62,
    50835 => -62,
    50836 => -62,
    50837 => -62,
    50838 => -62,
    50839 => -62,
    50840 => -62,
    50841 => -62,
    50842 => -62,
    50843 => -62,
    50844 => -62,
    50845 => -62,
    50846 => -62,
    50847 => -62,
    50848 => -62,
    50849 => -62,
    50850 => -62,
    50851 => -62,
    50852 => -62,
    50853 => -62,
    50854 => -62,
    50855 => -62,
    50856 => -62,
    50857 => -62,
    50858 => -62,
    50859 => -62,
    50860 => -62,
    50861 => -62,
    50862 => -62,
    50863 => -62,
    50864 => -62,
    50865 => -62,
    50866 => -62,
    50867 => -62,
    50868 => -62,
    50869 => -62,
    50870 => -62,
    50871 => -62,
    50872 => -62,
    50873 => -62,
    50874 => -62,
    50875 => -62,
    50876 => -62,
    50877 => -62,
    50878 => -62,
    50879 => -62,
    50880 => -62,
    50881 => -62,
    50882 => -62,
    50883 => -62,
    50884 => -62,
    50885 => -62,
    50886 => -62,
    50887 => -62,
    50888 => -62,
    50889 => -62,
    50890 => -62,
    50891 => -62,
    50892 => -62,
    50893 => -62,
    50894 => -62,
    50895 => -62,
    50896 => -62,
    50897 => -62,
    50898 => -62,
    50899 => -62,
    50900 => -62,
    50901 => -62,
    50902 => -62,
    50903 => -62,
    50904 => -62,
    50905 => -62,
    50906 => -62,
    50907 => -62,
    50908 => -62,
    50909 => -62,
    50910 => -62,
    50911 => -62,
    50912 => -62,
    50913 => -62,
    50914 => -62,
    50915 => -62,
    50916 => -62,
    50917 => -62,
    50918 => -62,
    50919 => -62,
    50920 => -62,
    50921 => -62,
    50922 => -62,
    50923 => -62,
    50924 => -62,
    50925 => -62,
    50926 => -62,
    50927 => -62,
    50928 => -62,
    50929 => -62,
    50930 => -62,
    50931 => -62,
    50932 => -62,
    50933 => -62,
    50934 => -62,
    50935 => -62,
    50936 => -62,
    50937 => -62,
    50938 => -62,
    50939 => -62,
    50940 => -62,
    50941 => -62,
    50942 => -62,
    50943 => -62,
    50944 => -62,
    50945 => -62,
    50946 => -62,
    50947 => -62,
    50948 => -62,
    50949 => -62,
    50950 => -62,
    50951 => -62,
    50952 => -62,
    50953 => -62,
    50954 => -62,
    50955 => -62,
    50956 => -62,
    50957 => -62,
    50958 => -62,
    50959 => -62,
    50960 => -62,
    50961 => -62,
    50962 => -62,
    50963 => -62,
    50964 => -62,
    50965 => -62,
    50966 => -62,
    50967 => -62,
    50968 => -62,
    50969 => -62,
    50970 => -62,
    50971 => -62,
    50972 => -62,
    50973 => -62,
    50974 => -62,
    50975 => -62,
    50976 => -62,
    50977 => -62,
    50978 => -62,
    50979 => -62,
    50980 => -62,
    50981 => -62,
    50982 => -62,
    50983 => -62,
    50984 => -62,
    50985 => -62,
    50986 => -62,
    50987 => -62,
    50988 => -62,
    50989 => -62,
    50990 => -62,
    50991 => -62,
    50992 => -62,
    50993 => -62,
    50994 => -62,
    50995 => -62,
    50996 => -62,
    50997 => -62,
    50998 => -62,
    50999 => -62,
    51000 => -62,
    51001 => -62,
    51002 => -62,
    51003 => -62,
    51004 => -62,
    51005 => -62,
    51006 => -62,
    51007 => -62,
    51008 => -62,
    51009 => -62,
    51010 => -62,
    51011 => -62,
    51012 => -62,
    51013 => -62,
    51014 => -62,
    51015 => -62,
    51016 => -62,
    51017 => -62,
    51018 => -62,
    51019 => -62,
    51020 => -62,
    51021 => -62,
    51022 => -62,
    51023 => -62,
    51024 => -62,
    51025 => -62,
    51026 => -62,
    51027 => -62,
    51028 => -62,
    51029 => -62,
    51030 => -62,
    51031 => -62,
    51032 => -62,
    51033 => -62,
    51034 => -62,
    51035 => -62,
    51036 => -62,
    51037 => -62,
    51038 => -62,
    51039 => -62,
    51040 => -62,
    51041 => -62,
    51042 => -62,
    51043 => -62,
    51044 => -62,
    51045 => -62,
    51046 => -62,
    51047 => -62,
    51048 => -62,
    51049 => -62,
    51050 => -62,
    51051 => -62,
    51052 => -62,
    51053 => -62,
    51054 => -62,
    51055 => -62,
    51056 => -62,
    51057 => -62,
    51058 => -62,
    51059 => -62,
    51060 => -62,
    51061 => -62,
    51062 => -62,
    51063 => -62,
    51064 => -62,
    51065 => -62,
    51066 => -62,
    51067 => -62,
    51068 => -62,
    51069 => -62,
    51070 => -62,
    51071 => -62,
    51072 => -62,
    51073 => -62,
    51074 => -62,
    51075 => -62,
    51076 => -62,
    51077 => -62,
    51078 => -62,
    51079 => -62,
    51080 => -62,
    51081 => -62,
    51082 => -62,
    51083 => -62,
    51084 => -62,
    51085 => -62,
    51086 => -62,
    51087 => -62,
    51088 => -62,
    51089 => -62,
    51090 => -62,
    51091 => -62,
    51092 => -62,
    51093 => -62,
    51094 => -62,
    51095 => -62,
    51096 => -62,
    51097 => -62,
    51098 => -62,
    51099 => -62,
    51100 => -62,
    51101 => -62,
    51102 => -62,
    51103 => -62,
    51104 => -62,
    51105 => -62,
    51106 => -62,
    51107 => -62,
    51108 => -62,
    51109 => -62,
    51110 => -62,
    51111 => -62,
    51112 => -62,
    51113 => -62,
    51114 => -62,
    51115 => -62,
    51116 => -62,
    51117 => -62,
    51118 => -62,
    51119 => -62,
    51120 => -62,
    51121 => -62,
    51122 => -62,
    51123 => -62,
    51124 => -62,
    51125 => -62,
    51126 => -62,
    51127 => -62,
    51128 => -62,
    51129 => -62,
    51130 => -62,
    51131 => -62,
    51132 => -62,
    51133 => -62,
    51134 => -62,
    51135 => -62,
    51136 => -62,
    51137 => -62,
    51138 => -62,
    51139 => -62,
    51140 => -62,
    51141 => -62,
    51142 => -62,
    51143 => -62,
    51144 => -62,
    51145 => -62,
    51146 => -62,
    51147 => -62,
    51148 => -62,
    51149 => -62,
    51150 => -62,
    51151 => -62,
    51152 => -62,
    51153 => -62,
    51154 => -62,
    51155 => -62,
    51156 => -62,
    51157 => -62,
    51158 => -62,
    51159 => -62,
    51160 => -62,
    51161 => -62,
    51162 => -62,
    51163 => -62,
    51164 => -62,
    51165 => -62,
    51166 => -62,
    51167 => -62,
    51168 => -62,
    51169 => -62,
    51170 => -62,
    51171 => -62,
    51172 => -62,
    51173 => -62,
    51174 => -62,
    51175 => -62,
    51176 => -62,
    51177 => -62,
    51178 => -62,
    51179 => -62,
    51180 => -62,
    51181 => -62,
    51182 => -62,
    51183 => -62,
    51184 => -62,
    51185 => -62,
    51186 => -62,
    51187 => -62,
    51188 => -62,
    51189 => -62,
    51190 => -62,
    51191 => -62,
    51192 => -62,
    51193 => -62,
    51194 => -62,
    51195 => -62,
    51196 => -62,
    51197 => -62,
    51198 => -62,
    51199 => -62,
    51200 => -62,
    51201 => -62,
    51202 => -62,
    51203 => -62,
    51204 => -62,
    51205 => -62,
    51206 => -62,
    51207 => -62,
    51208 => -62,
    51209 => -62,
    51210 => -62,
    51211 => -62,
    51212 => -62,
    51213 => -62,
    51214 => -62,
    51215 => -62,
    51216 => -62,
    51217 => -62,
    51218 => -62,
    51219 => -62,
    51220 => -62,
    51221 => -62,
    51222 => -62,
    51223 => -62,
    51224 => -62,
    51225 => -62,
    51226 => -62,
    51227 => -62,
    51228 => -62,
    51229 => -62,
    51230 => -62,
    51231 => -62,
    51232 => -62,
    51233 => -62,
    51234 => -62,
    51235 => -62,
    51236 => -62,
    51237 => -62,
    51238 => -62,
    51239 => -62,
    51240 => -62,
    51241 => -62,
    51242 => -62,
    51243 => -62,
    51244 => -62,
    51245 => -62,
    51246 => -62,
    51247 => -62,
    51248 => -62,
    51249 => -62,
    51250 => -62,
    51251 => -62,
    51252 => -62,
    51253 => -62,
    51254 => -62,
    51255 => -62,
    51256 => -62,
    51257 => -62,
    51258 => -62,
    51259 => -62,
    51260 => -62,
    51261 => -62,
    51262 => -62,
    51263 => -62,
    51264 => -62,
    51265 => -62,
    51266 => -62,
    51267 => -62,
    51268 => -62,
    51269 => -62,
    51270 => -62,
    51271 => -62,
    51272 => -62,
    51273 => -62,
    51274 => -62,
    51275 => -62,
    51276 => -62,
    51277 => -62,
    51278 => -62,
    51279 => -62,
    51280 => -62,
    51281 => -62,
    51282 => -62,
    51283 => -62,
    51284 => -62,
    51285 => -62,
    51286 => -62,
    51287 => -62,
    51288 => -62,
    51289 => -62,
    51290 => -62,
    51291 => -62,
    51292 => -62,
    51293 => -62,
    51294 => -62,
    51295 => -62,
    51296 => -62,
    51297 => -62,
    51298 => -62,
    51299 => -62,
    51300 => -62,
    51301 => -62,
    51302 => -62,
    51303 => -62,
    51304 => -62,
    51305 => -62,
    51306 => -62,
    51307 => -62,
    51308 => -62,
    51309 => -62,
    51310 => -62,
    51311 => -62,
    51312 => -62,
    51313 => -62,
    51314 => -62,
    51315 => -62,
    51316 => -62,
    51317 => -62,
    51318 => -62,
    51319 => -62,
    51320 => -62,
    51321 => -62,
    51322 => -62,
    51323 => -62,
    51324 => -62,
    51325 => -62,
    51326 => -62,
    51327 => -62,
    51328 => -62,
    51329 => -62,
    51330 => -62,
    51331 => -62,
    51332 => -62,
    51333 => -62,
    51334 => -62,
    51335 => -62,
    51336 => -62,
    51337 => -62,
    51338 => -62,
    51339 => -62,
    51340 => -62,
    51341 => -62,
    51342 => -62,
    51343 => -62,
    51344 => -62,
    51345 => -62,
    51346 => -62,
    51347 => -62,
    51348 => -62,
    51349 => -62,
    51350 => -62,
    51351 => -62,
    51352 => -62,
    51353 => -62,
    51354 => -62,
    51355 => -62,
    51356 => -62,
    51357 => -62,
    51358 => -62,
    51359 => -62,
    51360 => -62,
    51361 => -62,
    51362 => -62,
    51363 => -62,
    51364 => -62,
    51365 => -62,
    51366 => -62,
    51367 => -62,
    51368 => -62,
    51369 => -62,
    51370 => -62,
    51371 => -62,
    51372 => -62,
    51373 => -62,
    51374 => -62,
    51375 => -62,
    51376 => -62,
    51377 => -62,
    51378 => -62,
    51379 => -62,
    51380 => -62,
    51381 => -62,
    51382 => -62,
    51383 => -62,
    51384 => -62,
    51385 => -62,
    51386 => -62,
    51387 => -62,
    51388 => -62,
    51389 => -62,
    51390 => -62,
    51391 => -62,
    51392 => -62,
    51393 => -62,
    51394 => -62,
    51395 => -62,
    51396 => -62,
    51397 => -62,
    51398 => -62,
    51399 => -62,
    51400 => -62,
    51401 => -62,
    51402 => -62,
    51403 => -62,
    51404 => -62,
    51405 => -62,
    51406 => -62,
    51407 => -62,
    51408 => -62,
    51409 => -62,
    51410 => -62,
    51411 => -62,
    51412 => -62,
    51413 => -62,
    51414 => -62,
    51415 => -62,
    51416 => -62,
    51417 => -62,
    51418 => -62,
    51419 => -62,
    51420 => -62,
    51421 => -62,
    51422 => -62,
    51423 => -62,
    51424 => -62,
    51425 => -62,
    51426 => -62,
    51427 => -62,
    51428 => -62,
    51429 => -62,
    51430 => -62,
    51431 => -62,
    51432 => -62,
    51433 => -61,
    51434 => -61,
    51435 => -61,
    51436 => -61,
    51437 => -61,
    51438 => -61,
    51439 => -61,
    51440 => -61,
    51441 => -61,
    51442 => -61,
    51443 => -61,
    51444 => -61,
    51445 => -61,
    51446 => -61,
    51447 => -61,
    51448 => -61,
    51449 => -61,
    51450 => -61,
    51451 => -61,
    51452 => -61,
    51453 => -61,
    51454 => -61,
    51455 => -61,
    51456 => -61,
    51457 => -61,
    51458 => -61,
    51459 => -61,
    51460 => -61,
    51461 => -61,
    51462 => -61,
    51463 => -61,
    51464 => -61,
    51465 => -61,
    51466 => -61,
    51467 => -61,
    51468 => -61,
    51469 => -61,
    51470 => -61,
    51471 => -61,
    51472 => -61,
    51473 => -61,
    51474 => -61,
    51475 => -61,
    51476 => -61,
    51477 => -61,
    51478 => -61,
    51479 => -61,
    51480 => -61,
    51481 => -61,
    51482 => -61,
    51483 => -61,
    51484 => -61,
    51485 => -61,
    51486 => -61,
    51487 => -61,
    51488 => -61,
    51489 => -61,
    51490 => -61,
    51491 => -61,
    51492 => -61,
    51493 => -61,
    51494 => -61,
    51495 => -61,
    51496 => -61,
    51497 => -61,
    51498 => -61,
    51499 => -61,
    51500 => -61,
    51501 => -61,
    51502 => -61,
    51503 => -61,
    51504 => -61,
    51505 => -61,
    51506 => -61,
    51507 => -61,
    51508 => -61,
    51509 => -61,
    51510 => -61,
    51511 => -61,
    51512 => -61,
    51513 => -61,
    51514 => -61,
    51515 => -61,
    51516 => -61,
    51517 => -61,
    51518 => -61,
    51519 => -61,
    51520 => -61,
    51521 => -61,
    51522 => -61,
    51523 => -61,
    51524 => -61,
    51525 => -61,
    51526 => -61,
    51527 => -61,
    51528 => -61,
    51529 => -61,
    51530 => -61,
    51531 => -61,
    51532 => -61,
    51533 => -61,
    51534 => -61,
    51535 => -61,
    51536 => -61,
    51537 => -61,
    51538 => -61,
    51539 => -61,
    51540 => -61,
    51541 => -61,
    51542 => -61,
    51543 => -61,
    51544 => -61,
    51545 => -61,
    51546 => -61,
    51547 => -61,
    51548 => -61,
    51549 => -61,
    51550 => -61,
    51551 => -61,
    51552 => -61,
    51553 => -61,
    51554 => -61,
    51555 => -61,
    51556 => -61,
    51557 => -61,
    51558 => -61,
    51559 => -61,
    51560 => -61,
    51561 => -61,
    51562 => -61,
    51563 => -61,
    51564 => -61,
    51565 => -61,
    51566 => -61,
    51567 => -61,
    51568 => -61,
    51569 => -61,
    51570 => -61,
    51571 => -61,
    51572 => -61,
    51573 => -61,
    51574 => -61,
    51575 => -61,
    51576 => -61,
    51577 => -61,
    51578 => -61,
    51579 => -61,
    51580 => -61,
    51581 => -61,
    51582 => -61,
    51583 => -61,
    51584 => -61,
    51585 => -61,
    51586 => -61,
    51587 => -61,
    51588 => -61,
    51589 => -61,
    51590 => -61,
    51591 => -61,
    51592 => -61,
    51593 => -61,
    51594 => -61,
    51595 => -61,
    51596 => -61,
    51597 => -61,
    51598 => -61,
    51599 => -61,
    51600 => -61,
    51601 => -61,
    51602 => -61,
    51603 => -61,
    51604 => -61,
    51605 => -61,
    51606 => -61,
    51607 => -61,
    51608 => -61,
    51609 => -61,
    51610 => -61,
    51611 => -61,
    51612 => -61,
    51613 => -61,
    51614 => -61,
    51615 => -61,
    51616 => -61,
    51617 => -61,
    51618 => -61,
    51619 => -61,
    51620 => -61,
    51621 => -61,
    51622 => -61,
    51623 => -61,
    51624 => -61,
    51625 => -61,
    51626 => -61,
    51627 => -61,
    51628 => -61,
    51629 => -61,
    51630 => -61,
    51631 => -61,
    51632 => -61,
    51633 => -61,
    51634 => -61,
    51635 => -61,
    51636 => -61,
    51637 => -61,
    51638 => -61,
    51639 => -61,
    51640 => -61,
    51641 => -61,
    51642 => -61,
    51643 => -61,
    51644 => -61,
    51645 => -61,
    51646 => -61,
    51647 => -61,
    51648 => -61,
    51649 => -61,
    51650 => -61,
    51651 => -61,
    51652 => -61,
    51653 => -61,
    51654 => -61,
    51655 => -61,
    51656 => -61,
    51657 => -61,
    51658 => -61,
    51659 => -61,
    51660 => -61,
    51661 => -61,
    51662 => -61,
    51663 => -61,
    51664 => -61,
    51665 => -61,
    51666 => -61,
    51667 => -61,
    51668 => -61,
    51669 => -61,
    51670 => -61,
    51671 => -61,
    51672 => -61,
    51673 => -61,
    51674 => -61,
    51675 => -61,
    51676 => -61,
    51677 => -61,
    51678 => -61,
    51679 => -61,
    51680 => -61,
    51681 => -61,
    51682 => -61,
    51683 => -61,
    51684 => -61,
    51685 => -61,
    51686 => -61,
    51687 => -61,
    51688 => -61,
    51689 => -61,
    51690 => -61,
    51691 => -61,
    51692 => -61,
    51693 => -61,
    51694 => -61,
    51695 => -61,
    51696 => -61,
    51697 => -61,
    51698 => -61,
    51699 => -61,
    51700 => -61,
    51701 => -61,
    51702 => -61,
    51703 => -61,
    51704 => -61,
    51705 => -61,
    51706 => -61,
    51707 => -61,
    51708 => -61,
    51709 => -61,
    51710 => -61,
    51711 => -61,
    51712 => -61,
    51713 => -61,
    51714 => -61,
    51715 => -61,
    51716 => -61,
    51717 => -61,
    51718 => -61,
    51719 => -61,
    51720 => -61,
    51721 => -61,
    51722 => -61,
    51723 => -61,
    51724 => -61,
    51725 => -61,
    51726 => -61,
    51727 => -61,
    51728 => -61,
    51729 => -61,
    51730 => -61,
    51731 => -61,
    51732 => -61,
    51733 => -61,
    51734 => -61,
    51735 => -61,
    51736 => -61,
    51737 => -61,
    51738 => -61,
    51739 => -61,
    51740 => -61,
    51741 => -61,
    51742 => -61,
    51743 => -61,
    51744 => -61,
    51745 => -61,
    51746 => -61,
    51747 => -61,
    51748 => -61,
    51749 => -61,
    51750 => -61,
    51751 => -61,
    51752 => -61,
    51753 => -61,
    51754 => -61,
    51755 => -61,
    51756 => -61,
    51757 => -61,
    51758 => -61,
    51759 => -61,
    51760 => -61,
    51761 => -61,
    51762 => -61,
    51763 => -61,
    51764 => -61,
    51765 => -61,
    51766 => -61,
    51767 => -61,
    51768 => -61,
    51769 => -61,
    51770 => -61,
    51771 => -61,
    51772 => -61,
    51773 => -61,
    51774 => -61,
    51775 => -61,
    51776 => -61,
    51777 => -61,
    51778 => -61,
    51779 => -61,
    51780 => -61,
    51781 => -61,
    51782 => -61,
    51783 => -61,
    51784 => -61,
    51785 => -61,
    51786 => -61,
    51787 => -61,
    51788 => -61,
    51789 => -61,
    51790 => -61,
    51791 => -61,
    51792 => -61,
    51793 => -61,
    51794 => -61,
    51795 => -61,
    51796 => -61,
    51797 => -61,
    51798 => -61,
    51799 => -61,
    51800 => -61,
    51801 => -61,
    51802 => -61,
    51803 => -61,
    51804 => -61,
    51805 => -61,
    51806 => -61,
    51807 => -61,
    51808 => -61,
    51809 => -61,
    51810 => -61,
    51811 => -61,
    51812 => -61,
    51813 => -61,
    51814 => -61,
    51815 => -61,
    51816 => -61,
    51817 => -61,
    51818 => -61,
    51819 => -61,
    51820 => -61,
    51821 => -61,
    51822 => -61,
    51823 => -61,
    51824 => -61,
    51825 => -61,
    51826 => -61,
    51827 => -61,
    51828 => -61,
    51829 => -61,
    51830 => -61,
    51831 => -61,
    51832 => -61,
    51833 => -61,
    51834 => -61,
    51835 => -61,
    51836 => -61,
    51837 => -61,
    51838 => -61,
    51839 => -61,
    51840 => -61,
    51841 => -61,
    51842 => -61,
    51843 => -61,
    51844 => -61,
    51845 => -61,
    51846 => -61,
    51847 => -61,
    51848 => -61,
    51849 => -61,
    51850 => -61,
    51851 => -61,
    51852 => -61,
    51853 => -61,
    51854 => -61,
    51855 => -61,
    51856 => -61,
    51857 => -61,
    51858 => -61,
    51859 => -61,
    51860 => -61,
    51861 => -61,
    51862 => -61,
    51863 => -61,
    51864 => -61,
    51865 => -61,
    51866 => -61,
    51867 => -61,
    51868 => -61,
    51869 => -61,
    51870 => -61,
    51871 => -61,
    51872 => -61,
    51873 => -61,
    51874 => -61,
    51875 => -61,
    51876 => -61,
    51877 => -61,
    51878 => -61,
    51879 => -61,
    51880 => -61,
    51881 => -61,
    51882 => -61,
    51883 => -61,
    51884 => -61,
    51885 => -61,
    51886 => -61,
    51887 => -61,
    51888 => -61,
    51889 => -61,
    51890 => -61,
    51891 => -61,
    51892 => -61,
    51893 => -61,
    51894 => -61,
    51895 => -61,
    51896 => -61,
    51897 => -61,
    51898 => -61,
    51899 => -61,
    51900 => -61,
    51901 => -61,
    51902 => -61,
    51903 => -61,
    51904 => -61,
    51905 => -61,
    51906 => -61,
    51907 => -61,
    51908 => -61,
    51909 => -61,
    51910 => -61,
    51911 => -61,
    51912 => -61,
    51913 => -61,
    51914 => -61,
    51915 => -61,
    51916 => -61,
    51917 => -61,
    51918 => -61,
    51919 => -61,
    51920 => -61,
    51921 => -61,
    51922 => -61,
    51923 => -61,
    51924 => -61,
    51925 => -61,
    51926 => -61,
    51927 => -61,
    51928 => -61,
    51929 => -61,
    51930 => -61,
    51931 => -61,
    51932 => -61,
    51933 => -61,
    51934 => -61,
    51935 => -61,
    51936 => -61,
    51937 => -61,
    51938 => -61,
    51939 => -61,
    51940 => -61,
    51941 => -61,
    51942 => -61,
    51943 => -61,
    51944 => -61,
    51945 => -61,
    51946 => -61,
    51947 => -61,
    51948 => -61,
    51949 => -61,
    51950 => -61,
    51951 => -61,
    51952 => -61,
    51953 => -61,
    51954 => -61,
    51955 => -61,
    51956 => -61,
    51957 => -61,
    51958 => -61,
    51959 => -61,
    51960 => -61,
    51961 => -61,
    51962 => -61,
    51963 => -61,
    51964 => -61,
    51965 => -61,
    51966 => -61,
    51967 => -61,
    51968 => -61,
    51969 => -61,
    51970 => -61,
    51971 => -61,
    51972 => -61,
    51973 => -61,
    51974 => -61,
    51975 => -61,
    51976 => -61,
    51977 => -61,
    51978 => -61,
    51979 => -61,
    51980 => -61,
    51981 => -61,
    51982 => -61,
    51983 => -61,
    51984 => -61,
    51985 => -61,
    51986 => -61,
    51987 => -61,
    51988 => -61,
    51989 => -61,
    51990 => -61,
    51991 => -61,
    51992 => -61,
    51993 => -61,
    51994 => -61,
    51995 => -61,
    51996 => -61,
    51997 => -61,
    51998 => -61,
    51999 => -61,
    52000 => -61,
    52001 => -61,
    52002 => -61,
    52003 => -61,
    52004 => -61,
    52005 => -61,
    52006 => -61,
    52007 => -61,
    52008 => -61,
    52009 => -61,
    52010 => -61,
    52011 => -61,
    52012 => -61,
    52013 => -61,
    52014 => -61,
    52015 => -61,
    52016 => -61,
    52017 => -61,
    52018 => -61,
    52019 => -61,
    52020 => -61,
    52021 => -61,
    52022 => -61,
    52023 => -61,
    52024 => -61,
    52025 => -61,
    52026 => -61,
    52027 => -61,
    52028 => -61,
    52029 => -61,
    52030 => -61,
    52031 => -61,
    52032 => -61,
    52033 => -61,
    52034 => -61,
    52035 => -61,
    52036 => -61,
    52037 => -61,
    52038 => -61,
    52039 => -61,
    52040 => -61,
    52041 => -61,
    52042 => -61,
    52043 => -61,
    52044 => -61,
    52045 => -61,
    52046 => -61,
    52047 => -61,
    52048 => -61,
    52049 => -61,
    52050 => -61,
    52051 => -61,
    52052 => -61,
    52053 => -61,
    52054 => -61,
    52055 => -61,
    52056 => -61,
    52057 => -61,
    52058 => -61,
    52059 => -61,
    52060 => -61,
    52061 => -61,
    52062 => -61,
    52063 => -61,
    52064 => -61,
    52065 => -61,
    52066 => -61,
    52067 => -61,
    52068 => -61,
    52069 => -61,
    52070 => -61,
    52071 => -61,
    52072 => -61,
    52073 => -61,
    52074 => -61,
    52075 => -61,
    52076 => -61,
    52077 => -61,
    52078 => -61,
    52079 => -61,
    52080 => -61,
    52081 => -61,
    52082 => -61,
    52083 => -61,
    52084 => -61,
    52085 => -61,
    52086 => -61,
    52087 => -61,
    52088 => -61,
    52089 => -61,
    52090 => -61,
    52091 => -61,
    52092 => -61,
    52093 => -61,
    52094 => -61,
    52095 => -61,
    52096 => -61,
    52097 => -61,
    52098 => -61,
    52099 => -61,
    52100 => -61,
    52101 => -60,
    52102 => -60,
    52103 => -60,
    52104 => -60,
    52105 => -60,
    52106 => -60,
    52107 => -60,
    52108 => -60,
    52109 => -60,
    52110 => -60,
    52111 => -60,
    52112 => -60,
    52113 => -60,
    52114 => -60,
    52115 => -60,
    52116 => -60,
    52117 => -60,
    52118 => -60,
    52119 => -60,
    52120 => -60,
    52121 => -60,
    52122 => -60,
    52123 => -60,
    52124 => -60,
    52125 => -60,
    52126 => -60,
    52127 => -60,
    52128 => -60,
    52129 => -60,
    52130 => -60,
    52131 => -60,
    52132 => -60,
    52133 => -60,
    52134 => -60,
    52135 => -60,
    52136 => -60,
    52137 => -60,
    52138 => -60,
    52139 => -60,
    52140 => -60,
    52141 => -60,
    52142 => -60,
    52143 => -60,
    52144 => -60,
    52145 => -60,
    52146 => -60,
    52147 => -60,
    52148 => -60,
    52149 => -60,
    52150 => -60,
    52151 => -60,
    52152 => -60,
    52153 => -60,
    52154 => -60,
    52155 => -60,
    52156 => -60,
    52157 => -60,
    52158 => -60,
    52159 => -60,
    52160 => -60,
    52161 => -60,
    52162 => -60,
    52163 => -60,
    52164 => -60,
    52165 => -60,
    52166 => -60,
    52167 => -60,
    52168 => -60,
    52169 => -60,
    52170 => -60,
    52171 => -60,
    52172 => -60,
    52173 => -60,
    52174 => -60,
    52175 => -60,
    52176 => -60,
    52177 => -60,
    52178 => -60,
    52179 => -60,
    52180 => -60,
    52181 => -60,
    52182 => -60,
    52183 => -60,
    52184 => -60,
    52185 => -60,
    52186 => -60,
    52187 => -60,
    52188 => -60,
    52189 => -60,
    52190 => -60,
    52191 => -60,
    52192 => -60,
    52193 => -60,
    52194 => -60,
    52195 => -60,
    52196 => -60,
    52197 => -60,
    52198 => -60,
    52199 => -60,
    52200 => -60,
    52201 => -60,
    52202 => -60,
    52203 => -60,
    52204 => -60,
    52205 => -60,
    52206 => -60,
    52207 => -60,
    52208 => -60,
    52209 => -60,
    52210 => -60,
    52211 => -60,
    52212 => -60,
    52213 => -60,
    52214 => -60,
    52215 => -60,
    52216 => -60,
    52217 => -60,
    52218 => -60,
    52219 => -60,
    52220 => -60,
    52221 => -60,
    52222 => -60,
    52223 => -60,
    52224 => -60,
    52225 => -60,
    52226 => -60,
    52227 => -60,
    52228 => -60,
    52229 => -60,
    52230 => -60,
    52231 => -60,
    52232 => -60,
    52233 => -60,
    52234 => -60,
    52235 => -60,
    52236 => -60,
    52237 => -60,
    52238 => -60,
    52239 => -60,
    52240 => -60,
    52241 => -60,
    52242 => -60,
    52243 => -60,
    52244 => -60,
    52245 => -60,
    52246 => -60,
    52247 => -60,
    52248 => -60,
    52249 => -60,
    52250 => -60,
    52251 => -60,
    52252 => -60,
    52253 => -60,
    52254 => -60,
    52255 => -60,
    52256 => -60,
    52257 => -60,
    52258 => -60,
    52259 => -60,
    52260 => -60,
    52261 => -60,
    52262 => -60,
    52263 => -60,
    52264 => -60,
    52265 => -60,
    52266 => -60,
    52267 => -60,
    52268 => -60,
    52269 => -60,
    52270 => -60,
    52271 => -60,
    52272 => -60,
    52273 => -60,
    52274 => -60,
    52275 => -60,
    52276 => -60,
    52277 => -60,
    52278 => -60,
    52279 => -60,
    52280 => -60,
    52281 => -60,
    52282 => -60,
    52283 => -60,
    52284 => -60,
    52285 => -60,
    52286 => -60,
    52287 => -60,
    52288 => -60,
    52289 => -60,
    52290 => -60,
    52291 => -60,
    52292 => -60,
    52293 => -60,
    52294 => -60,
    52295 => -60,
    52296 => -60,
    52297 => -60,
    52298 => -60,
    52299 => -60,
    52300 => -60,
    52301 => -60,
    52302 => -60,
    52303 => -60,
    52304 => -60,
    52305 => -60,
    52306 => -60,
    52307 => -60,
    52308 => -60,
    52309 => -60,
    52310 => -60,
    52311 => -60,
    52312 => -60,
    52313 => -60,
    52314 => -60,
    52315 => -60,
    52316 => -60,
    52317 => -60,
    52318 => -60,
    52319 => -60,
    52320 => -60,
    52321 => -60,
    52322 => -60,
    52323 => -60,
    52324 => -60,
    52325 => -60,
    52326 => -60,
    52327 => -60,
    52328 => -60,
    52329 => -60,
    52330 => -60,
    52331 => -60,
    52332 => -60,
    52333 => -60,
    52334 => -60,
    52335 => -60,
    52336 => -60,
    52337 => -60,
    52338 => -60,
    52339 => -60,
    52340 => -60,
    52341 => -60,
    52342 => -60,
    52343 => -60,
    52344 => -60,
    52345 => -60,
    52346 => -60,
    52347 => -60,
    52348 => -60,
    52349 => -60,
    52350 => -60,
    52351 => -60,
    52352 => -60,
    52353 => -60,
    52354 => -60,
    52355 => -60,
    52356 => -60,
    52357 => -60,
    52358 => -60,
    52359 => -60,
    52360 => -60,
    52361 => -60,
    52362 => -60,
    52363 => -60,
    52364 => -60,
    52365 => -60,
    52366 => -60,
    52367 => -60,
    52368 => -60,
    52369 => -60,
    52370 => -60,
    52371 => -60,
    52372 => -60,
    52373 => -60,
    52374 => -60,
    52375 => -60,
    52376 => -60,
    52377 => -60,
    52378 => -60,
    52379 => -60,
    52380 => -60,
    52381 => -60,
    52382 => -60,
    52383 => -60,
    52384 => -60,
    52385 => -60,
    52386 => -60,
    52387 => -60,
    52388 => -60,
    52389 => -60,
    52390 => -60,
    52391 => -60,
    52392 => -60,
    52393 => -60,
    52394 => -60,
    52395 => -60,
    52396 => -60,
    52397 => -60,
    52398 => -60,
    52399 => -60,
    52400 => -60,
    52401 => -60,
    52402 => -60,
    52403 => -60,
    52404 => -60,
    52405 => -60,
    52406 => -60,
    52407 => -60,
    52408 => -60,
    52409 => -60,
    52410 => -60,
    52411 => -60,
    52412 => -60,
    52413 => -60,
    52414 => -60,
    52415 => -60,
    52416 => -60,
    52417 => -60,
    52418 => -60,
    52419 => -60,
    52420 => -60,
    52421 => -60,
    52422 => -60,
    52423 => -60,
    52424 => -60,
    52425 => -60,
    52426 => -60,
    52427 => -60,
    52428 => -60,
    52429 => -60,
    52430 => -60,
    52431 => -60,
    52432 => -60,
    52433 => -60,
    52434 => -60,
    52435 => -60,
    52436 => -60,
    52437 => -60,
    52438 => -60,
    52439 => -60,
    52440 => -60,
    52441 => -60,
    52442 => -60,
    52443 => -60,
    52444 => -60,
    52445 => -60,
    52446 => -60,
    52447 => -60,
    52448 => -60,
    52449 => -60,
    52450 => -60,
    52451 => -60,
    52452 => -60,
    52453 => -60,
    52454 => -60,
    52455 => -60,
    52456 => -60,
    52457 => -60,
    52458 => -60,
    52459 => -60,
    52460 => -60,
    52461 => -60,
    52462 => -60,
    52463 => -60,
    52464 => -60,
    52465 => -60,
    52466 => -60,
    52467 => -60,
    52468 => -60,
    52469 => -60,
    52470 => -60,
    52471 => -60,
    52472 => -60,
    52473 => -60,
    52474 => -60,
    52475 => -60,
    52476 => -60,
    52477 => -60,
    52478 => -60,
    52479 => -60,
    52480 => -60,
    52481 => -60,
    52482 => -60,
    52483 => -60,
    52484 => -60,
    52485 => -60,
    52486 => -60,
    52487 => -60,
    52488 => -60,
    52489 => -60,
    52490 => -60,
    52491 => -60,
    52492 => -60,
    52493 => -60,
    52494 => -60,
    52495 => -60,
    52496 => -60,
    52497 => -60,
    52498 => -60,
    52499 => -60,
    52500 => -60,
    52501 => -60,
    52502 => -60,
    52503 => -60,
    52504 => -60,
    52505 => -60,
    52506 => -60,
    52507 => -60,
    52508 => -60,
    52509 => -60,
    52510 => -60,
    52511 => -60,
    52512 => -60,
    52513 => -60,
    52514 => -60,
    52515 => -60,
    52516 => -60,
    52517 => -60,
    52518 => -60,
    52519 => -60,
    52520 => -60,
    52521 => -60,
    52522 => -60,
    52523 => -60,
    52524 => -60,
    52525 => -60,
    52526 => -60,
    52527 => -60,
    52528 => -60,
    52529 => -60,
    52530 => -60,
    52531 => -60,
    52532 => -60,
    52533 => -60,
    52534 => -60,
    52535 => -60,
    52536 => -60,
    52537 => -60,
    52538 => -60,
    52539 => -60,
    52540 => -60,
    52541 => -60,
    52542 => -60,
    52543 => -60,
    52544 => -60,
    52545 => -60,
    52546 => -60,
    52547 => -60,
    52548 => -60,
    52549 => -60,
    52550 => -60,
    52551 => -60,
    52552 => -60,
    52553 => -60,
    52554 => -60,
    52555 => -60,
    52556 => -60,
    52557 => -60,
    52558 => -60,
    52559 => -60,
    52560 => -60,
    52561 => -60,
    52562 => -60,
    52563 => -60,
    52564 => -60,
    52565 => -60,
    52566 => -60,
    52567 => -60,
    52568 => -60,
    52569 => -60,
    52570 => -60,
    52571 => -60,
    52572 => -60,
    52573 => -60,
    52574 => -60,
    52575 => -60,
    52576 => -60,
    52577 => -60,
    52578 => -60,
    52579 => -60,
    52580 => -60,
    52581 => -60,
    52582 => -60,
    52583 => -60,
    52584 => -60,
    52585 => -60,
    52586 => -60,
    52587 => -60,
    52588 => -60,
    52589 => -60,
    52590 => -60,
    52591 => -60,
    52592 => -60,
    52593 => -60,
    52594 => -60,
    52595 => -60,
    52596 => -60,
    52597 => -60,
    52598 => -60,
    52599 => -60,
    52600 => -60,
    52601 => -60,
    52602 => -60,
    52603 => -60,
    52604 => -60,
    52605 => -60,
    52606 => -60,
    52607 => -60,
    52608 => -60,
    52609 => -60,
    52610 => -60,
    52611 => -60,
    52612 => -60,
    52613 => -60,
    52614 => -60,
    52615 => -60,
    52616 => -60,
    52617 => -60,
    52618 => -60,
    52619 => -60,
    52620 => -60,
    52621 => -60,
    52622 => -60,
    52623 => -60,
    52624 => -60,
    52625 => -60,
    52626 => -60,
    52627 => -60,
    52628 => -60,
    52629 => -60,
    52630 => -60,
    52631 => -60,
    52632 => -60,
    52633 => -60,
    52634 => -60,
    52635 => -60,
    52636 => -60,
    52637 => -60,
    52638 => -60,
    52639 => -60,
    52640 => -60,
    52641 => -60,
    52642 => -60,
    52643 => -60,
    52644 => -60,
    52645 => -60,
    52646 => -59,
    52647 => -59,
    52648 => -59,
    52649 => -59,
    52650 => -59,
    52651 => -59,
    52652 => -59,
    52653 => -59,
    52654 => -59,
    52655 => -59,
    52656 => -59,
    52657 => -59,
    52658 => -59,
    52659 => -59,
    52660 => -59,
    52661 => -59,
    52662 => -59,
    52663 => -59,
    52664 => -59,
    52665 => -59,
    52666 => -59,
    52667 => -59,
    52668 => -59,
    52669 => -59,
    52670 => -59,
    52671 => -59,
    52672 => -59,
    52673 => -59,
    52674 => -59,
    52675 => -59,
    52676 => -59,
    52677 => -59,
    52678 => -59,
    52679 => -59,
    52680 => -59,
    52681 => -59,
    52682 => -59,
    52683 => -59,
    52684 => -59,
    52685 => -59,
    52686 => -59,
    52687 => -59,
    52688 => -59,
    52689 => -59,
    52690 => -59,
    52691 => -59,
    52692 => -59,
    52693 => -59,
    52694 => -59,
    52695 => -59,
    52696 => -59,
    52697 => -59,
    52698 => -59,
    52699 => -59,
    52700 => -59,
    52701 => -59,
    52702 => -59,
    52703 => -59,
    52704 => -59,
    52705 => -59,
    52706 => -59,
    52707 => -59,
    52708 => -59,
    52709 => -59,
    52710 => -59,
    52711 => -59,
    52712 => -59,
    52713 => -59,
    52714 => -59,
    52715 => -59,
    52716 => -59,
    52717 => -59,
    52718 => -59,
    52719 => -59,
    52720 => -59,
    52721 => -59,
    52722 => -59,
    52723 => -59,
    52724 => -59,
    52725 => -59,
    52726 => -59,
    52727 => -59,
    52728 => -59,
    52729 => -59,
    52730 => -59,
    52731 => -59,
    52732 => -59,
    52733 => -59,
    52734 => -59,
    52735 => -59,
    52736 => -59,
    52737 => -59,
    52738 => -59,
    52739 => -59,
    52740 => -59,
    52741 => -59,
    52742 => -59,
    52743 => -59,
    52744 => -59,
    52745 => -59,
    52746 => -59,
    52747 => -59,
    52748 => -59,
    52749 => -59,
    52750 => -59,
    52751 => -59,
    52752 => -59,
    52753 => -59,
    52754 => -59,
    52755 => -59,
    52756 => -59,
    52757 => -59,
    52758 => -59,
    52759 => -59,
    52760 => -59,
    52761 => -59,
    52762 => -59,
    52763 => -59,
    52764 => -59,
    52765 => -59,
    52766 => -59,
    52767 => -59,
    52768 => -59,
    52769 => -59,
    52770 => -59,
    52771 => -59,
    52772 => -59,
    52773 => -59,
    52774 => -59,
    52775 => -59,
    52776 => -59,
    52777 => -59,
    52778 => -59,
    52779 => -59,
    52780 => -59,
    52781 => -59,
    52782 => -59,
    52783 => -59,
    52784 => -59,
    52785 => -59,
    52786 => -59,
    52787 => -59,
    52788 => -59,
    52789 => -59,
    52790 => -59,
    52791 => -59,
    52792 => -59,
    52793 => -59,
    52794 => -59,
    52795 => -59,
    52796 => -59,
    52797 => -59,
    52798 => -59,
    52799 => -59,
    52800 => -59,
    52801 => -59,
    52802 => -59,
    52803 => -59,
    52804 => -59,
    52805 => -59,
    52806 => -59,
    52807 => -59,
    52808 => -59,
    52809 => -59,
    52810 => -59,
    52811 => -59,
    52812 => -59,
    52813 => -59,
    52814 => -59,
    52815 => -59,
    52816 => -59,
    52817 => -59,
    52818 => -59,
    52819 => -59,
    52820 => -59,
    52821 => -59,
    52822 => -59,
    52823 => -59,
    52824 => -59,
    52825 => -59,
    52826 => -59,
    52827 => -59,
    52828 => -59,
    52829 => -59,
    52830 => -59,
    52831 => -59,
    52832 => -59,
    52833 => -59,
    52834 => -59,
    52835 => -59,
    52836 => -59,
    52837 => -59,
    52838 => -59,
    52839 => -59,
    52840 => -59,
    52841 => -59,
    52842 => -59,
    52843 => -59,
    52844 => -59,
    52845 => -59,
    52846 => -59,
    52847 => -59,
    52848 => -59,
    52849 => -59,
    52850 => -59,
    52851 => -59,
    52852 => -59,
    52853 => -59,
    52854 => -59,
    52855 => -59,
    52856 => -59,
    52857 => -59,
    52858 => -59,
    52859 => -59,
    52860 => -59,
    52861 => -59,
    52862 => -59,
    52863 => -59,
    52864 => -59,
    52865 => -59,
    52866 => -59,
    52867 => -59,
    52868 => -59,
    52869 => -59,
    52870 => -59,
    52871 => -59,
    52872 => -59,
    52873 => -59,
    52874 => -59,
    52875 => -59,
    52876 => -59,
    52877 => -59,
    52878 => -59,
    52879 => -59,
    52880 => -59,
    52881 => -59,
    52882 => -59,
    52883 => -59,
    52884 => -59,
    52885 => -59,
    52886 => -59,
    52887 => -59,
    52888 => -59,
    52889 => -59,
    52890 => -59,
    52891 => -59,
    52892 => -59,
    52893 => -59,
    52894 => -59,
    52895 => -59,
    52896 => -59,
    52897 => -59,
    52898 => -59,
    52899 => -59,
    52900 => -59,
    52901 => -59,
    52902 => -59,
    52903 => -59,
    52904 => -59,
    52905 => -59,
    52906 => -59,
    52907 => -59,
    52908 => -59,
    52909 => -59,
    52910 => -59,
    52911 => -59,
    52912 => -59,
    52913 => -59,
    52914 => -59,
    52915 => -59,
    52916 => -59,
    52917 => -59,
    52918 => -59,
    52919 => -59,
    52920 => -59,
    52921 => -59,
    52922 => -59,
    52923 => -59,
    52924 => -59,
    52925 => -59,
    52926 => -59,
    52927 => -59,
    52928 => -59,
    52929 => -59,
    52930 => -59,
    52931 => -59,
    52932 => -59,
    52933 => -59,
    52934 => -59,
    52935 => -59,
    52936 => -59,
    52937 => -59,
    52938 => -59,
    52939 => -59,
    52940 => -59,
    52941 => -59,
    52942 => -59,
    52943 => -59,
    52944 => -59,
    52945 => -59,
    52946 => -59,
    52947 => -59,
    52948 => -59,
    52949 => -59,
    52950 => -59,
    52951 => -59,
    52952 => -59,
    52953 => -59,
    52954 => -59,
    52955 => -59,
    52956 => -59,
    52957 => -59,
    52958 => -59,
    52959 => -59,
    52960 => -59,
    52961 => -59,
    52962 => -59,
    52963 => -59,
    52964 => -59,
    52965 => -59,
    52966 => -59,
    52967 => -59,
    52968 => -59,
    52969 => -59,
    52970 => -59,
    52971 => -59,
    52972 => -59,
    52973 => -59,
    52974 => -59,
    52975 => -59,
    52976 => -59,
    52977 => -59,
    52978 => -59,
    52979 => -59,
    52980 => -59,
    52981 => -59,
    52982 => -59,
    52983 => -59,
    52984 => -59,
    52985 => -59,
    52986 => -59,
    52987 => -59,
    52988 => -59,
    52989 => -59,
    52990 => -59,
    52991 => -59,
    52992 => -59,
    52993 => -59,
    52994 => -59,
    52995 => -59,
    52996 => -59,
    52997 => -59,
    52998 => -59,
    52999 => -59,
    53000 => -59,
    53001 => -59,
    53002 => -59,
    53003 => -59,
    53004 => -59,
    53005 => -59,
    53006 => -59,
    53007 => -59,
    53008 => -59,
    53009 => -59,
    53010 => -59,
    53011 => -59,
    53012 => -59,
    53013 => -59,
    53014 => -59,
    53015 => -59,
    53016 => -59,
    53017 => -59,
    53018 => -59,
    53019 => -59,
    53020 => -59,
    53021 => -59,
    53022 => -59,
    53023 => -59,
    53024 => -59,
    53025 => -59,
    53026 => -59,
    53027 => -59,
    53028 => -59,
    53029 => -59,
    53030 => -59,
    53031 => -59,
    53032 => -59,
    53033 => -59,
    53034 => -59,
    53035 => -59,
    53036 => -59,
    53037 => -59,
    53038 => -59,
    53039 => -59,
    53040 => -59,
    53041 => -59,
    53042 => -59,
    53043 => -59,
    53044 => -59,
    53045 => -59,
    53046 => -59,
    53047 => -59,
    53048 => -59,
    53049 => -59,
    53050 => -59,
    53051 => -59,
    53052 => -59,
    53053 => -59,
    53054 => -59,
    53055 => -59,
    53056 => -59,
    53057 => -59,
    53058 => -59,
    53059 => -59,
    53060 => -59,
    53061 => -59,
    53062 => -59,
    53063 => -59,
    53064 => -59,
    53065 => -59,
    53066 => -59,
    53067 => -59,
    53068 => -59,
    53069 => -59,
    53070 => -59,
    53071 => -59,
    53072 => -59,
    53073 => -59,
    53074 => -59,
    53075 => -59,
    53076 => -59,
    53077 => -59,
    53078 => -59,
    53079 => -59,
    53080 => -59,
    53081 => -59,
    53082 => -59,
    53083 => -59,
    53084 => -59,
    53085 => -59,
    53086 => -59,
    53087 => -59,
    53088 => -59,
    53089 => -59,
    53090 => -59,
    53091 => -59,
    53092 => -59,
    53093 => -59,
    53094 => -59,
    53095 => -59,
    53096 => -59,
    53097 => -59,
    53098 => -59,
    53099 => -59,
    53100 => -59,
    53101 => -59,
    53102 => -59,
    53103 => -59,
    53104 => -59,
    53105 => -59,
    53106 => -59,
    53107 => -59,
    53108 => -59,
    53109 => -59,
    53110 => -59,
    53111 => -59,
    53112 => -59,
    53113 => -59,
    53114 => -59,
    53115 => -59,
    53116 => -59,
    53117 => -59,
    53118 => -59,
    53119 => -58,
    53120 => -58,
    53121 => -58,
    53122 => -58,
    53123 => -58,
    53124 => -58,
    53125 => -58,
    53126 => -58,
    53127 => -58,
    53128 => -58,
    53129 => -58,
    53130 => -58,
    53131 => -58,
    53132 => -58,
    53133 => -58,
    53134 => -58,
    53135 => -58,
    53136 => -58,
    53137 => -58,
    53138 => -58,
    53139 => -58,
    53140 => -58,
    53141 => -58,
    53142 => -58,
    53143 => -58,
    53144 => -58,
    53145 => -58,
    53146 => -58,
    53147 => -58,
    53148 => -58,
    53149 => -58,
    53150 => -58,
    53151 => -58,
    53152 => -58,
    53153 => -58,
    53154 => -58,
    53155 => -58,
    53156 => -58,
    53157 => -58,
    53158 => -58,
    53159 => -58,
    53160 => -58,
    53161 => -58,
    53162 => -58,
    53163 => -58,
    53164 => -58,
    53165 => -58,
    53166 => -58,
    53167 => -58,
    53168 => -58,
    53169 => -58,
    53170 => -58,
    53171 => -58,
    53172 => -58,
    53173 => -58,
    53174 => -58,
    53175 => -58,
    53176 => -58,
    53177 => -58,
    53178 => -58,
    53179 => -58,
    53180 => -58,
    53181 => -58,
    53182 => -58,
    53183 => -58,
    53184 => -58,
    53185 => -58,
    53186 => -58,
    53187 => -58,
    53188 => -58,
    53189 => -58,
    53190 => -58,
    53191 => -58,
    53192 => -58,
    53193 => -58,
    53194 => -58,
    53195 => -58,
    53196 => -58,
    53197 => -58,
    53198 => -58,
    53199 => -58,
    53200 => -58,
    53201 => -58,
    53202 => -58,
    53203 => -58,
    53204 => -58,
    53205 => -58,
    53206 => -58,
    53207 => -58,
    53208 => -58,
    53209 => -58,
    53210 => -58,
    53211 => -58,
    53212 => -58,
    53213 => -58,
    53214 => -58,
    53215 => -58,
    53216 => -58,
    53217 => -58,
    53218 => -58,
    53219 => -58,
    53220 => -58,
    53221 => -58,
    53222 => -58,
    53223 => -58,
    53224 => -58,
    53225 => -58,
    53226 => -58,
    53227 => -58,
    53228 => -58,
    53229 => -58,
    53230 => -58,
    53231 => -58,
    53232 => -58,
    53233 => -58,
    53234 => -58,
    53235 => -58,
    53236 => -58,
    53237 => -58,
    53238 => -58,
    53239 => -58,
    53240 => -58,
    53241 => -58,
    53242 => -58,
    53243 => -58,
    53244 => -58,
    53245 => -58,
    53246 => -58,
    53247 => -58,
    53248 => -58,
    53249 => -58,
    53250 => -58,
    53251 => -58,
    53252 => -58,
    53253 => -58,
    53254 => -58,
    53255 => -58,
    53256 => -58,
    53257 => -58,
    53258 => -58,
    53259 => -58,
    53260 => -58,
    53261 => -58,
    53262 => -58,
    53263 => -58,
    53264 => -58,
    53265 => -58,
    53266 => -58,
    53267 => -58,
    53268 => -58,
    53269 => -58,
    53270 => -58,
    53271 => -58,
    53272 => -58,
    53273 => -58,
    53274 => -58,
    53275 => -58,
    53276 => -58,
    53277 => -58,
    53278 => -58,
    53279 => -58,
    53280 => -58,
    53281 => -58,
    53282 => -58,
    53283 => -58,
    53284 => -58,
    53285 => -58,
    53286 => -58,
    53287 => -58,
    53288 => -58,
    53289 => -58,
    53290 => -58,
    53291 => -58,
    53292 => -58,
    53293 => -58,
    53294 => -58,
    53295 => -58,
    53296 => -58,
    53297 => -58,
    53298 => -58,
    53299 => -58,
    53300 => -58,
    53301 => -58,
    53302 => -58,
    53303 => -58,
    53304 => -58,
    53305 => -58,
    53306 => -58,
    53307 => -58,
    53308 => -58,
    53309 => -58,
    53310 => -58,
    53311 => -58,
    53312 => -58,
    53313 => -58,
    53314 => -58,
    53315 => -58,
    53316 => -58,
    53317 => -58,
    53318 => -58,
    53319 => -58,
    53320 => -58,
    53321 => -58,
    53322 => -58,
    53323 => -58,
    53324 => -58,
    53325 => -58,
    53326 => -58,
    53327 => -58,
    53328 => -58,
    53329 => -58,
    53330 => -58,
    53331 => -58,
    53332 => -58,
    53333 => -58,
    53334 => -58,
    53335 => -58,
    53336 => -58,
    53337 => -58,
    53338 => -58,
    53339 => -58,
    53340 => -58,
    53341 => -58,
    53342 => -58,
    53343 => -58,
    53344 => -58,
    53345 => -58,
    53346 => -58,
    53347 => -58,
    53348 => -58,
    53349 => -58,
    53350 => -58,
    53351 => -58,
    53352 => -58,
    53353 => -58,
    53354 => -58,
    53355 => -58,
    53356 => -58,
    53357 => -58,
    53358 => -58,
    53359 => -58,
    53360 => -58,
    53361 => -58,
    53362 => -58,
    53363 => -58,
    53364 => -58,
    53365 => -58,
    53366 => -58,
    53367 => -58,
    53368 => -58,
    53369 => -58,
    53370 => -58,
    53371 => -58,
    53372 => -58,
    53373 => -58,
    53374 => -58,
    53375 => -58,
    53376 => -58,
    53377 => -58,
    53378 => -58,
    53379 => -58,
    53380 => -58,
    53381 => -58,
    53382 => -58,
    53383 => -58,
    53384 => -58,
    53385 => -58,
    53386 => -58,
    53387 => -58,
    53388 => -58,
    53389 => -58,
    53390 => -58,
    53391 => -58,
    53392 => -58,
    53393 => -58,
    53394 => -58,
    53395 => -58,
    53396 => -58,
    53397 => -58,
    53398 => -58,
    53399 => -58,
    53400 => -58,
    53401 => -58,
    53402 => -58,
    53403 => -58,
    53404 => -58,
    53405 => -58,
    53406 => -58,
    53407 => -58,
    53408 => -58,
    53409 => -58,
    53410 => -58,
    53411 => -58,
    53412 => -58,
    53413 => -58,
    53414 => -58,
    53415 => -58,
    53416 => -58,
    53417 => -58,
    53418 => -58,
    53419 => -58,
    53420 => -58,
    53421 => -58,
    53422 => -58,
    53423 => -58,
    53424 => -58,
    53425 => -58,
    53426 => -58,
    53427 => -58,
    53428 => -58,
    53429 => -58,
    53430 => -58,
    53431 => -58,
    53432 => -58,
    53433 => -58,
    53434 => -58,
    53435 => -58,
    53436 => -58,
    53437 => -58,
    53438 => -58,
    53439 => -58,
    53440 => -58,
    53441 => -58,
    53442 => -58,
    53443 => -58,
    53444 => -58,
    53445 => -58,
    53446 => -58,
    53447 => -58,
    53448 => -58,
    53449 => -58,
    53450 => -58,
    53451 => -58,
    53452 => -58,
    53453 => -58,
    53454 => -58,
    53455 => -58,
    53456 => -58,
    53457 => -58,
    53458 => -58,
    53459 => -58,
    53460 => -58,
    53461 => -58,
    53462 => -58,
    53463 => -58,
    53464 => -58,
    53465 => -58,
    53466 => -58,
    53467 => -58,
    53468 => -58,
    53469 => -58,
    53470 => -58,
    53471 => -58,
    53472 => -58,
    53473 => -58,
    53474 => -58,
    53475 => -58,
    53476 => -58,
    53477 => -58,
    53478 => -58,
    53479 => -58,
    53480 => -58,
    53481 => -58,
    53482 => -58,
    53483 => -58,
    53484 => -58,
    53485 => -58,
    53486 => -58,
    53487 => -58,
    53488 => -58,
    53489 => -58,
    53490 => -58,
    53491 => -58,
    53492 => -58,
    53493 => -58,
    53494 => -58,
    53495 => -58,
    53496 => -58,
    53497 => -58,
    53498 => -58,
    53499 => -58,
    53500 => -58,
    53501 => -58,
    53502 => -58,
    53503 => -58,
    53504 => -58,
    53505 => -58,
    53506 => -58,
    53507 => -58,
    53508 => -58,
    53509 => -58,
    53510 => -58,
    53511 => -58,
    53512 => -58,
    53513 => -58,
    53514 => -58,
    53515 => -58,
    53516 => -58,
    53517 => -58,
    53518 => -58,
    53519 => -58,
    53520 => -58,
    53521 => -58,
    53522 => -58,
    53523 => -58,
    53524 => -58,
    53525 => -58,
    53526 => -58,
    53527 => -58,
    53528 => -58,
    53529 => -58,
    53530 => -58,
    53531 => -58,
    53532 => -58,
    53533 => -58,
    53534 => -58,
    53535 => -58,
    53536 => -58,
    53537 => -58,
    53538 => -58,
    53539 => -58,
    53540 => -58,
    53541 => -58,
    53542 => -58,
    53543 => -57,
    53544 => -57,
    53545 => -57,
    53546 => -57,
    53547 => -57,
    53548 => -57,
    53549 => -57,
    53550 => -57,
    53551 => -57,
    53552 => -57,
    53553 => -57,
    53554 => -57,
    53555 => -57,
    53556 => -57,
    53557 => -57,
    53558 => -57,
    53559 => -57,
    53560 => -57,
    53561 => -57,
    53562 => -57,
    53563 => -57,
    53564 => -57,
    53565 => -57,
    53566 => -57,
    53567 => -57,
    53568 => -57,
    53569 => -57,
    53570 => -57,
    53571 => -57,
    53572 => -57,
    53573 => -57,
    53574 => -57,
    53575 => -57,
    53576 => -57,
    53577 => -57,
    53578 => -57,
    53579 => -57,
    53580 => -57,
    53581 => -57,
    53582 => -57,
    53583 => -57,
    53584 => -57,
    53585 => -57,
    53586 => -57,
    53587 => -57,
    53588 => -57,
    53589 => -57,
    53590 => -57,
    53591 => -57,
    53592 => -57,
    53593 => -57,
    53594 => -57,
    53595 => -57,
    53596 => -57,
    53597 => -57,
    53598 => -57,
    53599 => -57,
    53600 => -57,
    53601 => -57,
    53602 => -57,
    53603 => -57,
    53604 => -57,
    53605 => -57,
    53606 => -57,
    53607 => -57,
    53608 => -57,
    53609 => -57,
    53610 => -57,
    53611 => -57,
    53612 => -57,
    53613 => -57,
    53614 => -57,
    53615 => -57,
    53616 => -57,
    53617 => -57,
    53618 => -57,
    53619 => -57,
    53620 => -57,
    53621 => -57,
    53622 => -57,
    53623 => -57,
    53624 => -57,
    53625 => -57,
    53626 => -57,
    53627 => -57,
    53628 => -57,
    53629 => -57,
    53630 => -57,
    53631 => -57,
    53632 => -57,
    53633 => -57,
    53634 => -57,
    53635 => -57,
    53636 => -57,
    53637 => -57,
    53638 => -57,
    53639 => -57,
    53640 => -57,
    53641 => -57,
    53642 => -57,
    53643 => -57,
    53644 => -57,
    53645 => -57,
    53646 => -57,
    53647 => -57,
    53648 => -57,
    53649 => -57,
    53650 => -57,
    53651 => -57,
    53652 => -57,
    53653 => -57,
    53654 => -57,
    53655 => -57,
    53656 => -57,
    53657 => -57,
    53658 => -57,
    53659 => -57,
    53660 => -57,
    53661 => -57,
    53662 => -57,
    53663 => -57,
    53664 => -57,
    53665 => -57,
    53666 => -57,
    53667 => -57,
    53668 => -57,
    53669 => -57,
    53670 => -57,
    53671 => -57,
    53672 => -57,
    53673 => -57,
    53674 => -57,
    53675 => -57,
    53676 => -57,
    53677 => -57,
    53678 => -57,
    53679 => -57,
    53680 => -57,
    53681 => -57,
    53682 => -57,
    53683 => -57,
    53684 => -57,
    53685 => -57,
    53686 => -57,
    53687 => -57,
    53688 => -57,
    53689 => -57,
    53690 => -57,
    53691 => -57,
    53692 => -57,
    53693 => -57,
    53694 => -57,
    53695 => -57,
    53696 => -57,
    53697 => -57,
    53698 => -57,
    53699 => -57,
    53700 => -57,
    53701 => -57,
    53702 => -57,
    53703 => -57,
    53704 => -57,
    53705 => -57,
    53706 => -57,
    53707 => -57,
    53708 => -57,
    53709 => -57,
    53710 => -57,
    53711 => -57,
    53712 => -57,
    53713 => -57,
    53714 => -57,
    53715 => -57,
    53716 => -57,
    53717 => -57,
    53718 => -57,
    53719 => -57,
    53720 => -57,
    53721 => -57,
    53722 => -57,
    53723 => -57,
    53724 => -57,
    53725 => -57,
    53726 => -57,
    53727 => -57,
    53728 => -57,
    53729 => -57,
    53730 => -57,
    53731 => -57,
    53732 => -57,
    53733 => -57,
    53734 => -57,
    53735 => -57,
    53736 => -57,
    53737 => -57,
    53738 => -57,
    53739 => -57,
    53740 => -57,
    53741 => -57,
    53742 => -57,
    53743 => -57,
    53744 => -57,
    53745 => -57,
    53746 => -57,
    53747 => -57,
    53748 => -57,
    53749 => -57,
    53750 => -57,
    53751 => -57,
    53752 => -57,
    53753 => -57,
    53754 => -57,
    53755 => -57,
    53756 => -57,
    53757 => -57,
    53758 => -57,
    53759 => -57,
    53760 => -57,
    53761 => -57,
    53762 => -57,
    53763 => -57,
    53764 => -57,
    53765 => -57,
    53766 => -57,
    53767 => -57,
    53768 => -57,
    53769 => -57,
    53770 => -57,
    53771 => -57,
    53772 => -57,
    53773 => -57,
    53774 => -57,
    53775 => -57,
    53776 => -57,
    53777 => -57,
    53778 => -57,
    53779 => -57,
    53780 => -57,
    53781 => -57,
    53782 => -57,
    53783 => -57,
    53784 => -57,
    53785 => -57,
    53786 => -57,
    53787 => -57,
    53788 => -57,
    53789 => -57,
    53790 => -57,
    53791 => -57,
    53792 => -57,
    53793 => -57,
    53794 => -57,
    53795 => -57,
    53796 => -57,
    53797 => -57,
    53798 => -57,
    53799 => -57,
    53800 => -57,
    53801 => -57,
    53802 => -57,
    53803 => -57,
    53804 => -57,
    53805 => -57,
    53806 => -57,
    53807 => -57,
    53808 => -57,
    53809 => -57,
    53810 => -57,
    53811 => -57,
    53812 => -57,
    53813 => -57,
    53814 => -57,
    53815 => -57,
    53816 => -57,
    53817 => -57,
    53818 => -57,
    53819 => -57,
    53820 => -57,
    53821 => -57,
    53822 => -57,
    53823 => -57,
    53824 => -57,
    53825 => -57,
    53826 => -57,
    53827 => -57,
    53828 => -57,
    53829 => -57,
    53830 => -57,
    53831 => -57,
    53832 => -57,
    53833 => -57,
    53834 => -57,
    53835 => -57,
    53836 => -57,
    53837 => -57,
    53838 => -57,
    53839 => -57,
    53840 => -57,
    53841 => -57,
    53842 => -57,
    53843 => -57,
    53844 => -57,
    53845 => -57,
    53846 => -57,
    53847 => -57,
    53848 => -57,
    53849 => -57,
    53850 => -57,
    53851 => -57,
    53852 => -57,
    53853 => -57,
    53854 => -57,
    53855 => -57,
    53856 => -57,
    53857 => -57,
    53858 => -57,
    53859 => -57,
    53860 => -57,
    53861 => -57,
    53862 => -57,
    53863 => -57,
    53864 => -57,
    53865 => -57,
    53866 => -57,
    53867 => -57,
    53868 => -57,
    53869 => -57,
    53870 => -57,
    53871 => -57,
    53872 => -57,
    53873 => -57,
    53874 => -57,
    53875 => -57,
    53876 => -57,
    53877 => -57,
    53878 => -57,
    53879 => -57,
    53880 => -57,
    53881 => -57,
    53882 => -57,
    53883 => -57,
    53884 => -57,
    53885 => -57,
    53886 => -57,
    53887 => -57,
    53888 => -57,
    53889 => -57,
    53890 => -57,
    53891 => -57,
    53892 => -57,
    53893 => -57,
    53894 => -57,
    53895 => -57,
    53896 => -57,
    53897 => -57,
    53898 => -57,
    53899 => -57,
    53900 => -57,
    53901 => -57,
    53902 => -57,
    53903 => -57,
    53904 => -57,
    53905 => -57,
    53906 => -57,
    53907 => -57,
    53908 => -57,
    53909 => -57,
    53910 => -57,
    53911 => -57,
    53912 => -57,
    53913 => -57,
    53914 => -57,
    53915 => -57,
    53916 => -57,
    53917 => -57,
    53918 => -57,
    53919 => -57,
    53920 => -57,
    53921 => -57,
    53922 => -57,
    53923 => -57,
    53924 => -57,
    53925 => -57,
    53926 => -57,
    53927 => -57,
    53928 => -57,
    53929 => -57,
    53930 => -57,
    53931 => -57,
    53932 => -56,
    53933 => -56,
    53934 => -56,
    53935 => -56,
    53936 => -56,
    53937 => -56,
    53938 => -56,
    53939 => -56,
    53940 => -56,
    53941 => -56,
    53942 => -56,
    53943 => -56,
    53944 => -56,
    53945 => -56,
    53946 => -56,
    53947 => -56,
    53948 => -56,
    53949 => -56,
    53950 => -56,
    53951 => -56,
    53952 => -56,
    53953 => -56,
    53954 => -56,
    53955 => -56,
    53956 => -56,
    53957 => -56,
    53958 => -56,
    53959 => -56,
    53960 => -56,
    53961 => -56,
    53962 => -56,
    53963 => -56,
    53964 => -56,
    53965 => -56,
    53966 => -56,
    53967 => -56,
    53968 => -56,
    53969 => -56,
    53970 => -56,
    53971 => -56,
    53972 => -56,
    53973 => -56,
    53974 => -56,
    53975 => -56,
    53976 => -56,
    53977 => -56,
    53978 => -56,
    53979 => -56,
    53980 => -56,
    53981 => -56,
    53982 => -56,
    53983 => -56,
    53984 => -56,
    53985 => -56,
    53986 => -56,
    53987 => -56,
    53988 => -56,
    53989 => -56,
    53990 => -56,
    53991 => -56,
    53992 => -56,
    53993 => -56,
    53994 => -56,
    53995 => -56,
    53996 => -56,
    53997 => -56,
    53998 => -56,
    53999 => -56,
    54000 => -56,
    54001 => -56,
    54002 => -56,
    54003 => -56,
    54004 => -56,
    54005 => -56,
    54006 => -56,
    54007 => -56,
    54008 => -56,
    54009 => -56,
    54010 => -56,
    54011 => -56,
    54012 => -56,
    54013 => -56,
    54014 => -56,
    54015 => -56,
    54016 => -56,
    54017 => -56,
    54018 => -56,
    54019 => -56,
    54020 => -56,
    54021 => -56,
    54022 => -56,
    54023 => -56,
    54024 => -56,
    54025 => -56,
    54026 => -56,
    54027 => -56,
    54028 => -56,
    54029 => -56,
    54030 => -56,
    54031 => -56,
    54032 => -56,
    54033 => -56,
    54034 => -56,
    54035 => -56,
    54036 => -56,
    54037 => -56,
    54038 => -56,
    54039 => -56,
    54040 => -56,
    54041 => -56,
    54042 => -56,
    54043 => -56,
    54044 => -56,
    54045 => -56,
    54046 => -56,
    54047 => -56,
    54048 => -56,
    54049 => -56,
    54050 => -56,
    54051 => -56,
    54052 => -56,
    54053 => -56,
    54054 => -56,
    54055 => -56,
    54056 => -56,
    54057 => -56,
    54058 => -56,
    54059 => -56,
    54060 => -56,
    54061 => -56,
    54062 => -56,
    54063 => -56,
    54064 => -56,
    54065 => -56,
    54066 => -56,
    54067 => -56,
    54068 => -56,
    54069 => -56,
    54070 => -56,
    54071 => -56,
    54072 => -56,
    54073 => -56,
    54074 => -56,
    54075 => -56,
    54076 => -56,
    54077 => -56,
    54078 => -56,
    54079 => -56,
    54080 => -56,
    54081 => -56,
    54082 => -56,
    54083 => -56,
    54084 => -56,
    54085 => -56,
    54086 => -56,
    54087 => -56,
    54088 => -56,
    54089 => -56,
    54090 => -56,
    54091 => -56,
    54092 => -56,
    54093 => -56,
    54094 => -56,
    54095 => -56,
    54096 => -56,
    54097 => -56,
    54098 => -56,
    54099 => -56,
    54100 => -56,
    54101 => -56,
    54102 => -56,
    54103 => -56,
    54104 => -56,
    54105 => -56,
    54106 => -56,
    54107 => -56,
    54108 => -56,
    54109 => -56,
    54110 => -56,
    54111 => -56,
    54112 => -56,
    54113 => -56,
    54114 => -56,
    54115 => -56,
    54116 => -56,
    54117 => -56,
    54118 => -56,
    54119 => -56,
    54120 => -56,
    54121 => -56,
    54122 => -56,
    54123 => -56,
    54124 => -56,
    54125 => -56,
    54126 => -56,
    54127 => -56,
    54128 => -56,
    54129 => -56,
    54130 => -56,
    54131 => -56,
    54132 => -56,
    54133 => -56,
    54134 => -56,
    54135 => -56,
    54136 => -56,
    54137 => -56,
    54138 => -56,
    54139 => -56,
    54140 => -56,
    54141 => -56,
    54142 => -56,
    54143 => -56,
    54144 => -56,
    54145 => -56,
    54146 => -56,
    54147 => -56,
    54148 => -56,
    54149 => -56,
    54150 => -56,
    54151 => -56,
    54152 => -56,
    54153 => -56,
    54154 => -56,
    54155 => -56,
    54156 => -56,
    54157 => -56,
    54158 => -56,
    54159 => -56,
    54160 => -56,
    54161 => -56,
    54162 => -56,
    54163 => -56,
    54164 => -56,
    54165 => -56,
    54166 => -56,
    54167 => -56,
    54168 => -56,
    54169 => -56,
    54170 => -56,
    54171 => -56,
    54172 => -56,
    54173 => -56,
    54174 => -56,
    54175 => -56,
    54176 => -56,
    54177 => -56,
    54178 => -56,
    54179 => -56,
    54180 => -56,
    54181 => -56,
    54182 => -56,
    54183 => -56,
    54184 => -56,
    54185 => -56,
    54186 => -56,
    54187 => -56,
    54188 => -56,
    54189 => -56,
    54190 => -56,
    54191 => -56,
    54192 => -56,
    54193 => -56,
    54194 => -56,
    54195 => -56,
    54196 => -56,
    54197 => -56,
    54198 => -56,
    54199 => -56,
    54200 => -56,
    54201 => -56,
    54202 => -56,
    54203 => -56,
    54204 => -56,
    54205 => -56,
    54206 => -56,
    54207 => -56,
    54208 => -56,
    54209 => -56,
    54210 => -56,
    54211 => -56,
    54212 => -56,
    54213 => -56,
    54214 => -56,
    54215 => -56,
    54216 => -56,
    54217 => -56,
    54218 => -56,
    54219 => -56,
    54220 => -56,
    54221 => -56,
    54222 => -56,
    54223 => -56,
    54224 => -56,
    54225 => -56,
    54226 => -56,
    54227 => -56,
    54228 => -56,
    54229 => -56,
    54230 => -56,
    54231 => -56,
    54232 => -56,
    54233 => -56,
    54234 => -56,
    54235 => -56,
    54236 => -56,
    54237 => -56,
    54238 => -56,
    54239 => -56,
    54240 => -56,
    54241 => -56,
    54242 => -56,
    54243 => -56,
    54244 => -56,
    54245 => -56,
    54246 => -56,
    54247 => -56,
    54248 => -56,
    54249 => -56,
    54250 => -56,
    54251 => -56,
    54252 => -56,
    54253 => -56,
    54254 => -56,
    54255 => -56,
    54256 => -56,
    54257 => -56,
    54258 => -56,
    54259 => -56,
    54260 => -56,
    54261 => -56,
    54262 => -56,
    54263 => -56,
    54264 => -56,
    54265 => -56,
    54266 => -56,
    54267 => -56,
    54268 => -56,
    54269 => -56,
    54270 => -56,
    54271 => -56,
    54272 => -56,
    54273 => -56,
    54274 => -56,
    54275 => -56,
    54276 => -56,
    54277 => -56,
    54278 => -56,
    54279 => -56,
    54280 => -56,
    54281 => -56,
    54282 => -56,
    54283 => -56,
    54284 => -56,
    54285 => -56,
    54286 => -56,
    54287 => -56,
    54288 => -56,
    54289 => -56,
    54290 => -56,
    54291 => -56,
    54292 => -56,
    54293 => -56,
    54294 => -55,
    54295 => -55,
    54296 => -55,
    54297 => -55,
    54298 => -55,
    54299 => -55,
    54300 => -55,
    54301 => -55,
    54302 => -55,
    54303 => -55,
    54304 => -55,
    54305 => -55,
    54306 => -55,
    54307 => -55,
    54308 => -55,
    54309 => -55,
    54310 => -55,
    54311 => -55,
    54312 => -55,
    54313 => -55,
    54314 => -55,
    54315 => -55,
    54316 => -55,
    54317 => -55,
    54318 => -55,
    54319 => -55,
    54320 => -55,
    54321 => -55,
    54322 => -55,
    54323 => -55,
    54324 => -55,
    54325 => -55,
    54326 => -55,
    54327 => -55,
    54328 => -55,
    54329 => -55,
    54330 => -55,
    54331 => -55,
    54332 => -55,
    54333 => -55,
    54334 => -55,
    54335 => -55,
    54336 => -55,
    54337 => -55,
    54338 => -55,
    54339 => -55,
    54340 => -55,
    54341 => -55,
    54342 => -55,
    54343 => -55,
    54344 => -55,
    54345 => -55,
    54346 => -55,
    54347 => -55,
    54348 => -55,
    54349 => -55,
    54350 => -55,
    54351 => -55,
    54352 => -55,
    54353 => -55,
    54354 => -55,
    54355 => -55,
    54356 => -55,
    54357 => -55,
    54358 => -55,
    54359 => -55,
    54360 => -55,
    54361 => -55,
    54362 => -55,
    54363 => -55,
    54364 => -55,
    54365 => -55,
    54366 => -55,
    54367 => -55,
    54368 => -55,
    54369 => -55,
    54370 => -55,
    54371 => -55,
    54372 => -55,
    54373 => -55,
    54374 => -55,
    54375 => -55,
    54376 => -55,
    54377 => -55,
    54378 => -55,
    54379 => -55,
    54380 => -55,
    54381 => -55,
    54382 => -55,
    54383 => -55,
    54384 => -55,
    54385 => -55,
    54386 => -55,
    54387 => -55,
    54388 => -55,
    54389 => -55,
    54390 => -55,
    54391 => -55,
    54392 => -55,
    54393 => -55,
    54394 => -55,
    54395 => -55,
    54396 => -55,
    54397 => -55,
    54398 => -55,
    54399 => -55,
    54400 => -55,
    54401 => -55,
    54402 => -55,
    54403 => -55,
    54404 => -55,
    54405 => -55,
    54406 => -55,
    54407 => -55,
    54408 => -55,
    54409 => -55,
    54410 => -55,
    54411 => -55,
    54412 => -55,
    54413 => -55,
    54414 => -55,
    54415 => -55,
    54416 => -55,
    54417 => -55,
    54418 => -55,
    54419 => -55,
    54420 => -55,
    54421 => -55,
    54422 => -55,
    54423 => -55,
    54424 => -55,
    54425 => -55,
    54426 => -55,
    54427 => -55,
    54428 => -55,
    54429 => -55,
    54430 => -55,
    54431 => -55,
    54432 => -55,
    54433 => -55,
    54434 => -55,
    54435 => -55,
    54436 => -55,
    54437 => -55,
    54438 => -55,
    54439 => -55,
    54440 => -55,
    54441 => -55,
    54442 => -55,
    54443 => -55,
    54444 => -55,
    54445 => -55,
    54446 => -55,
    54447 => -55,
    54448 => -55,
    54449 => -55,
    54450 => -55,
    54451 => -55,
    54452 => -55,
    54453 => -55,
    54454 => -55,
    54455 => -55,
    54456 => -55,
    54457 => -55,
    54458 => -55,
    54459 => -55,
    54460 => -55,
    54461 => -55,
    54462 => -55,
    54463 => -55,
    54464 => -55,
    54465 => -55,
    54466 => -55,
    54467 => -55,
    54468 => -55,
    54469 => -55,
    54470 => -55,
    54471 => -55,
    54472 => -55,
    54473 => -55,
    54474 => -55,
    54475 => -55,
    54476 => -55,
    54477 => -55,
    54478 => -55,
    54479 => -55,
    54480 => -55,
    54481 => -55,
    54482 => -55,
    54483 => -55,
    54484 => -55,
    54485 => -55,
    54486 => -55,
    54487 => -55,
    54488 => -55,
    54489 => -55,
    54490 => -55,
    54491 => -55,
    54492 => -55,
    54493 => -55,
    54494 => -55,
    54495 => -55,
    54496 => -55,
    54497 => -55,
    54498 => -55,
    54499 => -55,
    54500 => -55,
    54501 => -55,
    54502 => -55,
    54503 => -55,
    54504 => -55,
    54505 => -55,
    54506 => -55,
    54507 => -55,
    54508 => -55,
    54509 => -55,
    54510 => -55,
    54511 => -55,
    54512 => -55,
    54513 => -55,
    54514 => -55,
    54515 => -55,
    54516 => -55,
    54517 => -55,
    54518 => -55,
    54519 => -55,
    54520 => -55,
    54521 => -55,
    54522 => -55,
    54523 => -55,
    54524 => -55,
    54525 => -55,
    54526 => -55,
    54527 => -55,
    54528 => -55,
    54529 => -55,
    54530 => -55,
    54531 => -55,
    54532 => -55,
    54533 => -55,
    54534 => -55,
    54535 => -55,
    54536 => -55,
    54537 => -55,
    54538 => -55,
    54539 => -55,
    54540 => -55,
    54541 => -55,
    54542 => -55,
    54543 => -55,
    54544 => -55,
    54545 => -55,
    54546 => -55,
    54547 => -55,
    54548 => -55,
    54549 => -55,
    54550 => -55,
    54551 => -55,
    54552 => -55,
    54553 => -55,
    54554 => -55,
    54555 => -55,
    54556 => -55,
    54557 => -55,
    54558 => -55,
    54559 => -55,
    54560 => -55,
    54561 => -55,
    54562 => -55,
    54563 => -55,
    54564 => -55,
    54565 => -55,
    54566 => -55,
    54567 => -55,
    54568 => -55,
    54569 => -55,
    54570 => -55,
    54571 => -55,
    54572 => -55,
    54573 => -55,
    54574 => -55,
    54575 => -55,
    54576 => -55,
    54577 => -55,
    54578 => -55,
    54579 => -55,
    54580 => -55,
    54581 => -55,
    54582 => -55,
    54583 => -55,
    54584 => -55,
    54585 => -55,
    54586 => -55,
    54587 => -55,
    54588 => -55,
    54589 => -55,
    54590 => -55,
    54591 => -55,
    54592 => -55,
    54593 => -55,
    54594 => -55,
    54595 => -55,
    54596 => -55,
    54597 => -55,
    54598 => -55,
    54599 => -55,
    54600 => -55,
    54601 => -55,
    54602 => -55,
    54603 => -55,
    54604 => -55,
    54605 => -55,
    54606 => -55,
    54607 => -55,
    54608 => -55,
    54609 => -55,
    54610 => -55,
    54611 => -55,
    54612 => -55,
    54613 => -55,
    54614 => -55,
    54615 => -55,
    54616 => -55,
    54617 => -55,
    54618 => -55,
    54619 => -55,
    54620 => -55,
    54621 => -55,
    54622 => -55,
    54623 => -55,
    54624 => -55,
    54625 => -55,
    54626 => -55,
    54627 => -55,
    54628 => -55,
    54629 => -55,
    54630 => -55,
    54631 => -55,
    54632 => -55,
    54633 => -55,
    54634 => -54,
    54635 => -54,
    54636 => -54,
    54637 => -54,
    54638 => -54,
    54639 => -54,
    54640 => -54,
    54641 => -54,
    54642 => -54,
    54643 => -54,
    54644 => -54,
    54645 => -54,
    54646 => -54,
    54647 => -54,
    54648 => -54,
    54649 => -54,
    54650 => -54,
    54651 => -54,
    54652 => -54,
    54653 => -54,
    54654 => -54,
    54655 => -54,
    54656 => -54,
    54657 => -54,
    54658 => -54,
    54659 => -54,
    54660 => -54,
    54661 => -54,
    54662 => -54,
    54663 => -54,
    54664 => -54,
    54665 => -54,
    54666 => -54,
    54667 => -54,
    54668 => -54,
    54669 => -54,
    54670 => -54,
    54671 => -54,
    54672 => -54,
    54673 => -54,
    54674 => -54,
    54675 => -54,
    54676 => -54,
    54677 => -54,
    54678 => -54,
    54679 => -54,
    54680 => -54,
    54681 => -54,
    54682 => -54,
    54683 => -54,
    54684 => -54,
    54685 => -54,
    54686 => -54,
    54687 => -54,
    54688 => -54,
    54689 => -54,
    54690 => -54,
    54691 => -54,
    54692 => -54,
    54693 => -54,
    54694 => -54,
    54695 => -54,
    54696 => -54,
    54697 => -54,
    54698 => -54,
    54699 => -54,
    54700 => -54,
    54701 => -54,
    54702 => -54,
    54703 => -54,
    54704 => -54,
    54705 => -54,
    54706 => -54,
    54707 => -54,
    54708 => -54,
    54709 => -54,
    54710 => -54,
    54711 => -54,
    54712 => -54,
    54713 => -54,
    54714 => -54,
    54715 => -54,
    54716 => -54,
    54717 => -54,
    54718 => -54,
    54719 => -54,
    54720 => -54,
    54721 => -54,
    54722 => -54,
    54723 => -54,
    54724 => -54,
    54725 => -54,
    54726 => -54,
    54727 => -54,
    54728 => -54,
    54729 => -54,
    54730 => -54,
    54731 => -54,
    54732 => -54,
    54733 => -54,
    54734 => -54,
    54735 => -54,
    54736 => -54,
    54737 => -54,
    54738 => -54,
    54739 => -54,
    54740 => -54,
    54741 => -54,
    54742 => -54,
    54743 => -54,
    54744 => -54,
    54745 => -54,
    54746 => -54,
    54747 => -54,
    54748 => -54,
    54749 => -54,
    54750 => -54,
    54751 => -54,
    54752 => -54,
    54753 => -54,
    54754 => -54,
    54755 => -54,
    54756 => -54,
    54757 => -54,
    54758 => -54,
    54759 => -54,
    54760 => -54,
    54761 => -54,
    54762 => -54,
    54763 => -54,
    54764 => -54,
    54765 => -54,
    54766 => -54,
    54767 => -54,
    54768 => -54,
    54769 => -54,
    54770 => -54,
    54771 => -54,
    54772 => -54,
    54773 => -54,
    54774 => -54,
    54775 => -54,
    54776 => -54,
    54777 => -54,
    54778 => -54,
    54779 => -54,
    54780 => -54,
    54781 => -54,
    54782 => -54,
    54783 => -54,
    54784 => -54,
    54785 => -54,
    54786 => -54,
    54787 => -54,
    54788 => -54,
    54789 => -54,
    54790 => -54,
    54791 => -54,
    54792 => -54,
    54793 => -54,
    54794 => -54,
    54795 => -54,
    54796 => -54,
    54797 => -54,
    54798 => -54,
    54799 => -54,
    54800 => -54,
    54801 => -54,
    54802 => -54,
    54803 => -54,
    54804 => -54,
    54805 => -54,
    54806 => -54,
    54807 => -54,
    54808 => -54,
    54809 => -54,
    54810 => -54,
    54811 => -54,
    54812 => -54,
    54813 => -54,
    54814 => -54,
    54815 => -54,
    54816 => -54,
    54817 => -54,
    54818 => -54,
    54819 => -54,
    54820 => -54,
    54821 => -54,
    54822 => -54,
    54823 => -54,
    54824 => -54,
    54825 => -54,
    54826 => -54,
    54827 => -54,
    54828 => -54,
    54829 => -54,
    54830 => -54,
    54831 => -54,
    54832 => -54,
    54833 => -54,
    54834 => -54,
    54835 => -54,
    54836 => -54,
    54837 => -54,
    54838 => -54,
    54839 => -54,
    54840 => -54,
    54841 => -54,
    54842 => -54,
    54843 => -54,
    54844 => -54,
    54845 => -54,
    54846 => -54,
    54847 => -54,
    54848 => -54,
    54849 => -54,
    54850 => -54,
    54851 => -54,
    54852 => -54,
    54853 => -54,
    54854 => -54,
    54855 => -54,
    54856 => -54,
    54857 => -54,
    54858 => -54,
    54859 => -54,
    54860 => -54,
    54861 => -54,
    54862 => -54,
    54863 => -54,
    54864 => -54,
    54865 => -54,
    54866 => -54,
    54867 => -54,
    54868 => -54,
    54869 => -54,
    54870 => -54,
    54871 => -54,
    54872 => -54,
    54873 => -54,
    54874 => -54,
    54875 => -54,
    54876 => -54,
    54877 => -54,
    54878 => -54,
    54879 => -54,
    54880 => -54,
    54881 => -54,
    54882 => -54,
    54883 => -54,
    54884 => -54,
    54885 => -54,
    54886 => -54,
    54887 => -54,
    54888 => -54,
    54889 => -54,
    54890 => -54,
    54891 => -54,
    54892 => -54,
    54893 => -54,
    54894 => -54,
    54895 => -54,
    54896 => -54,
    54897 => -54,
    54898 => -54,
    54899 => -54,
    54900 => -54,
    54901 => -54,
    54902 => -54,
    54903 => -54,
    54904 => -54,
    54905 => -54,
    54906 => -54,
    54907 => -54,
    54908 => -54,
    54909 => -54,
    54910 => -54,
    54911 => -54,
    54912 => -54,
    54913 => -54,
    54914 => -54,
    54915 => -54,
    54916 => -54,
    54917 => -54,
    54918 => -54,
    54919 => -54,
    54920 => -54,
    54921 => -54,
    54922 => -54,
    54923 => -54,
    54924 => -54,
    54925 => -54,
    54926 => -54,
    54927 => -54,
    54928 => -54,
    54929 => -54,
    54930 => -54,
    54931 => -54,
    54932 => -54,
    54933 => -54,
    54934 => -54,
    54935 => -54,
    54936 => -54,
    54937 => -54,
    54938 => -54,
    54939 => -54,
    54940 => -54,
    54941 => -54,
    54942 => -54,
    54943 => -54,
    54944 => -54,
    54945 => -54,
    54946 => -54,
    54947 => -54,
    54948 => -54,
    54949 => -54,
    54950 => -54,
    54951 => -54,
    54952 => -54,
    54953 => -54,
    54954 => -54,
    54955 => -53,
    54956 => -53,
    54957 => -53,
    54958 => -53,
    54959 => -53,
    54960 => -53,
    54961 => -53,
    54962 => -53,
    54963 => -53,
    54964 => -53,
    54965 => -53,
    54966 => -53,
    54967 => -53,
    54968 => -53,
    54969 => -53,
    54970 => -53,
    54971 => -53,
    54972 => -53,
    54973 => -53,
    54974 => -53,
    54975 => -53,
    54976 => -53,
    54977 => -53,
    54978 => -53,
    54979 => -53,
    54980 => -53,
    54981 => -53,
    54982 => -53,
    54983 => -53,
    54984 => -53,
    54985 => -53,
    54986 => -53,
    54987 => -53,
    54988 => -53,
    54989 => -53,
    54990 => -53,
    54991 => -53,
    54992 => -53,
    54993 => -53,
    54994 => -53,
    54995 => -53,
    54996 => -53,
    54997 => -53,
    54998 => -53,
    54999 => -53,
    55000 => -53,
    55001 => -53,
    55002 => -53,
    55003 => -53,
    55004 => -53,
    55005 => -53,
    55006 => -53,
    55007 => -53,
    55008 => -53,
    55009 => -53,
    55010 => -53,
    55011 => -53,
    55012 => -53,
    55013 => -53,
    55014 => -53,
    55015 => -53,
    55016 => -53,
    55017 => -53,
    55018 => -53,
    55019 => -53,
    55020 => -53,
    55021 => -53,
    55022 => -53,
    55023 => -53,
    55024 => -53,
    55025 => -53,
    55026 => -53,
    55027 => -53,
    55028 => -53,
    55029 => -53,
    55030 => -53,
    55031 => -53,
    55032 => -53,
    55033 => -53,
    55034 => -53,
    55035 => -53,
    55036 => -53,
    55037 => -53,
    55038 => -53,
    55039 => -53,
    55040 => -53,
    55041 => -53,
    55042 => -53,
    55043 => -53,
    55044 => -53,
    55045 => -53,
    55046 => -53,
    55047 => -53,
    55048 => -53,
    55049 => -53,
    55050 => -53,
    55051 => -53,
    55052 => -53,
    55053 => -53,
    55054 => -53,
    55055 => -53,
    55056 => -53,
    55057 => -53,
    55058 => -53,
    55059 => -53,
    55060 => -53,
    55061 => -53,
    55062 => -53,
    55063 => -53,
    55064 => -53,
    55065 => -53,
    55066 => -53,
    55067 => -53,
    55068 => -53,
    55069 => -53,
    55070 => -53,
    55071 => -53,
    55072 => -53,
    55073 => -53,
    55074 => -53,
    55075 => -53,
    55076 => -53,
    55077 => -53,
    55078 => -53,
    55079 => -53,
    55080 => -53,
    55081 => -53,
    55082 => -53,
    55083 => -53,
    55084 => -53,
    55085 => -53,
    55086 => -53,
    55087 => -53,
    55088 => -53,
    55089 => -53,
    55090 => -53,
    55091 => -53,
    55092 => -53,
    55093 => -53,
    55094 => -53,
    55095 => -53,
    55096 => -53,
    55097 => -53,
    55098 => -53,
    55099 => -53,
    55100 => -53,
    55101 => -53,
    55102 => -53,
    55103 => -53,
    55104 => -53,
    55105 => -53,
    55106 => -53,
    55107 => -53,
    55108 => -53,
    55109 => -53,
    55110 => -53,
    55111 => -53,
    55112 => -53,
    55113 => -53,
    55114 => -53,
    55115 => -53,
    55116 => -53,
    55117 => -53,
    55118 => -53,
    55119 => -53,
    55120 => -53,
    55121 => -53,
    55122 => -53,
    55123 => -53,
    55124 => -53,
    55125 => -53,
    55126 => -53,
    55127 => -53,
    55128 => -53,
    55129 => -53,
    55130 => -53,
    55131 => -53,
    55132 => -53,
    55133 => -53,
    55134 => -53,
    55135 => -53,
    55136 => -53,
    55137 => -53,
    55138 => -53,
    55139 => -53,
    55140 => -53,
    55141 => -53,
    55142 => -53,
    55143 => -53,
    55144 => -53,
    55145 => -53,
    55146 => -53,
    55147 => -53,
    55148 => -53,
    55149 => -53,
    55150 => -53,
    55151 => -53,
    55152 => -53,
    55153 => -53,
    55154 => -53,
    55155 => -53,
    55156 => -53,
    55157 => -53,
    55158 => -53,
    55159 => -53,
    55160 => -53,
    55161 => -53,
    55162 => -53,
    55163 => -53,
    55164 => -53,
    55165 => -53,
    55166 => -53,
    55167 => -53,
    55168 => -53,
    55169 => -53,
    55170 => -53,
    55171 => -53,
    55172 => -53,
    55173 => -53,
    55174 => -53,
    55175 => -53,
    55176 => -53,
    55177 => -53,
    55178 => -53,
    55179 => -53,
    55180 => -53,
    55181 => -53,
    55182 => -53,
    55183 => -53,
    55184 => -53,
    55185 => -53,
    55186 => -53,
    55187 => -53,
    55188 => -53,
    55189 => -53,
    55190 => -53,
    55191 => -53,
    55192 => -53,
    55193 => -53,
    55194 => -53,
    55195 => -53,
    55196 => -53,
    55197 => -53,
    55198 => -53,
    55199 => -53,
    55200 => -53,
    55201 => -53,
    55202 => -53,
    55203 => -53,
    55204 => -53,
    55205 => -53,
    55206 => -53,
    55207 => -53,
    55208 => -53,
    55209 => -53,
    55210 => -53,
    55211 => -53,
    55212 => -53,
    55213 => -53,
    55214 => -53,
    55215 => -53,
    55216 => -53,
    55217 => -53,
    55218 => -53,
    55219 => -53,
    55220 => -53,
    55221 => -53,
    55222 => -53,
    55223 => -53,
    55224 => -53,
    55225 => -53,
    55226 => -53,
    55227 => -53,
    55228 => -53,
    55229 => -53,
    55230 => -53,
    55231 => -53,
    55232 => -53,
    55233 => -53,
    55234 => -53,
    55235 => -53,
    55236 => -53,
    55237 => -53,
    55238 => -53,
    55239 => -53,
    55240 => -53,
    55241 => -53,
    55242 => -53,
    55243 => -53,
    55244 => -53,
    55245 => -53,
    55246 => -53,
    55247 => -53,
    55248 => -53,
    55249 => -53,
    55250 => -53,
    55251 => -53,
    55252 => -53,
    55253 => -53,
    55254 => -53,
    55255 => -53,
    55256 => -53,
    55257 => -53,
    55258 => -53,
    55259 => -53,
    55260 => -53,
    55261 => -52,
    55262 => -52,
    55263 => -52,
    55264 => -52,
    55265 => -52,
    55266 => -52,
    55267 => -52,
    55268 => -52,
    55269 => -52,
    55270 => -52,
    55271 => -52,
    55272 => -52,
    55273 => -52,
    55274 => -52,
    55275 => -52,
    55276 => -52,
    55277 => -52,
    55278 => -52,
    55279 => -52,
    55280 => -52,
    55281 => -52,
    55282 => -52,
    55283 => -52,
    55284 => -52,
    55285 => -52,
    55286 => -52,
    55287 => -52,
    55288 => -52,
    55289 => -52,
    55290 => -52,
    55291 => -52,
    55292 => -52,
    55293 => -52,
    55294 => -52,
    55295 => -52,
    55296 => -52,
    55297 => -52,
    55298 => -52,
    55299 => -52,
    55300 => -52,
    55301 => -52,
    55302 => -52,
    55303 => -52,
    55304 => -52,
    55305 => -52,
    55306 => -52,
    55307 => -52,
    55308 => -52,
    55309 => -52,
    55310 => -52,
    55311 => -52,
    55312 => -52,
    55313 => -52,
    55314 => -52,
    55315 => -52,
    55316 => -52,
    55317 => -52,
    55318 => -52,
    55319 => -52,
    55320 => -52,
    55321 => -52,
    55322 => -52,
    55323 => -52,
    55324 => -52,
    55325 => -52,
    55326 => -52,
    55327 => -52,
    55328 => -52,
    55329 => -52,
    55330 => -52,
    55331 => -52,
    55332 => -52,
    55333 => -52,
    55334 => -52,
    55335 => -52,
    55336 => -52,
    55337 => -52,
    55338 => -52,
    55339 => -52,
    55340 => -52,
    55341 => -52,
    55342 => -52,
    55343 => -52,
    55344 => -52,
    55345 => -52,
    55346 => -52,
    55347 => -52,
    55348 => -52,
    55349 => -52,
    55350 => -52,
    55351 => -52,
    55352 => -52,
    55353 => -52,
    55354 => -52,
    55355 => -52,
    55356 => -52,
    55357 => -52,
    55358 => -52,
    55359 => -52,
    55360 => -52,
    55361 => -52,
    55362 => -52,
    55363 => -52,
    55364 => -52,
    55365 => -52,
    55366 => -52,
    55367 => -52,
    55368 => -52,
    55369 => -52,
    55370 => -52,
    55371 => -52,
    55372 => -52,
    55373 => -52,
    55374 => -52,
    55375 => -52,
    55376 => -52,
    55377 => -52,
    55378 => -52,
    55379 => -52,
    55380 => -52,
    55381 => -52,
    55382 => -52,
    55383 => -52,
    55384 => -52,
    55385 => -52,
    55386 => -52,
    55387 => -52,
    55388 => -52,
    55389 => -52,
    55390 => -52,
    55391 => -52,
    55392 => -52,
    55393 => -52,
    55394 => -52,
    55395 => -52,
    55396 => -52,
    55397 => -52,
    55398 => -52,
    55399 => -52,
    55400 => -52,
    55401 => -52,
    55402 => -52,
    55403 => -52,
    55404 => -52,
    55405 => -52,
    55406 => -52,
    55407 => -52,
    55408 => -52,
    55409 => -52,
    55410 => -52,
    55411 => -52,
    55412 => -52,
    55413 => -52,
    55414 => -52,
    55415 => -52,
    55416 => -52,
    55417 => -52,
    55418 => -52,
    55419 => -52,
    55420 => -52,
    55421 => -52,
    55422 => -52,
    55423 => -52,
    55424 => -52,
    55425 => -52,
    55426 => -52,
    55427 => -52,
    55428 => -52,
    55429 => -52,
    55430 => -52,
    55431 => -52,
    55432 => -52,
    55433 => -52,
    55434 => -52,
    55435 => -52,
    55436 => -52,
    55437 => -52,
    55438 => -52,
    55439 => -52,
    55440 => -52,
    55441 => -52,
    55442 => -52,
    55443 => -52,
    55444 => -52,
    55445 => -52,
    55446 => -52,
    55447 => -52,
    55448 => -52,
    55449 => -52,
    55450 => -52,
    55451 => -52,
    55452 => -52,
    55453 => -52,
    55454 => -52,
    55455 => -52,
    55456 => -52,
    55457 => -52,
    55458 => -52,
    55459 => -52,
    55460 => -52,
    55461 => -52,
    55462 => -52,
    55463 => -52,
    55464 => -52,
    55465 => -52,
    55466 => -52,
    55467 => -52,
    55468 => -52,
    55469 => -52,
    55470 => -52,
    55471 => -52,
    55472 => -52,
    55473 => -52,
    55474 => -52,
    55475 => -52,
    55476 => -52,
    55477 => -52,
    55478 => -52,
    55479 => -52,
    55480 => -52,
    55481 => -52,
    55482 => -52,
    55483 => -52,
    55484 => -52,
    55485 => -52,
    55486 => -52,
    55487 => -52,
    55488 => -52,
    55489 => -52,
    55490 => -52,
    55491 => -52,
    55492 => -52,
    55493 => -52,
    55494 => -52,
    55495 => -52,
    55496 => -52,
    55497 => -52,
    55498 => -52,
    55499 => -52,
    55500 => -52,
    55501 => -52,
    55502 => -52,
    55503 => -52,
    55504 => -52,
    55505 => -52,
    55506 => -52,
    55507 => -52,
    55508 => -52,
    55509 => -52,
    55510 => -52,
    55511 => -52,
    55512 => -52,
    55513 => -52,
    55514 => -52,
    55515 => -52,
    55516 => -52,
    55517 => -52,
    55518 => -52,
    55519 => -52,
    55520 => -52,
    55521 => -52,
    55522 => -52,
    55523 => -52,
    55524 => -52,
    55525 => -52,
    55526 => -52,
    55527 => -52,
    55528 => -52,
    55529 => -52,
    55530 => -52,
    55531 => -52,
    55532 => -52,
    55533 => -52,
    55534 => -52,
    55535 => -52,
    55536 => -52,
    55537 => -52,
    55538 => -52,
    55539 => -52,
    55540 => -52,
    55541 => -52,
    55542 => -52,
    55543 => -52,
    55544 => -52,
    55545 => -52,
    55546 => -52,
    55547 => -52,
    55548 => -52,
    55549 => -52,
    55550 => -52,
    55551 => -52,
    55552 => -52,
    55553 => -52,
    55554 => -52,
    55555 => -51,
    55556 => -51,
    55557 => -51,
    55558 => -51,
    55559 => -51,
    55560 => -51,
    55561 => -51,
    55562 => -51,
    55563 => -51,
    55564 => -51,
    55565 => -51,
    55566 => -51,
    55567 => -51,
    55568 => -51,
    55569 => -51,
    55570 => -51,
    55571 => -51,
    55572 => -51,
    55573 => -51,
    55574 => -51,
    55575 => -51,
    55576 => -51,
    55577 => -51,
    55578 => -51,
    55579 => -51,
    55580 => -51,
    55581 => -51,
    55582 => -51,
    55583 => -51,
    55584 => -51,
    55585 => -51,
    55586 => -51,
    55587 => -51,
    55588 => -51,
    55589 => -51,
    55590 => -51,
    55591 => -51,
    55592 => -51,
    55593 => -51,
    55594 => -51,
    55595 => -51,
    55596 => -51,
    55597 => -51,
    55598 => -51,
    55599 => -51,
    55600 => -51,
    55601 => -51,
    55602 => -51,
    55603 => -51,
    55604 => -51,
    55605 => -51,
    55606 => -51,
    55607 => -51,
    55608 => -51,
    55609 => -51,
    55610 => -51,
    55611 => -51,
    55612 => -51,
    55613 => -51,
    55614 => -51,
    55615 => -51,
    55616 => -51,
    55617 => -51,
    55618 => -51,
    55619 => -51,
    55620 => -51,
    55621 => -51,
    55622 => -51,
    55623 => -51,
    55624 => -51,
    55625 => -51,
    55626 => -51,
    55627 => -51,
    55628 => -51,
    55629 => -51,
    55630 => -51,
    55631 => -51,
    55632 => -51,
    55633 => -51,
    55634 => -51,
    55635 => -51,
    55636 => -51,
    55637 => -51,
    55638 => -51,
    55639 => -51,
    55640 => -51,
    55641 => -51,
    55642 => -51,
    55643 => -51,
    55644 => -51,
    55645 => -51,
    55646 => -51,
    55647 => -51,
    55648 => -51,
    55649 => -51,
    55650 => -51,
    55651 => -51,
    55652 => -51,
    55653 => -51,
    55654 => -51,
    55655 => -51,
    55656 => -51,
    55657 => -51,
    55658 => -51,
    55659 => -51,
    55660 => -51,
    55661 => -51,
    55662 => -51,
    55663 => -51,
    55664 => -51,
    55665 => -51,
    55666 => -51,
    55667 => -51,
    55668 => -51,
    55669 => -51,
    55670 => -51,
    55671 => -51,
    55672 => -51,
    55673 => -51,
    55674 => -51,
    55675 => -51,
    55676 => -51,
    55677 => -51,
    55678 => -51,
    55679 => -51,
    55680 => -51,
    55681 => -51,
    55682 => -51,
    55683 => -51,
    55684 => -51,
    55685 => -51,
    55686 => -51,
    55687 => -51,
    55688 => -51,
    55689 => -51,
    55690 => -51,
    55691 => -51,
    55692 => -51,
    55693 => -51,
    55694 => -51,
    55695 => -51,
    55696 => -51,
    55697 => -51,
    55698 => -51,
    55699 => -51,
    55700 => -51,
    55701 => -51,
    55702 => -51,
    55703 => -51,
    55704 => -51,
    55705 => -51,
    55706 => -51,
    55707 => -51,
    55708 => -51,
    55709 => -51,
    55710 => -51,
    55711 => -51,
    55712 => -51,
    55713 => -51,
    55714 => -51,
    55715 => -51,
    55716 => -51,
    55717 => -51,
    55718 => -51,
    55719 => -51,
    55720 => -51,
    55721 => -51,
    55722 => -51,
    55723 => -51,
    55724 => -51,
    55725 => -51,
    55726 => -51,
    55727 => -51,
    55728 => -51,
    55729 => -51,
    55730 => -51,
    55731 => -51,
    55732 => -51,
    55733 => -51,
    55734 => -51,
    55735 => -51,
    55736 => -51,
    55737 => -51,
    55738 => -51,
    55739 => -51,
    55740 => -51,
    55741 => -51,
    55742 => -51,
    55743 => -51,
    55744 => -51,
    55745 => -51,
    55746 => -51,
    55747 => -51,
    55748 => -51,
    55749 => -51,
    55750 => -51,
    55751 => -51,
    55752 => -51,
    55753 => -51,
    55754 => -51,
    55755 => -51,
    55756 => -51,
    55757 => -51,
    55758 => -51,
    55759 => -51,
    55760 => -51,
    55761 => -51,
    55762 => -51,
    55763 => -51,
    55764 => -51,
    55765 => -51,
    55766 => -51,
    55767 => -51,
    55768 => -51,
    55769 => -51,
    55770 => -51,
    55771 => -51,
    55772 => -51,
    55773 => -51,
    55774 => -51,
    55775 => -51,
    55776 => -51,
    55777 => -51,
    55778 => -51,
    55779 => -51,
    55780 => -51,
    55781 => -51,
    55782 => -51,
    55783 => -51,
    55784 => -51,
    55785 => -51,
    55786 => -51,
    55787 => -51,
    55788 => -51,
    55789 => -51,
    55790 => -51,
    55791 => -51,
    55792 => -51,
    55793 => -51,
    55794 => -51,
    55795 => -51,
    55796 => -51,
    55797 => -51,
    55798 => -51,
    55799 => -51,
    55800 => -51,
    55801 => -51,
    55802 => -51,
    55803 => -51,
    55804 => -51,
    55805 => -51,
    55806 => -51,
    55807 => -51,
    55808 => -51,
    55809 => -51,
    55810 => -51,
    55811 => -51,
    55812 => -51,
    55813 => -51,
    55814 => -51,
    55815 => -51,
    55816 => -51,
    55817 => -51,
    55818 => -51,
    55819 => -51,
    55820 => -51,
    55821 => -51,
    55822 => -51,
    55823 => -51,
    55824 => -51,
    55825 => -51,
    55826 => -51,
    55827 => -51,
    55828 => -51,
    55829 => -51,
    55830 => -51,
    55831 => -51,
    55832 => -51,
    55833 => -51,
    55834 => -51,
    55835 => -51,
    55836 => -51,
    55837 => -50,
    55838 => -50,
    55839 => -50,
    55840 => -50,
    55841 => -50,
    55842 => -50,
    55843 => -50,
    55844 => -50,
    55845 => -50,
    55846 => -50,
    55847 => -50,
    55848 => -50,
    55849 => -50,
    55850 => -50,
    55851 => -50,
    55852 => -50,
    55853 => -50,
    55854 => -50,
    55855 => -50,
    55856 => -50,
    55857 => -50,
    55858 => -50,
    55859 => -50,
    55860 => -50,
    55861 => -50,
    55862 => -50,
    55863 => -50,
    55864 => -50,
    55865 => -50,
    55866 => -50,
    55867 => -50,
    55868 => -50,
    55869 => -50,
    55870 => -50,
    55871 => -50,
    55872 => -50,
    55873 => -50,
    55874 => -50,
    55875 => -50,
    55876 => -50,
    55877 => -50,
    55878 => -50,
    55879 => -50,
    55880 => -50,
    55881 => -50,
    55882 => -50,
    55883 => -50,
    55884 => -50,
    55885 => -50,
    55886 => -50,
    55887 => -50,
    55888 => -50,
    55889 => -50,
    55890 => -50,
    55891 => -50,
    55892 => -50,
    55893 => -50,
    55894 => -50,
    55895 => -50,
    55896 => -50,
    55897 => -50,
    55898 => -50,
    55899 => -50,
    55900 => -50,
    55901 => -50,
    55902 => -50,
    55903 => -50,
    55904 => -50,
    55905 => -50,
    55906 => -50,
    55907 => -50,
    55908 => -50,
    55909 => -50,
    55910 => -50,
    55911 => -50,
    55912 => -50,
    55913 => -50,
    55914 => -50,
    55915 => -50,
    55916 => -50,
    55917 => -50,
    55918 => -50,
    55919 => -50,
    55920 => -50,
    55921 => -50,
    55922 => -50,
    55923 => -50,
    55924 => -50,
    55925 => -50,
    55926 => -50,
    55927 => -50,
    55928 => -50,
    55929 => -50,
    55930 => -50,
    55931 => -50,
    55932 => -50,
    55933 => -50,
    55934 => -50,
    55935 => -50,
    55936 => -50,
    55937 => -50,
    55938 => -50,
    55939 => -50,
    55940 => -50,
    55941 => -50,
    55942 => -50,
    55943 => -50,
    55944 => -50,
    55945 => -50,
    55946 => -50,
    55947 => -50,
    55948 => -50,
    55949 => -50,
    55950 => -50,
    55951 => -50,
    55952 => -50,
    55953 => -50,
    55954 => -50,
    55955 => -50,
    55956 => -50,
    55957 => -50,
    55958 => -50,
    55959 => -50,
    55960 => -50,
    55961 => -50,
    55962 => -50,
    55963 => -50,
    55964 => -50,
    55965 => -50,
    55966 => -50,
    55967 => -50,
    55968 => -50,
    55969 => -50,
    55970 => -50,
    55971 => -50,
    55972 => -50,
    55973 => -50,
    55974 => -50,
    55975 => -50,
    55976 => -50,
    55977 => -50,
    55978 => -50,
    55979 => -50,
    55980 => -50,
    55981 => -50,
    55982 => -50,
    55983 => -50,
    55984 => -50,
    55985 => -50,
    55986 => -50,
    55987 => -50,
    55988 => -50,
    55989 => -50,
    55990 => -50,
    55991 => -50,
    55992 => -50,
    55993 => -50,
    55994 => -50,
    55995 => -50,
    55996 => -50,
    55997 => -50,
    55998 => -50,
    55999 => -50,
    56000 => -50,
    56001 => -50,
    56002 => -50,
    56003 => -50,
    56004 => -50,
    56005 => -50,
    56006 => -50,
    56007 => -50,
    56008 => -50,
    56009 => -50,
    56010 => -50,
    56011 => -50,
    56012 => -50,
    56013 => -50,
    56014 => -50,
    56015 => -50,
    56016 => -50,
    56017 => -50,
    56018 => -50,
    56019 => -50,
    56020 => -50,
    56021 => -50,
    56022 => -50,
    56023 => -50,
    56024 => -50,
    56025 => -50,
    56026 => -50,
    56027 => -50,
    56028 => -50,
    56029 => -50,
    56030 => -50,
    56031 => -50,
    56032 => -50,
    56033 => -50,
    56034 => -50,
    56035 => -50,
    56036 => -50,
    56037 => -50,
    56038 => -50,
    56039 => -50,
    56040 => -50,
    56041 => -50,
    56042 => -50,
    56043 => -50,
    56044 => -50,
    56045 => -50,
    56046 => -50,
    56047 => -50,
    56048 => -50,
    56049 => -50,
    56050 => -50,
    56051 => -50,
    56052 => -50,
    56053 => -50,
    56054 => -50,
    56055 => -50,
    56056 => -50,
    56057 => -50,
    56058 => -50,
    56059 => -50,
    56060 => -50,
    56061 => -50,
    56062 => -50,
    56063 => -50,
    56064 => -50,
    56065 => -50,
    56066 => -50,
    56067 => -50,
    56068 => -50,
    56069 => -50,
    56070 => -50,
    56071 => -50,
    56072 => -50,
    56073 => -50,
    56074 => -50,
    56075 => -50,
    56076 => -50,
    56077 => -50,
    56078 => -50,
    56079 => -50,
    56080 => -50,
    56081 => -50,
    56082 => -50,
    56083 => -50,
    56084 => -50,
    56085 => -50,
    56086 => -50,
    56087 => -50,
    56088 => -50,
    56089 => -50,
    56090 => -50,
    56091 => -50,
    56092 => -50,
    56093 => -50,
    56094 => -50,
    56095 => -50,
    56096 => -50,
    56097 => -50,
    56098 => -50,
    56099 => -50,
    56100 => -50,
    56101 => -50,
    56102 => -50,
    56103 => -50,
    56104 => -50,
    56105 => -50,
    56106 => -50,
    56107 => -50,
    56108 => -50,
    56109 => -49,
    56110 => -49,
    56111 => -49,
    56112 => -49,
    56113 => -49,
    56114 => -49,
    56115 => -49,
    56116 => -49,
    56117 => -49,
    56118 => -49,
    56119 => -49,
    56120 => -49,
    56121 => -49,
    56122 => -49,
    56123 => -49,
    56124 => -49,
    56125 => -49,
    56126 => -49,
    56127 => -49,
    56128 => -49,
    56129 => -49,
    56130 => -49,
    56131 => -49,
    56132 => -49,
    56133 => -49,
    56134 => -49,
    56135 => -49,
    56136 => -49,
    56137 => -49,
    56138 => -49,
    56139 => -49,
    56140 => -49,
    56141 => -49,
    56142 => -49,
    56143 => -49,
    56144 => -49,
    56145 => -49,
    56146 => -49,
    56147 => -49,
    56148 => -49,
    56149 => -49,
    56150 => -49,
    56151 => -49,
    56152 => -49,
    56153 => -49,
    56154 => -49,
    56155 => -49,
    56156 => -49,
    56157 => -49,
    56158 => -49,
    56159 => -49,
    56160 => -49,
    56161 => -49,
    56162 => -49,
    56163 => -49,
    56164 => -49,
    56165 => -49,
    56166 => -49,
    56167 => -49,
    56168 => -49,
    56169 => -49,
    56170 => -49,
    56171 => -49,
    56172 => -49,
    56173 => -49,
    56174 => -49,
    56175 => -49,
    56176 => -49,
    56177 => -49,
    56178 => -49,
    56179 => -49,
    56180 => -49,
    56181 => -49,
    56182 => -49,
    56183 => -49,
    56184 => -49,
    56185 => -49,
    56186 => -49,
    56187 => -49,
    56188 => -49,
    56189 => -49,
    56190 => -49,
    56191 => -49,
    56192 => -49,
    56193 => -49,
    56194 => -49,
    56195 => -49,
    56196 => -49,
    56197 => -49,
    56198 => -49,
    56199 => -49,
    56200 => -49,
    56201 => -49,
    56202 => -49,
    56203 => -49,
    56204 => -49,
    56205 => -49,
    56206 => -49,
    56207 => -49,
    56208 => -49,
    56209 => -49,
    56210 => -49,
    56211 => -49,
    56212 => -49,
    56213 => -49,
    56214 => -49,
    56215 => -49,
    56216 => -49,
    56217 => -49,
    56218 => -49,
    56219 => -49,
    56220 => -49,
    56221 => -49,
    56222 => -49,
    56223 => -49,
    56224 => -49,
    56225 => -49,
    56226 => -49,
    56227 => -49,
    56228 => -49,
    56229 => -49,
    56230 => -49,
    56231 => -49,
    56232 => -49,
    56233 => -49,
    56234 => -49,
    56235 => -49,
    56236 => -49,
    56237 => -49,
    56238 => -49,
    56239 => -49,
    56240 => -49,
    56241 => -49,
    56242 => -49,
    56243 => -49,
    56244 => -49,
    56245 => -49,
    56246 => -49,
    56247 => -49,
    56248 => -49,
    56249 => -49,
    56250 => -49,
    56251 => -49,
    56252 => -49,
    56253 => -49,
    56254 => -49,
    56255 => -49,
    56256 => -49,
    56257 => -49,
    56258 => -49,
    56259 => -49,
    56260 => -49,
    56261 => -49,
    56262 => -49,
    56263 => -49,
    56264 => -49,
    56265 => -49,
    56266 => -49,
    56267 => -49,
    56268 => -49,
    56269 => -49,
    56270 => -49,
    56271 => -49,
    56272 => -49,
    56273 => -49,
    56274 => -49,
    56275 => -49,
    56276 => -49,
    56277 => -49,
    56278 => -49,
    56279 => -49,
    56280 => -49,
    56281 => -49,
    56282 => -49,
    56283 => -49,
    56284 => -49,
    56285 => -49,
    56286 => -49,
    56287 => -49,
    56288 => -49,
    56289 => -49,
    56290 => -49,
    56291 => -49,
    56292 => -49,
    56293 => -49,
    56294 => -49,
    56295 => -49,
    56296 => -49,
    56297 => -49,
    56298 => -49,
    56299 => -49,
    56300 => -49,
    56301 => -49,
    56302 => -49,
    56303 => -49,
    56304 => -49,
    56305 => -49,
    56306 => -49,
    56307 => -49,
    56308 => -49,
    56309 => -49,
    56310 => -49,
    56311 => -49,
    56312 => -49,
    56313 => -49,
    56314 => -49,
    56315 => -49,
    56316 => -49,
    56317 => -49,
    56318 => -49,
    56319 => -49,
    56320 => -49,
    56321 => -49,
    56322 => -49,
    56323 => -49,
    56324 => -49,
    56325 => -49,
    56326 => -49,
    56327 => -49,
    56328 => -49,
    56329 => -49,
    56330 => -49,
    56331 => -49,
    56332 => -49,
    56333 => -49,
    56334 => -49,
    56335 => -49,
    56336 => -49,
    56337 => -49,
    56338 => -49,
    56339 => -49,
    56340 => -49,
    56341 => -49,
    56342 => -49,
    56343 => -49,
    56344 => -49,
    56345 => -49,
    56346 => -49,
    56347 => -49,
    56348 => -49,
    56349 => -49,
    56350 => -49,
    56351 => -49,
    56352 => -49,
    56353 => -49,
    56354 => -49,
    56355 => -49,
    56356 => -49,
    56357 => -49,
    56358 => -49,
    56359 => -49,
    56360 => -49,
    56361 => -49,
    56362 => -49,
    56363 => -49,
    56364 => -49,
    56365 => -49,
    56366 => -49,
    56367 => -49,
    56368 => -49,
    56369 => -49,
    56370 => -49,
    56371 => -49,
    56372 => -48,
    56373 => -48,
    56374 => -48,
    56375 => -48,
    56376 => -48,
    56377 => -48,
    56378 => -48,
    56379 => -48,
    56380 => -48,
    56381 => -48,
    56382 => -48,
    56383 => -48,
    56384 => -48,
    56385 => -48,
    56386 => -48,
    56387 => -48,
    56388 => -48,
    56389 => -48,
    56390 => -48,
    56391 => -48,
    56392 => -48,
    56393 => -48,
    56394 => -48,
    56395 => -48,
    56396 => -48,
    56397 => -48,
    56398 => -48,
    56399 => -48,
    56400 => -48,
    56401 => -48,
    56402 => -48,
    56403 => -48,
    56404 => -48,
    56405 => -48,
    56406 => -48,
    56407 => -48,
    56408 => -48,
    56409 => -48,
    56410 => -48,
    56411 => -48,
    56412 => -48,
    56413 => -48,
    56414 => -48,
    56415 => -48,
    56416 => -48,
    56417 => -48,
    56418 => -48,
    56419 => -48,
    56420 => -48,
    56421 => -48,
    56422 => -48,
    56423 => -48,
    56424 => -48,
    56425 => -48,
    56426 => -48,
    56427 => -48,
    56428 => -48,
    56429 => -48,
    56430 => -48,
    56431 => -48,
    56432 => -48,
    56433 => -48,
    56434 => -48,
    56435 => -48,
    56436 => -48,
    56437 => -48,
    56438 => -48,
    56439 => -48,
    56440 => -48,
    56441 => -48,
    56442 => -48,
    56443 => -48,
    56444 => -48,
    56445 => -48,
    56446 => -48,
    56447 => -48,
    56448 => -48,
    56449 => -48,
    56450 => -48,
    56451 => -48,
    56452 => -48,
    56453 => -48,
    56454 => -48,
    56455 => -48,
    56456 => -48,
    56457 => -48,
    56458 => -48,
    56459 => -48,
    56460 => -48,
    56461 => -48,
    56462 => -48,
    56463 => -48,
    56464 => -48,
    56465 => -48,
    56466 => -48,
    56467 => -48,
    56468 => -48,
    56469 => -48,
    56470 => -48,
    56471 => -48,
    56472 => -48,
    56473 => -48,
    56474 => -48,
    56475 => -48,
    56476 => -48,
    56477 => -48,
    56478 => -48,
    56479 => -48,
    56480 => -48,
    56481 => -48,
    56482 => -48,
    56483 => -48,
    56484 => -48,
    56485 => -48,
    56486 => -48,
    56487 => -48,
    56488 => -48,
    56489 => -48,
    56490 => -48,
    56491 => -48,
    56492 => -48,
    56493 => -48,
    56494 => -48,
    56495 => -48,
    56496 => -48,
    56497 => -48,
    56498 => -48,
    56499 => -48,
    56500 => -48,
    56501 => -48,
    56502 => -48,
    56503 => -48,
    56504 => -48,
    56505 => -48,
    56506 => -48,
    56507 => -48,
    56508 => -48,
    56509 => -48,
    56510 => -48,
    56511 => -48,
    56512 => -48,
    56513 => -48,
    56514 => -48,
    56515 => -48,
    56516 => -48,
    56517 => -48,
    56518 => -48,
    56519 => -48,
    56520 => -48,
    56521 => -48,
    56522 => -48,
    56523 => -48,
    56524 => -48,
    56525 => -48,
    56526 => -48,
    56527 => -48,
    56528 => -48,
    56529 => -48,
    56530 => -48,
    56531 => -48,
    56532 => -48,
    56533 => -48,
    56534 => -48,
    56535 => -48,
    56536 => -48,
    56537 => -48,
    56538 => -48,
    56539 => -48,
    56540 => -48,
    56541 => -48,
    56542 => -48,
    56543 => -48,
    56544 => -48,
    56545 => -48,
    56546 => -48,
    56547 => -48,
    56548 => -48,
    56549 => -48,
    56550 => -48,
    56551 => -48,
    56552 => -48,
    56553 => -48,
    56554 => -48,
    56555 => -48,
    56556 => -48,
    56557 => -48,
    56558 => -48,
    56559 => -48,
    56560 => -48,
    56561 => -48,
    56562 => -48,
    56563 => -48,
    56564 => -48,
    56565 => -48,
    56566 => -48,
    56567 => -48,
    56568 => -48,
    56569 => -48,
    56570 => -48,
    56571 => -48,
    56572 => -48,
    56573 => -48,
    56574 => -48,
    56575 => -48,
    56576 => -48,
    56577 => -48,
    56578 => -48,
    56579 => -48,
    56580 => -48,
    56581 => -48,
    56582 => -48,
    56583 => -48,
    56584 => -48,
    56585 => -48,
    56586 => -48,
    56587 => -48,
    56588 => -48,
    56589 => -48,
    56590 => -48,
    56591 => -48,
    56592 => -48,
    56593 => -48,
    56594 => -48,
    56595 => -48,
    56596 => -48,
    56597 => -48,
    56598 => -48,
    56599 => -48,
    56600 => -48,
    56601 => -48,
    56602 => -48,
    56603 => -48,
    56604 => -48,
    56605 => -48,
    56606 => -48,
    56607 => -48,
    56608 => -48,
    56609 => -48,
    56610 => -48,
    56611 => -48,
    56612 => -48,
    56613 => -48,
    56614 => -48,
    56615 => -48,
    56616 => -48,
    56617 => -48,
    56618 => -48,
    56619 => -48,
    56620 => -48,
    56621 => -48,
    56622 => -48,
    56623 => -48,
    56624 => -48,
    56625 => -48,
    56626 => -48,
    56627 => -48,
    56628 => -47,
    56629 => -47,
    56630 => -47,
    56631 => -47,
    56632 => -47,
    56633 => -47,
    56634 => -47,
    56635 => -47,
    56636 => -47,
    56637 => -47,
    56638 => -47,
    56639 => -47,
    56640 => -47,
    56641 => -47,
    56642 => -47,
    56643 => -47,
    56644 => -47,
    56645 => -47,
    56646 => -47,
    56647 => -47,
    56648 => -47,
    56649 => -47,
    56650 => -47,
    56651 => -47,
    56652 => -47,
    56653 => -47,
    56654 => -47,
    56655 => -47,
    56656 => -47,
    56657 => -47,
    56658 => -47,
    56659 => -47,
    56660 => -47,
    56661 => -47,
    56662 => -47,
    56663 => -47,
    56664 => -47,
    56665 => -47,
    56666 => -47,
    56667 => -47,
    56668 => -47,
    56669 => -47,
    56670 => -47,
    56671 => -47,
    56672 => -47,
    56673 => -47,
    56674 => -47,
    56675 => -47,
    56676 => -47,
    56677 => -47,
    56678 => -47,
    56679 => -47,
    56680 => -47,
    56681 => -47,
    56682 => -47,
    56683 => -47,
    56684 => -47,
    56685 => -47,
    56686 => -47,
    56687 => -47,
    56688 => -47,
    56689 => -47,
    56690 => -47,
    56691 => -47,
    56692 => -47,
    56693 => -47,
    56694 => -47,
    56695 => -47,
    56696 => -47,
    56697 => -47,
    56698 => -47,
    56699 => -47,
    56700 => -47,
    56701 => -47,
    56702 => -47,
    56703 => -47,
    56704 => -47,
    56705 => -47,
    56706 => -47,
    56707 => -47,
    56708 => -47,
    56709 => -47,
    56710 => -47,
    56711 => -47,
    56712 => -47,
    56713 => -47,
    56714 => -47,
    56715 => -47,
    56716 => -47,
    56717 => -47,
    56718 => -47,
    56719 => -47,
    56720 => -47,
    56721 => -47,
    56722 => -47,
    56723 => -47,
    56724 => -47,
    56725 => -47,
    56726 => -47,
    56727 => -47,
    56728 => -47,
    56729 => -47,
    56730 => -47,
    56731 => -47,
    56732 => -47,
    56733 => -47,
    56734 => -47,
    56735 => -47,
    56736 => -47,
    56737 => -47,
    56738 => -47,
    56739 => -47,
    56740 => -47,
    56741 => -47,
    56742 => -47,
    56743 => -47,
    56744 => -47,
    56745 => -47,
    56746 => -47,
    56747 => -47,
    56748 => -47,
    56749 => -47,
    56750 => -47,
    56751 => -47,
    56752 => -47,
    56753 => -47,
    56754 => -47,
    56755 => -47,
    56756 => -47,
    56757 => -47,
    56758 => -47,
    56759 => -47,
    56760 => -47,
    56761 => -47,
    56762 => -47,
    56763 => -47,
    56764 => -47,
    56765 => -47,
    56766 => -47,
    56767 => -47,
    56768 => -47,
    56769 => -47,
    56770 => -47,
    56771 => -47,
    56772 => -47,
    56773 => -47,
    56774 => -47,
    56775 => -47,
    56776 => -47,
    56777 => -47,
    56778 => -47,
    56779 => -47,
    56780 => -47,
    56781 => -47,
    56782 => -47,
    56783 => -47,
    56784 => -47,
    56785 => -47,
    56786 => -47,
    56787 => -47,
    56788 => -47,
    56789 => -47,
    56790 => -47,
    56791 => -47,
    56792 => -47,
    56793 => -47,
    56794 => -47,
    56795 => -47,
    56796 => -47,
    56797 => -47,
    56798 => -47,
    56799 => -47,
    56800 => -47,
    56801 => -47,
    56802 => -47,
    56803 => -47,
    56804 => -47,
    56805 => -47,
    56806 => -47,
    56807 => -47,
    56808 => -47,
    56809 => -47,
    56810 => -47,
    56811 => -47,
    56812 => -47,
    56813 => -47,
    56814 => -47,
    56815 => -47,
    56816 => -47,
    56817 => -47,
    56818 => -47,
    56819 => -47,
    56820 => -47,
    56821 => -47,
    56822 => -47,
    56823 => -47,
    56824 => -47,
    56825 => -47,
    56826 => -47,
    56827 => -47,
    56828 => -47,
    56829 => -47,
    56830 => -47,
    56831 => -47,
    56832 => -47,
    56833 => -47,
    56834 => -47,
    56835 => -47,
    56836 => -47,
    56837 => -47,
    56838 => -47,
    56839 => -47,
    56840 => -47,
    56841 => -47,
    56842 => -47,
    56843 => -47,
    56844 => -47,
    56845 => -47,
    56846 => -47,
    56847 => -47,
    56848 => -47,
    56849 => -47,
    56850 => -47,
    56851 => -47,
    56852 => -47,
    56853 => -47,
    56854 => -47,
    56855 => -47,
    56856 => -47,
    56857 => -47,
    56858 => -47,
    56859 => -47,
    56860 => -47,
    56861 => -47,
    56862 => -47,
    56863 => -47,
    56864 => -47,
    56865 => -47,
    56866 => -47,
    56867 => -47,
    56868 => -47,
    56869 => -47,
    56870 => -47,
    56871 => -47,
    56872 => -47,
    56873 => -47,
    56874 => -47,
    56875 => -47,
    56876 => -47,
    56877 => -46,
    56878 => -46,
    56879 => -46,
    56880 => -46,
    56881 => -46,
    56882 => -46,
    56883 => -46,
    56884 => -46,
    56885 => -46,
    56886 => -46,
    56887 => -46,
    56888 => -46,
    56889 => -46,
    56890 => -46,
    56891 => -46,
    56892 => -46,
    56893 => -46,
    56894 => -46,
    56895 => -46,
    56896 => -46,
    56897 => -46,
    56898 => -46,
    56899 => -46,
    56900 => -46,
    56901 => -46,
    56902 => -46,
    56903 => -46,
    56904 => -46,
    56905 => -46,
    56906 => -46,
    56907 => -46,
    56908 => -46,
    56909 => -46,
    56910 => -46,
    56911 => -46,
    56912 => -46,
    56913 => -46,
    56914 => -46,
    56915 => -46,
    56916 => -46,
    56917 => -46,
    56918 => -46,
    56919 => -46,
    56920 => -46,
    56921 => -46,
    56922 => -46,
    56923 => -46,
    56924 => -46,
    56925 => -46,
    56926 => -46,
    56927 => -46,
    56928 => -46,
    56929 => -46,
    56930 => -46,
    56931 => -46,
    56932 => -46,
    56933 => -46,
    56934 => -46,
    56935 => -46,
    56936 => -46,
    56937 => -46,
    56938 => -46,
    56939 => -46,
    56940 => -46,
    56941 => -46,
    56942 => -46,
    56943 => -46,
    56944 => -46,
    56945 => -46,
    56946 => -46,
    56947 => -46,
    56948 => -46,
    56949 => -46,
    56950 => -46,
    56951 => -46,
    56952 => -46,
    56953 => -46,
    56954 => -46,
    56955 => -46,
    56956 => -46,
    56957 => -46,
    56958 => -46,
    56959 => -46,
    56960 => -46,
    56961 => -46,
    56962 => -46,
    56963 => -46,
    56964 => -46,
    56965 => -46,
    56966 => -46,
    56967 => -46,
    56968 => -46,
    56969 => -46,
    56970 => -46,
    56971 => -46,
    56972 => -46,
    56973 => -46,
    56974 => -46,
    56975 => -46,
    56976 => -46,
    56977 => -46,
    56978 => -46,
    56979 => -46,
    56980 => -46,
    56981 => -46,
    56982 => -46,
    56983 => -46,
    56984 => -46,
    56985 => -46,
    56986 => -46,
    56987 => -46,
    56988 => -46,
    56989 => -46,
    56990 => -46,
    56991 => -46,
    56992 => -46,
    56993 => -46,
    56994 => -46,
    56995 => -46,
    56996 => -46,
    56997 => -46,
    56998 => -46,
    56999 => -46,
    57000 => -46,
    57001 => -46,
    57002 => -46,
    57003 => -46,
    57004 => -46,
    57005 => -46,
    57006 => -46,
    57007 => -46,
    57008 => -46,
    57009 => -46,
    57010 => -46,
    57011 => -46,
    57012 => -46,
    57013 => -46,
    57014 => -46,
    57015 => -46,
    57016 => -46,
    57017 => -46,
    57018 => -46,
    57019 => -46,
    57020 => -46,
    57021 => -46,
    57022 => -46,
    57023 => -46,
    57024 => -46,
    57025 => -46,
    57026 => -46,
    57027 => -46,
    57028 => -46,
    57029 => -46,
    57030 => -46,
    57031 => -46,
    57032 => -46,
    57033 => -46,
    57034 => -46,
    57035 => -46,
    57036 => -46,
    57037 => -46,
    57038 => -46,
    57039 => -46,
    57040 => -46,
    57041 => -46,
    57042 => -46,
    57043 => -46,
    57044 => -46,
    57045 => -46,
    57046 => -46,
    57047 => -46,
    57048 => -46,
    57049 => -46,
    57050 => -46,
    57051 => -46,
    57052 => -46,
    57053 => -46,
    57054 => -46,
    57055 => -46,
    57056 => -46,
    57057 => -46,
    57058 => -46,
    57059 => -46,
    57060 => -46,
    57061 => -46,
    57062 => -46,
    57063 => -46,
    57064 => -46,
    57065 => -46,
    57066 => -46,
    57067 => -46,
    57068 => -46,
    57069 => -46,
    57070 => -46,
    57071 => -46,
    57072 => -46,
    57073 => -46,
    57074 => -46,
    57075 => -46,
    57076 => -46,
    57077 => -46,
    57078 => -46,
    57079 => -46,
    57080 => -46,
    57081 => -46,
    57082 => -46,
    57083 => -46,
    57084 => -46,
    57085 => -46,
    57086 => -46,
    57087 => -46,
    57088 => -46,
    57089 => -46,
    57090 => -46,
    57091 => -46,
    57092 => -46,
    57093 => -46,
    57094 => -46,
    57095 => -46,
    57096 => -46,
    57097 => -46,
    57098 => -46,
    57099 => -46,
    57100 => -46,
    57101 => -46,
    57102 => -46,
    57103 => -46,
    57104 => -46,
    57105 => -46,
    57106 => -46,
    57107 => -46,
    57108 => -46,
    57109 => -46,
    57110 => -46,
    57111 => -46,
    57112 => -46,
    57113 => -46,
    57114 => -46,
    57115 => -46,
    57116 => -46,
    57117 => -46,
    57118 => -46,
    57119 => -45,
    57120 => -45,
    57121 => -45,
    57122 => -45,
    57123 => -45,
    57124 => -45,
    57125 => -45,
    57126 => -45,
    57127 => -45,
    57128 => -45,
    57129 => -45,
    57130 => -45,
    57131 => -45,
    57132 => -45,
    57133 => -45,
    57134 => -45,
    57135 => -45,
    57136 => -45,
    57137 => -45,
    57138 => -45,
    57139 => -45,
    57140 => -45,
    57141 => -45,
    57142 => -45,
    57143 => -45,
    57144 => -45,
    57145 => -45,
    57146 => -45,
    57147 => -45,
    57148 => -45,
    57149 => -45,
    57150 => -45,
    57151 => -45,
    57152 => -45,
    57153 => -45,
    57154 => -45,
    57155 => -45,
    57156 => -45,
    57157 => -45,
    57158 => -45,
    57159 => -45,
    57160 => -45,
    57161 => -45,
    57162 => -45,
    57163 => -45,
    57164 => -45,
    57165 => -45,
    57166 => -45,
    57167 => -45,
    57168 => -45,
    57169 => -45,
    57170 => -45,
    57171 => -45,
    57172 => -45,
    57173 => -45,
    57174 => -45,
    57175 => -45,
    57176 => -45,
    57177 => -45,
    57178 => -45,
    57179 => -45,
    57180 => -45,
    57181 => -45,
    57182 => -45,
    57183 => -45,
    57184 => -45,
    57185 => -45,
    57186 => -45,
    57187 => -45,
    57188 => -45,
    57189 => -45,
    57190 => -45,
    57191 => -45,
    57192 => -45,
    57193 => -45,
    57194 => -45,
    57195 => -45,
    57196 => -45,
    57197 => -45,
    57198 => -45,
    57199 => -45,
    57200 => -45,
    57201 => -45,
    57202 => -45,
    57203 => -45,
    57204 => -45,
    57205 => -45,
    57206 => -45,
    57207 => -45,
    57208 => -45,
    57209 => -45,
    57210 => -45,
    57211 => -45,
    57212 => -45,
    57213 => -45,
    57214 => -45,
    57215 => -45,
    57216 => -45,
    57217 => -45,
    57218 => -45,
    57219 => -45,
    57220 => -45,
    57221 => -45,
    57222 => -45,
    57223 => -45,
    57224 => -45,
    57225 => -45,
    57226 => -45,
    57227 => -45,
    57228 => -45,
    57229 => -45,
    57230 => -45,
    57231 => -45,
    57232 => -45,
    57233 => -45,
    57234 => -45,
    57235 => -45,
    57236 => -45,
    57237 => -45,
    57238 => -45,
    57239 => -45,
    57240 => -45,
    57241 => -45,
    57242 => -45,
    57243 => -45,
    57244 => -45,
    57245 => -45,
    57246 => -45,
    57247 => -45,
    57248 => -45,
    57249 => -45,
    57250 => -45,
    57251 => -45,
    57252 => -45,
    57253 => -45,
    57254 => -45,
    57255 => -45,
    57256 => -45,
    57257 => -45,
    57258 => -45,
    57259 => -45,
    57260 => -45,
    57261 => -45,
    57262 => -45,
    57263 => -45,
    57264 => -45,
    57265 => -45,
    57266 => -45,
    57267 => -45,
    57268 => -45,
    57269 => -45,
    57270 => -45,
    57271 => -45,
    57272 => -45,
    57273 => -45,
    57274 => -45,
    57275 => -45,
    57276 => -45,
    57277 => -45,
    57278 => -45,
    57279 => -45,
    57280 => -45,
    57281 => -45,
    57282 => -45,
    57283 => -45,
    57284 => -45,
    57285 => -45,
    57286 => -45,
    57287 => -45,
    57288 => -45,
    57289 => -45,
    57290 => -45,
    57291 => -45,
    57292 => -45,
    57293 => -45,
    57294 => -45,
    57295 => -45,
    57296 => -45,
    57297 => -45,
    57298 => -45,
    57299 => -45,
    57300 => -45,
    57301 => -45,
    57302 => -45,
    57303 => -45,
    57304 => -45,
    57305 => -45,
    57306 => -45,
    57307 => -45,
    57308 => -45,
    57309 => -45,
    57310 => -45,
    57311 => -45,
    57312 => -45,
    57313 => -45,
    57314 => -45,
    57315 => -45,
    57316 => -45,
    57317 => -45,
    57318 => -45,
    57319 => -45,
    57320 => -45,
    57321 => -45,
    57322 => -45,
    57323 => -45,
    57324 => -45,
    57325 => -45,
    57326 => -45,
    57327 => -45,
    57328 => -45,
    57329 => -45,
    57330 => -45,
    57331 => -45,
    57332 => -45,
    57333 => -45,
    57334 => -45,
    57335 => -45,
    57336 => -45,
    57337 => -45,
    57338 => -45,
    57339 => -45,
    57340 => -45,
    57341 => -45,
    57342 => -45,
    57343 => -45,
    57344 => -45,
    57345 => -45,
    57346 => -45,
    57347 => -45,
    57348 => -45,
    57349 => -45,
    57350 => -45,
    57351 => -45,
    57352 => -45,
    57353 => -45,
    57354 => -45,
    57355 => -45,
    57356 => -44,
    57357 => -44,
    57358 => -44,
    57359 => -44,
    57360 => -44,
    57361 => -44,
    57362 => -44,
    57363 => -44,
    57364 => -44,
    57365 => -44,
    57366 => -44,
    57367 => -44,
    57368 => -44,
    57369 => -44,
    57370 => -44,
    57371 => -44,
    57372 => -44,
    57373 => -44,
    57374 => -44,
    57375 => -44,
    57376 => -44,
    57377 => -44,
    57378 => -44,
    57379 => -44,
    57380 => -44,
    57381 => -44,
    57382 => -44,
    57383 => -44,
    57384 => -44,
    57385 => -44,
    57386 => -44,
    57387 => -44,
    57388 => -44,
    57389 => -44,
    57390 => -44,
    57391 => -44,
    57392 => -44,
    57393 => -44,
    57394 => -44,
    57395 => -44,
    57396 => -44,
    57397 => -44,
    57398 => -44,
    57399 => -44,
    57400 => -44,
    57401 => -44,
    57402 => -44,
    57403 => -44,
    57404 => -44,
    57405 => -44,
    57406 => -44,
    57407 => -44,
    57408 => -44,
    57409 => -44,
    57410 => -44,
    57411 => -44,
    57412 => -44,
    57413 => -44,
    57414 => -44,
    57415 => -44,
    57416 => -44,
    57417 => -44,
    57418 => -44,
    57419 => -44,
    57420 => -44,
    57421 => -44,
    57422 => -44,
    57423 => -44,
    57424 => -44,
    57425 => -44,
    57426 => -44,
    57427 => -44,
    57428 => -44,
    57429 => -44,
    57430 => -44,
    57431 => -44,
    57432 => -44,
    57433 => -44,
    57434 => -44,
    57435 => -44,
    57436 => -44,
    57437 => -44,
    57438 => -44,
    57439 => -44,
    57440 => -44,
    57441 => -44,
    57442 => -44,
    57443 => -44,
    57444 => -44,
    57445 => -44,
    57446 => -44,
    57447 => -44,
    57448 => -44,
    57449 => -44,
    57450 => -44,
    57451 => -44,
    57452 => -44,
    57453 => -44,
    57454 => -44,
    57455 => -44,
    57456 => -44,
    57457 => -44,
    57458 => -44,
    57459 => -44,
    57460 => -44,
    57461 => -44,
    57462 => -44,
    57463 => -44,
    57464 => -44,
    57465 => -44,
    57466 => -44,
    57467 => -44,
    57468 => -44,
    57469 => -44,
    57470 => -44,
    57471 => -44,
    57472 => -44,
    57473 => -44,
    57474 => -44,
    57475 => -44,
    57476 => -44,
    57477 => -44,
    57478 => -44,
    57479 => -44,
    57480 => -44,
    57481 => -44,
    57482 => -44,
    57483 => -44,
    57484 => -44,
    57485 => -44,
    57486 => -44,
    57487 => -44,
    57488 => -44,
    57489 => -44,
    57490 => -44,
    57491 => -44,
    57492 => -44,
    57493 => -44,
    57494 => -44,
    57495 => -44,
    57496 => -44,
    57497 => -44,
    57498 => -44,
    57499 => -44,
    57500 => -44,
    57501 => -44,
    57502 => -44,
    57503 => -44,
    57504 => -44,
    57505 => -44,
    57506 => -44,
    57507 => -44,
    57508 => -44,
    57509 => -44,
    57510 => -44,
    57511 => -44,
    57512 => -44,
    57513 => -44,
    57514 => -44,
    57515 => -44,
    57516 => -44,
    57517 => -44,
    57518 => -44,
    57519 => -44,
    57520 => -44,
    57521 => -44,
    57522 => -44,
    57523 => -44,
    57524 => -44,
    57525 => -44,
    57526 => -44,
    57527 => -44,
    57528 => -44,
    57529 => -44,
    57530 => -44,
    57531 => -44,
    57532 => -44,
    57533 => -44,
    57534 => -44,
    57535 => -44,
    57536 => -44,
    57537 => -44,
    57538 => -44,
    57539 => -44,
    57540 => -44,
    57541 => -44,
    57542 => -44,
    57543 => -44,
    57544 => -44,
    57545 => -44,
    57546 => -44,
    57547 => -44,
    57548 => -44,
    57549 => -44,
    57550 => -44,
    57551 => -44,
    57552 => -44,
    57553 => -44,
    57554 => -44,
    57555 => -44,
    57556 => -44,
    57557 => -44,
    57558 => -44,
    57559 => -44,
    57560 => -44,
    57561 => -44,
    57562 => -44,
    57563 => -44,
    57564 => -44,
    57565 => -44,
    57566 => -44,
    57567 => -44,
    57568 => -44,
    57569 => -44,
    57570 => -44,
    57571 => -44,
    57572 => -44,
    57573 => -44,
    57574 => -44,
    57575 => -44,
    57576 => -44,
    57577 => -44,
    57578 => -44,
    57579 => -44,
    57580 => -44,
    57581 => -44,
    57582 => -44,
    57583 => -44,
    57584 => -44,
    57585 => -44,
    57586 => -44,
    57587 => -43,
    57588 => -43,
    57589 => -43,
    57590 => -43,
    57591 => -43,
    57592 => -43,
    57593 => -43,
    57594 => -43,
    57595 => -43,
    57596 => -43,
    57597 => -43,
    57598 => -43,
    57599 => -43,
    57600 => -43,
    57601 => -43,
    57602 => -43,
    57603 => -43,
    57604 => -43,
    57605 => -43,
    57606 => -43,
    57607 => -43,
    57608 => -43,
    57609 => -43,
    57610 => -43,
    57611 => -43,
    57612 => -43,
    57613 => -43,
    57614 => -43,
    57615 => -43,
    57616 => -43,
    57617 => -43,
    57618 => -43,
    57619 => -43,
    57620 => -43,
    57621 => -43,
    57622 => -43,
    57623 => -43,
    57624 => -43,
    57625 => -43,
    57626 => -43,
    57627 => -43,
    57628 => -43,
    57629 => -43,
    57630 => -43,
    57631 => -43,
    57632 => -43,
    57633 => -43,
    57634 => -43,
    57635 => -43,
    57636 => -43,
    57637 => -43,
    57638 => -43,
    57639 => -43,
    57640 => -43,
    57641 => -43,
    57642 => -43,
    57643 => -43,
    57644 => -43,
    57645 => -43,
    57646 => -43,
    57647 => -43,
    57648 => -43,
    57649 => -43,
    57650 => -43,
    57651 => -43,
    57652 => -43,
    57653 => -43,
    57654 => -43,
    57655 => -43,
    57656 => -43,
    57657 => -43,
    57658 => -43,
    57659 => -43,
    57660 => -43,
    57661 => -43,
    57662 => -43,
    57663 => -43,
    57664 => -43,
    57665 => -43,
    57666 => -43,
    57667 => -43,
    57668 => -43,
    57669 => -43,
    57670 => -43,
    57671 => -43,
    57672 => -43,
    57673 => -43,
    57674 => -43,
    57675 => -43,
    57676 => -43,
    57677 => -43,
    57678 => -43,
    57679 => -43,
    57680 => -43,
    57681 => -43,
    57682 => -43,
    57683 => -43,
    57684 => -43,
    57685 => -43,
    57686 => -43,
    57687 => -43,
    57688 => -43,
    57689 => -43,
    57690 => -43,
    57691 => -43,
    57692 => -43,
    57693 => -43,
    57694 => -43,
    57695 => -43,
    57696 => -43,
    57697 => -43,
    57698 => -43,
    57699 => -43,
    57700 => -43,
    57701 => -43,
    57702 => -43,
    57703 => -43,
    57704 => -43,
    57705 => -43,
    57706 => -43,
    57707 => -43,
    57708 => -43,
    57709 => -43,
    57710 => -43,
    57711 => -43,
    57712 => -43,
    57713 => -43,
    57714 => -43,
    57715 => -43,
    57716 => -43,
    57717 => -43,
    57718 => -43,
    57719 => -43,
    57720 => -43,
    57721 => -43,
    57722 => -43,
    57723 => -43,
    57724 => -43,
    57725 => -43,
    57726 => -43,
    57727 => -43,
    57728 => -43,
    57729 => -43,
    57730 => -43,
    57731 => -43,
    57732 => -43,
    57733 => -43,
    57734 => -43,
    57735 => -43,
    57736 => -43,
    57737 => -43,
    57738 => -43,
    57739 => -43,
    57740 => -43,
    57741 => -43,
    57742 => -43,
    57743 => -43,
    57744 => -43,
    57745 => -43,
    57746 => -43,
    57747 => -43,
    57748 => -43,
    57749 => -43,
    57750 => -43,
    57751 => -43,
    57752 => -43,
    57753 => -43,
    57754 => -43,
    57755 => -43,
    57756 => -43,
    57757 => -43,
    57758 => -43,
    57759 => -43,
    57760 => -43,
    57761 => -43,
    57762 => -43,
    57763 => -43,
    57764 => -43,
    57765 => -43,
    57766 => -43,
    57767 => -43,
    57768 => -43,
    57769 => -43,
    57770 => -43,
    57771 => -43,
    57772 => -43,
    57773 => -43,
    57774 => -43,
    57775 => -43,
    57776 => -43,
    57777 => -43,
    57778 => -43,
    57779 => -43,
    57780 => -43,
    57781 => -43,
    57782 => -43,
    57783 => -43,
    57784 => -43,
    57785 => -43,
    57786 => -43,
    57787 => -43,
    57788 => -43,
    57789 => -43,
    57790 => -43,
    57791 => -43,
    57792 => -43,
    57793 => -43,
    57794 => -43,
    57795 => -43,
    57796 => -43,
    57797 => -43,
    57798 => -43,
    57799 => -43,
    57800 => -43,
    57801 => -43,
    57802 => -43,
    57803 => -43,
    57804 => -43,
    57805 => -43,
    57806 => -43,
    57807 => -43,
    57808 => -43,
    57809 => -43,
    57810 => -43,
    57811 => -43,
    57812 => -43,
    57813 => -43,
    57814 => -42,
    57815 => -42,
    57816 => -42,
    57817 => -42,
    57818 => -42,
    57819 => -42,
    57820 => -42,
    57821 => -42,
    57822 => -42,
    57823 => -42,
    57824 => -42,
    57825 => -42,
    57826 => -42,
    57827 => -42,
    57828 => -42,
    57829 => -42,
    57830 => -42,
    57831 => -42,
    57832 => -42,
    57833 => -42,
    57834 => -42,
    57835 => -42,
    57836 => -42,
    57837 => -42,
    57838 => -42,
    57839 => -42,
    57840 => -42,
    57841 => -42,
    57842 => -42,
    57843 => -42,
    57844 => -42,
    57845 => -42,
    57846 => -42,
    57847 => -42,
    57848 => -42,
    57849 => -42,
    57850 => -42,
    57851 => -42,
    57852 => -42,
    57853 => -42,
    57854 => -42,
    57855 => -42,
    57856 => -42,
    57857 => -42,
    57858 => -42,
    57859 => -42,
    57860 => -42,
    57861 => -42,
    57862 => -42,
    57863 => -42,
    57864 => -42,
    57865 => -42,
    57866 => -42,
    57867 => -42,
    57868 => -42,
    57869 => -42,
    57870 => -42,
    57871 => -42,
    57872 => -42,
    57873 => -42,
    57874 => -42,
    57875 => -42,
    57876 => -42,
    57877 => -42,
    57878 => -42,
    57879 => -42,
    57880 => -42,
    57881 => -42,
    57882 => -42,
    57883 => -42,
    57884 => -42,
    57885 => -42,
    57886 => -42,
    57887 => -42,
    57888 => -42,
    57889 => -42,
    57890 => -42,
    57891 => -42,
    57892 => -42,
    57893 => -42,
    57894 => -42,
    57895 => -42,
    57896 => -42,
    57897 => -42,
    57898 => -42,
    57899 => -42,
    57900 => -42,
    57901 => -42,
    57902 => -42,
    57903 => -42,
    57904 => -42,
    57905 => -42,
    57906 => -42,
    57907 => -42,
    57908 => -42,
    57909 => -42,
    57910 => -42,
    57911 => -42,
    57912 => -42,
    57913 => -42,
    57914 => -42,
    57915 => -42,
    57916 => -42,
    57917 => -42,
    57918 => -42,
    57919 => -42,
    57920 => -42,
    57921 => -42,
    57922 => -42,
    57923 => -42,
    57924 => -42,
    57925 => -42,
    57926 => -42,
    57927 => -42,
    57928 => -42,
    57929 => -42,
    57930 => -42,
    57931 => -42,
    57932 => -42,
    57933 => -42,
    57934 => -42,
    57935 => -42,
    57936 => -42,
    57937 => -42,
    57938 => -42,
    57939 => -42,
    57940 => -42,
    57941 => -42,
    57942 => -42,
    57943 => -42,
    57944 => -42,
    57945 => -42,
    57946 => -42,
    57947 => -42,
    57948 => -42,
    57949 => -42,
    57950 => -42,
    57951 => -42,
    57952 => -42,
    57953 => -42,
    57954 => -42,
    57955 => -42,
    57956 => -42,
    57957 => -42,
    57958 => -42,
    57959 => -42,
    57960 => -42,
    57961 => -42,
    57962 => -42,
    57963 => -42,
    57964 => -42,
    57965 => -42,
    57966 => -42,
    57967 => -42,
    57968 => -42,
    57969 => -42,
    57970 => -42,
    57971 => -42,
    57972 => -42,
    57973 => -42,
    57974 => -42,
    57975 => -42,
    57976 => -42,
    57977 => -42,
    57978 => -42,
    57979 => -42,
    57980 => -42,
    57981 => -42,
    57982 => -42,
    57983 => -42,
    57984 => -42,
    57985 => -42,
    57986 => -42,
    57987 => -42,
    57988 => -42,
    57989 => -42,
    57990 => -42,
    57991 => -42,
    57992 => -42,
    57993 => -42,
    57994 => -42,
    57995 => -42,
    57996 => -42,
    57997 => -42,
    57998 => -42,
    57999 => -42,
    58000 => -42,
    58001 => -42,
    58002 => -42,
    58003 => -42,
    58004 => -42,
    58005 => -42,
    58006 => -42,
    58007 => -42,
    58008 => -42,
    58009 => -42,
    58010 => -42,
    58011 => -42,
    58012 => -42,
    58013 => -42,
    58014 => -42,
    58015 => -42,
    58016 => -42,
    58017 => -42,
    58018 => -42,
    58019 => -42,
    58020 => -42,
    58021 => -42,
    58022 => -42,
    58023 => -42,
    58024 => -42,
    58025 => -42,
    58026 => -42,
    58027 => -42,
    58028 => -42,
    58029 => -42,
    58030 => -42,
    58031 => -42,
    58032 => -42,
    58033 => -42,
    58034 => -42,
    58035 => -42,
    58036 => -41,
    58037 => -41,
    58038 => -41,
    58039 => -41,
    58040 => -41,
    58041 => -41,
    58042 => -41,
    58043 => -41,
    58044 => -41,
    58045 => -41,
    58046 => -41,
    58047 => -41,
    58048 => -41,
    58049 => -41,
    58050 => -41,
    58051 => -41,
    58052 => -41,
    58053 => -41,
    58054 => -41,
    58055 => -41,
    58056 => -41,
    58057 => -41,
    58058 => -41,
    58059 => -41,
    58060 => -41,
    58061 => -41,
    58062 => -41,
    58063 => -41,
    58064 => -41,
    58065 => -41,
    58066 => -41,
    58067 => -41,
    58068 => -41,
    58069 => -41,
    58070 => -41,
    58071 => -41,
    58072 => -41,
    58073 => -41,
    58074 => -41,
    58075 => -41,
    58076 => -41,
    58077 => -41,
    58078 => -41,
    58079 => -41,
    58080 => -41,
    58081 => -41,
    58082 => -41,
    58083 => -41,
    58084 => -41,
    58085 => -41,
    58086 => -41,
    58087 => -41,
    58088 => -41,
    58089 => -41,
    58090 => -41,
    58091 => -41,
    58092 => -41,
    58093 => -41,
    58094 => -41,
    58095 => -41,
    58096 => -41,
    58097 => -41,
    58098 => -41,
    58099 => -41,
    58100 => -41,
    58101 => -41,
    58102 => -41,
    58103 => -41,
    58104 => -41,
    58105 => -41,
    58106 => -41,
    58107 => -41,
    58108 => -41,
    58109 => -41,
    58110 => -41,
    58111 => -41,
    58112 => -41,
    58113 => -41,
    58114 => -41,
    58115 => -41,
    58116 => -41,
    58117 => -41,
    58118 => -41,
    58119 => -41,
    58120 => -41,
    58121 => -41,
    58122 => -41,
    58123 => -41,
    58124 => -41,
    58125 => -41,
    58126 => -41,
    58127 => -41,
    58128 => -41,
    58129 => -41,
    58130 => -41,
    58131 => -41,
    58132 => -41,
    58133 => -41,
    58134 => -41,
    58135 => -41,
    58136 => -41,
    58137 => -41,
    58138 => -41,
    58139 => -41,
    58140 => -41,
    58141 => -41,
    58142 => -41,
    58143 => -41,
    58144 => -41,
    58145 => -41,
    58146 => -41,
    58147 => -41,
    58148 => -41,
    58149 => -41,
    58150 => -41,
    58151 => -41,
    58152 => -41,
    58153 => -41,
    58154 => -41,
    58155 => -41,
    58156 => -41,
    58157 => -41,
    58158 => -41,
    58159 => -41,
    58160 => -41,
    58161 => -41,
    58162 => -41,
    58163 => -41,
    58164 => -41,
    58165 => -41,
    58166 => -41,
    58167 => -41,
    58168 => -41,
    58169 => -41,
    58170 => -41,
    58171 => -41,
    58172 => -41,
    58173 => -41,
    58174 => -41,
    58175 => -41,
    58176 => -41,
    58177 => -41,
    58178 => -41,
    58179 => -41,
    58180 => -41,
    58181 => -41,
    58182 => -41,
    58183 => -41,
    58184 => -41,
    58185 => -41,
    58186 => -41,
    58187 => -41,
    58188 => -41,
    58189 => -41,
    58190 => -41,
    58191 => -41,
    58192 => -41,
    58193 => -41,
    58194 => -41,
    58195 => -41,
    58196 => -41,
    58197 => -41,
    58198 => -41,
    58199 => -41,
    58200 => -41,
    58201 => -41,
    58202 => -41,
    58203 => -41,
    58204 => -41,
    58205 => -41,
    58206 => -41,
    58207 => -41,
    58208 => -41,
    58209 => -41,
    58210 => -41,
    58211 => -41,
    58212 => -41,
    58213 => -41,
    58214 => -41,
    58215 => -41,
    58216 => -41,
    58217 => -41,
    58218 => -41,
    58219 => -41,
    58220 => -41,
    58221 => -41,
    58222 => -41,
    58223 => -41,
    58224 => -41,
    58225 => -41,
    58226 => -41,
    58227 => -41,
    58228 => -41,
    58229 => -41,
    58230 => -41,
    58231 => -41,
    58232 => -41,
    58233 => -41,
    58234 => -41,
    58235 => -41,
    58236 => -41,
    58237 => -41,
    58238 => -41,
    58239 => -41,
    58240 => -41,
    58241 => -41,
    58242 => -41,
    58243 => -41,
    58244 => -41,
    58245 => -41,
    58246 => -41,
    58247 => -41,
    58248 => -41,
    58249 => -41,
    58250 => -41,
    58251 => -41,
    58252 => -41,
    58253 => -41,
    58254 => -40,
    58255 => -40,
    58256 => -40,
    58257 => -40,
    58258 => -40,
    58259 => -40,
    58260 => -40,
    58261 => -40,
    58262 => -40,
    58263 => -40,
    58264 => -40,
    58265 => -40,
    58266 => -40,
    58267 => -40,
    58268 => -40,
    58269 => -40,
    58270 => -40,
    58271 => -40,
    58272 => -40,
    58273 => -40,
    58274 => -40,
    58275 => -40,
    58276 => -40,
    58277 => -40,
    58278 => -40,
    58279 => -40,
    58280 => -40,
    58281 => -40,
    58282 => -40,
    58283 => -40,
    58284 => -40,
    58285 => -40,
    58286 => -40,
    58287 => -40,
    58288 => -40,
    58289 => -40,
    58290 => -40,
    58291 => -40,
    58292 => -40,
    58293 => -40,
    58294 => -40,
    58295 => -40,
    58296 => -40,
    58297 => -40,
    58298 => -40,
    58299 => -40,
    58300 => -40,
    58301 => -40,
    58302 => -40,
    58303 => -40,
    58304 => -40,
    58305 => -40,
    58306 => -40,
    58307 => -40,
    58308 => -40,
    58309 => -40,
    58310 => -40,
    58311 => -40,
    58312 => -40,
    58313 => -40,
    58314 => -40,
    58315 => -40,
    58316 => -40,
    58317 => -40,
    58318 => -40,
    58319 => -40,
    58320 => -40,
    58321 => -40,
    58322 => -40,
    58323 => -40,
    58324 => -40,
    58325 => -40,
    58326 => -40,
    58327 => -40,
    58328 => -40,
    58329 => -40,
    58330 => -40,
    58331 => -40,
    58332 => -40,
    58333 => -40,
    58334 => -40,
    58335 => -40,
    58336 => -40,
    58337 => -40,
    58338 => -40,
    58339 => -40,
    58340 => -40,
    58341 => -40,
    58342 => -40,
    58343 => -40,
    58344 => -40,
    58345 => -40,
    58346 => -40,
    58347 => -40,
    58348 => -40,
    58349 => -40,
    58350 => -40,
    58351 => -40,
    58352 => -40,
    58353 => -40,
    58354 => -40,
    58355 => -40,
    58356 => -40,
    58357 => -40,
    58358 => -40,
    58359 => -40,
    58360 => -40,
    58361 => -40,
    58362 => -40,
    58363 => -40,
    58364 => -40,
    58365 => -40,
    58366 => -40,
    58367 => -40,
    58368 => -40,
    58369 => -40,
    58370 => -40,
    58371 => -40,
    58372 => -40,
    58373 => -40,
    58374 => -40,
    58375 => -40,
    58376 => -40,
    58377 => -40,
    58378 => -40,
    58379 => -40,
    58380 => -40,
    58381 => -40,
    58382 => -40,
    58383 => -40,
    58384 => -40,
    58385 => -40,
    58386 => -40,
    58387 => -40,
    58388 => -40,
    58389 => -40,
    58390 => -40,
    58391 => -40,
    58392 => -40,
    58393 => -40,
    58394 => -40,
    58395 => -40,
    58396 => -40,
    58397 => -40,
    58398 => -40,
    58399 => -40,
    58400 => -40,
    58401 => -40,
    58402 => -40,
    58403 => -40,
    58404 => -40,
    58405 => -40,
    58406 => -40,
    58407 => -40,
    58408 => -40,
    58409 => -40,
    58410 => -40,
    58411 => -40,
    58412 => -40,
    58413 => -40,
    58414 => -40,
    58415 => -40,
    58416 => -40,
    58417 => -40,
    58418 => -40,
    58419 => -40,
    58420 => -40,
    58421 => -40,
    58422 => -40,
    58423 => -40,
    58424 => -40,
    58425 => -40,
    58426 => -40,
    58427 => -40,
    58428 => -40,
    58429 => -40,
    58430 => -40,
    58431 => -40,
    58432 => -40,
    58433 => -40,
    58434 => -40,
    58435 => -40,
    58436 => -40,
    58437 => -40,
    58438 => -40,
    58439 => -40,
    58440 => -40,
    58441 => -40,
    58442 => -40,
    58443 => -40,
    58444 => -40,
    58445 => -40,
    58446 => -40,
    58447 => -40,
    58448 => -40,
    58449 => -40,
    58450 => -40,
    58451 => -40,
    58452 => -40,
    58453 => -40,
    58454 => -40,
    58455 => -40,
    58456 => -40,
    58457 => -40,
    58458 => -40,
    58459 => -40,
    58460 => -40,
    58461 => -40,
    58462 => -40,
    58463 => -40,
    58464 => -40,
    58465 => -40,
    58466 => -40,
    58467 => -40,
    58468 => -39,
    58469 => -39,
    58470 => -39,
    58471 => -39,
    58472 => -39,
    58473 => -39,
    58474 => -39,
    58475 => -39,
    58476 => -39,
    58477 => -39,
    58478 => -39,
    58479 => -39,
    58480 => -39,
    58481 => -39,
    58482 => -39,
    58483 => -39,
    58484 => -39,
    58485 => -39,
    58486 => -39,
    58487 => -39,
    58488 => -39,
    58489 => -39,
    58490 => -39,
    58491 => -39,
    58492 => -39,
    58493 => -39,
    58494 => -39,
    58495 => -39,
    58496 => -39,
    58497 => -39,
    58498 => -39,
    58499 => -39,
    58500 => -39,
    58501 => -39,
    58502 => -39,
    58503 => -39,
    58504 => -39,
    58505 => -39,
    58506 => -39,
    58507 => -39,
    58508 => -39,
    58509 => -39,
    58510 => -39,
    58511 => -39,
    58512 => -39,
    58513 => -39,
    58514 => -39,
    58515 => -39,
    58516 => -39,
    58517 => -39,
    58518 => -39,
    58519 => -39,
    58520 => -39,
    58521 => -39,
    58522 => -39,
    58523 => -39,
    58524 => -39,
    58525 => -39,
    58526 => -39,
    58527 => -39,
    58528 => -39,
    58529 => -39,
    58530 => -39,
    58531 => -39,
    58532 => -39,
    58533 => -39,
    58534 => -39,
    58535 => -39,
    58536 => -39,
    58537 => -39,
    58538 => -39,
    58539 => -39,
    58540 => -39,
    58541 => -39,
    58542 => -39,
    58543 => -39,
    58544 => -39,
    58545 => -39,
    58546 => -39,
    58547 => -39,
    58548 => -39,
    58549 => -39,
    58550 => -39,
    58551 => -39,
    58552 => -39,
    58553 => -39,
    58554 => -39,
    58555 => -39,
    58556 => -39,
    58557 => -39,
    58558 => -39,
    58559 => -39,
    58560 => -39,
    58561 => -39,
    58562 => -39,
    58563 => -39,
    58564 => -39,
    58565 => -39,
    58566 => -39,
    58567 => -39,
    58568 => -39,
    58569 => -39,
    58570 => -39,
    58571 => -39,
    58572 => -39,
    58573 => -39,
    58574 => -39,
    58575 => -39,
    58576 => -39,
    58577 => -39,
    58578 => -39,
    58579 => -39,
    58580 => -39,
    58581 => -39,
    58582 => -39,
    58583 => -39,
    58584 => -39,
    58585 => -39,
    58586 => -39,
    58587 => -39,
    58588 => -39,
    58589 => -39,
    58590 => -39,
    58591 => -39,
    58592 => -39,
    58593 => -39,
    58594 => -39,
    58595 => -39,
    58596 => -39,
    58597 => -39,
    58598 => -39,
    58599 => -39,
    58600 => -39,
    58601 => -39,
    58602 => -39,
    58603 => -39,
    58604 => -39,
    58605 => -39,
    58606 => -39,
    58607 => -39,
    58608 => -39,
    58609 => -39,
    58610 => -39,
    58611 => -39,
    58612 => -39,
    58613 => -39,
    58614 => -39,
    58615 => -39,
    58616 => -39,
    58617 => -39,
    58618 => -39,
    58619 => -39,
    58620 => -39,
    58621 => -39,
    58622 => -39,
    58623 => -39,
    58624 => -39,
    58625 => -39,
    58626 => -39,
    58627 => -39,
    58628 => -39,
    58629 => -39,
    58630 => -39,
    58631 => -39,
    58632 => -39,
    58633 => -39,
    58634 => -39,
    58635 => -39,
    58636 => -39,
    58637 => -39,
    58638 => -39,
    58639 => -39,
    58640 => -39,
    58641 => -39,
    58642 => -39,
    58643 => -39,
    58644 => -39,
    58645 => -39,
    58646 => -39,
    58647 => -39,
    58648 => -39,
    58649 => -39,
    58650 => -39,
    58651 => -39,
    58652 => -39,
    58653 => -39,
    58654 => -39,
    58655 => -39,
    58656 => -39,
    58657 => -39,
    58658 => -39,
    58659 => -39,
    58660 => -39,
    58661 => -39,
    58662 => -39,
    58663 => -39,
    58664 => -39,
    58665 => -39,
    58666 => -39,
    58667 => -39,
    58668 => -39,
    58669 => -39,
    58670 => -39,
    58671 => -39,
    58672 => -39,
    58673 => -39,
    58674 => -39,
    58675 => -39,
    58676 => -39,
    58677 => -39,
    58678 => -39,
    58679 => -38,
    58680 => -38,
    58681 => -38,
    58682 => -38,
    58683 => -38,
    58684 => -38,
    58685 => -38,
    58686 => -38,
    58687 => -38,
    58688 => -38,
    58689 => -38,
    58690 => -38,
    58691 => -38,
    58692 => -38,
    58693 => -38,
    58694 => -38,
    58695 => -38,
    58696 => -38,
    58697 => -38,
    58698 => -38,
    58699 => -38,
    58700 => -38,
    58701 => -38,
    58702 => -38,
    58703 => -38,
    58704 => -38,
    58705 => -38,
    58706 => -38,
    58707 => -38,
    58708 => -38,
    58709 => -38,
    58710 => -38,
    58711 => -38,
    58712 => -38,
    58713 => -38,
    58714 => -38,
    58715 => -38,
    58716 => -38,
    58717 => -38,
    58718 => -38,
    58719 => -38,
    58720 => -38,
    58721 => -38,
    58722 => -38,
    58723 => -38,
    58724 => -38,
    58725 => -38,
    58726 => -38,
    58727 => -38,
    58728 => -38,
    58729 => -38,
    58730 => -38,
    58731 => -38,
    58732 => -38,
    58733 => -38,
    58734 => -38,
    58735 => -38,
    58736 => -38,
    58737 => -38,
    58738 => -38,
    58739 => -38,
    58740 => -38,
    58741 => -38,
    58742 => -38,
    58743 => -38,
    58744 => -38,
    58745 => -38,
    58746 => -38,
    58747 => -38,
    58748 => -38,
    58749 => -38,
    58750 => -38,
    58751 => -38,
    58752 => -38,
    58753 => -38,
    58754 => -38,
    58755 => -38,
    58756 => -38,
    58757 => -38,
    58758 => -38,
    58759 => -38,
    58760 => -38,
    58761 => -38,
    58762 => -38,
    58763 => -38,
    58764 => -38,
    58765 => -38,
    58766 => -38,
    58767 => -38,
    58768 => -38,
    58769 => -38,
    58770 => -38,
    58771 => -38,
    58772 => -38,
    58773 => -38,
    58774 => -38,
    58775 => -38,
    58776 => -38,
    58777 => -38,
    58778 => -38,
    58779 => -38,
    58780 => -38,
    58781 => -38,
    58782 => -38,
    58783 => -38,
    58784 => -38,
    58785 => -38,
    58786 => -38,
    58787 => -38,
    58788 => -38,
    58789 => -38,
    58790 => -38,
    58791 => -38,
    58792 => -38,
    58793 => -38,
    58794 => -38,
    58795 => -38,
    58796 => -38,
    58797 => -38,
    58798 => -38,
    58799 => -38,
    58800 => -38,
    58801 => -38,
    58802 => -38,
    58803 => -38,
    58804 => -38,
    58805 => -38,
    58806 => -38,
    58807 => -38,
    58808 => -38,
    58809 => -38,
    58810 => -38,
    58811 => -38,
    58812 => -38,
    58813 => -38,
    58814 => -38,
    58815 => -38,
    58816 => -38,
    58817 => -38,
    58818 => -38,
    58819 => -38,
    58820 => -38,
    58821 => -38,
    58822 => -38,
    58823 => -38,
    58824 => -38,
    58825 => -38,
    58826 => -38,
    58827 => -38,
    58828 => -38,
    58829 => -38,
    58830 => -38,
    58831 => -38,
    58832 => -38,
    58833 => -38,
    58834 => -38,
    58835 => -38,
    58836 => -38,
    58837 => -38,
    58838 => -38,
    58839 => -38,
    58840 => -38,
    58841 => -38,
    58842 => -38,
    58843 => -38,
    58844 => -38,
    58845 => -38,
    58846 => -38,
    58847 => -38,
    58848 => -38,
    58849 => -38,
    58850 => -38,
    58851 => -38,
    58852 => -38,
    58853 => -38,
    58854 => -38,
    58855 => -38,
    58856 => -38,
    58857 => -38,
    58858 => -38,
    58859 => -38,
    58860 => -38,
    58861 => -38,
    58862 => -38,
    58863 => -38,
    58864 => -38,
    58865 => -38,
    58866 => -38,
    58867 => -38,
    58868 => -38,
    58869 => -38,
    58870 => -38,
    58871 => -38,
    58872 => -38,
    58873 => -38,
    58874 => -38,
    58875 => -38,
    58876 => -38,
    58877 => -38,
    58878 => -38,
    58879 => -38,
    58880 => -38,
    58881 => -38,
    58882 => -38,
    58883 => -38,
    58884 => -38,
    58885 => -38,
    58886 => -37,
    58887 => -37,
    58888 => -37,
    58889 => -37,
    58890 => -37,
    58891 => -37,
    58892 => -37,
    58893 => -37,
    58894 => -37,
    58895 => -37,
    58896 => -37,
    58897 => -37,
    58898 => -37,
    58899 => -37,
    58900 => -37,
    58901 => -37,
    58902 => -37,
    58903 => -37,
    58904 => -37,
    58905 => -37,
    58906 => -37,
    58907 => -37,
    58908 => -37,
    58909 => -37,
    58910 => -37,
    58911 => -37,
    58912 => -37,
    58913 => -37,
    58914 => -37,
    58915 => -37,
    58916 => -37,
    58917 => -37,
    58918 => -37,
    58919 => -37,
    58920 => -37,
    58921 => -37,
    58922 => -37,
    58923 => -37,
    58924 => -37,
    58925 => -37,
    58926 => -37,
    58927 => -37,
    58928 => -37,
    58929 => -37,
    58930 => -37,
    58931 => -37,
    58932 => -37,
    58933 => -37,
    58934 => -37,
    58935 => -37,
    58936 => -37,
    58937 => -37,
    58938 => -37,
    58939 => -37,
    58940 => -37,
    58941 => -37,
    58942 => -37,
    58943 => -37,
    58944 => -37,
    58945 => -37,
    58946 => -37,
    58947 => -37,
    58948 => -37,
    58949 => -37,
    58950 => -37,
    58951 => -37,
    58952 => -37,
    58953 => -37,
    58954 => -37,
    58955 => -37,
    58956 => -37,
    58957 => -37,
    58958 => -37,
    58959 => -37,
    58960 => -37,
    58961 => -37,
    58962 => -37,
    58963 => -37,
    58964 => -37,
    58965 => -37,
    58966 => -37,
    58967 => -37,
    58968 => -37,
    58969 => -37,
    58970 => -37,
    58971 => -37,
    58972 => -37,
    58973 => -37,
    58974 => -37,
    58975 => -37,
    58976 => -37,
    58977 => -37,
    58978 => -37,
    58979 => -37,
    58980 => -37,
    58981 => -37,
    58982 => -37,
    58983 => -37,
    58984 => -37,
    58985 => -37,
    58986 => -37,
    58987 => -37,
    58988 => -37,
    58989 => -37,
    58990 => -37,
    58991 => -37,
    58992 => -37,
    58993 => -37,
    58994 => -37,
    58995 => -37,
    58996 => -37,
    58997 => -37,
    58998 => -37,
    58999 => -37,
    59000 => -37,
    59001 => -37,
    59002 => -37,
    59003 => -37,
    59004 => -37,
    59005 => -37,
    59006 => -37,
    59007 => -37,
    59008 => -37,
    59009 => -37,
    59010 => -37,
    59011 => -37,
    59012 => -37,
    59013 => -37,
    59014 => -37,
    59015 => -37,
    59016 => -37,
    59017 => -37,
    59018 => -37,
    59019 => -37,
    59020 => -37,
    59021 => -37,
    59022 => -37,
    59023 => -37,
    59024 => -37,
    59025 => -37,
    59026 => -37,
    59027 => -37,
    59028 => -37,
    59029 => -37,
    59030 => -37,
    59031 => -37,
    59032 => -37,
    59033 => -37,
    59034 => -37,
    59035 => -37,
    59036 => -37,
    59037 => -37,
    59038 => -37,
    59039 => -37,
    59040 => -37,
    59041 => -37,
    59042 => -37,
    59043 => -37,
    59044 => -37,
    59045 => -37,
    59046 => -37,
    59047 => -37,
    59048 => -37,
    59049 => -37,
    59050 => -37,
    59051 => -37,
    59052 => -37,
    59053 => -37,
    59054 => -37,
    59055 => -37,
    59056 => -37,
    59057 => -37,
    59058 => -37,
    59059 => -37,
    59060 => -37,
    59061 => -37,
    59062 => -37,
    59063 => -37,
    59064 => -37,
    59065 => -37,
    59066 => -37,
    59067 => -37,
    59068 => -37,
    59069 => -37,
    59070 => -37,
    59071 => -37,
    59072 => -37,
    59073 => -37,
    59074 => -37,
    59075 => -37,
    59076 => -37,
    59077 => -37,
    59078 => -37,
    59079 => -37,
    59080 => -37,
    59081 => -37,
    59082 => -37,
    59083 => -37,
    59084 => -37,
    59085 => -37,
    59086 => -37,
    59087 => -37,
    59088 => -37,
    59089 => -37,
    59090 => -37,
    59091 => -36,
    59092 => -36,
    59093 => -36,
    59094 => -36,
    59095 => -36,
    59096 => -36,
    59097 => -36,
    59098 => -36,
    59099 => -36,
    59100 => -36,
    59101 => -36,
    59102 => -36,
    59103 => -36,
    59104 => -36,
    59105 => -36,
    59106 => -36,
    59107 => -36,
    59108 => -36,
    59109 => -36,
    59110 => -36,
    59111 => -36,
    59112 => -36,
    59113 => -36,
    59114 => -36,
    59115 => -36,
    59116 => -36,
    59117 => -36,
    59118 => -36,
    59119 => -36,
    59120 => -36,
    59121 => -36,
    59122 => -36,
    59123 => -36,
    59124 => -36,
    59125 => -36,
    59126 => -36,
    59127 => -36,
    59128 => -36,
    59129 => -36,
    59130 => -36,
    59131 => -36,
    59132 => -36,
    59133 => -36,
    59134 => -36,
    59135 => -36,
    59136 => -36,
    59137 => -36,
    59138 => -36,
    59139 => -36,
    59140 => -36,
    59141 => -36,
    59142 => -36,
    59143 => -36,
    59144 => -36,
    59145 => -36,
    59146 => -36,
    59147 => -36,
    59148 => -36,
    59149 => -36,
    59150 => -36,
    59151 => -36,
    59152 => -36,
    59153 => -36,
    59154 => -36,
    59155 => -36,
    59156 => -36,
    59157 => -36,
    59158 => -36,
    59159 => -36,
    59160 => -36,
    59161 => -36,
    59162 => -36,
    59163 => -36,
    59164 => -36,
    59165 => -36,
    59166 => -36,
    59167 => -36,
    59168 => -36,
    59169 => -36,
    59170 => -36,
    59171 => -36,
    59172 => -36,
    59173 => -36,
    59174 => -36,
    59175 => -36,
    59176 => -36,
    59177 => -36,
    59178 => -36,
    59179 => -36,
    59180 => -36,
    59181 => -36,
    59182 => -36,
    59183 => -36,
    59184 => -36,
    59185 => -36,
    59186 => -36,
    59187 => -36,
    59188 => -36,
    59189 => -36,
    59190 => -36,
    59191 => -36,
    59192 => -36,
    59193 => -36,
    59194 => -36,
    59195 => -36,
    59196 => -36,
    59197 => -36,
    59198 => -36,
    59199 => -36,
    59200 => -36,
    59201 => -36,
    59202 => -36,
    59203 => -36,
    59204 => -36,
    59205 => -36,
    59206 => -36,
    59207 => -36,
    59208 => -36,
    59209 => -36,
    59210 => -36,
    59211 => -36,
    59212 => -36,
    59213 => -36,
    59214 => -36,
    59215 => -36,
    59216 => -36,
    59217 => -36,
    59218 => -36,
    59219 => -36,
    59220 => -36,
    59221 => -36,
    59222 => -36,
    59223 => -36,
    59224 => -36,
    59225 => -36,
    59226 => -36,
    59227 => -36,
    59228 => -36,
    59229 => -36,
    59230 => -36,
    59231 => -36,
    59232 => -36,
    59233 => -36,
    59234 => -36,
    59235 => -36,
    59236 => -36,
    59237 => -36,
    59238 => -36,
    59239 => -36,
    59240 => -36,
    59241 => -36,
    59242 => -36,
    59243 => -36,
    59244 => -36,
    59245 => -36,
    59246 => -36,
    59247 => -36,
    59248 => -36,
    59249 => -36,
    59250 => -36,
    59251 => -36,
    59252 => -36,
    59253 => -36,
    59254 => -36,
    59255 => -36,
    59256 => -36,
    59257 => -36,
    59258 => -36,
    59259 => -36,
    59260 => -36,
    59261 => -36,
    59262 => -36,
    59263 => -36,
    59264 => -36,
    59265 => -36,
    59266 => -36,
    59267 => -36,
    59268 => -36,
    59269 => -36,
    59270 => -36,
    59271 => -36,
    59272 => -36,
    59273 => -36,
    59274 => -36,
    59275 => -36,
    59276 => -36,
    59277 => -36,
    59278 => -36,
    59279 => -36,
    59280 => -36,
    59281 => -36,
    59282 => -36,
    59283 => -36,
    59284 => -36,
    59285 => -36,
    59286 => -36,
    59287 => -36,
    59288 => -36,
    59289 => -36,
    59290 => -36,
    59291 => -36,
    59292 => -36,
    59293 => -35,
    59294 => -35,
    59295 => -35,
    59296 => -35,
    59297 => -35,
    59298 => -35,
    59299 => -35,
    59300 => -35,
    59301 => -35,
    59302 => -35,
    59303 => -35,
    59304 => -35,
    59305 => -35,
    59306 => -35,
    59307 => -35,
    59308 => -35,
    59309 => -35,
    59310 => -35,
    59311 => -35,
    59312 => -35,
    59313 => -35,
    59314 => -35,
    59315 => -35,
    59316 => -35,
    59317 => -35,
    59318 => -35,
    59319 => -35,
    59320 => -35,
    59321 => -35,
    59322 => -35,
    59323 => -35,
    59324 => -35,
    59325 => -35,
    59326 => -35,
    59327 => -35,
    59328 => -35,
    59329 => -35,
    59330 => -35,
    59331 => -35,
    59332 => -35,
    59333 => -35,
    59334 => -35,
    59335 => -35,
    59336 => -35,
    59337 => -35,
    59338 => -35,
    59339 => -35,
    59340 => -35,
    59341 => -35,
    59342 => -35,
    59343 => -35,
    59344 => -35,
    59345 => -35,
    59346 => -35,
    59347 => -35,
    59348 => -35,
    59349 => -35,
    59350 => -35,
    59351 => -35,
    59352 => -35,
    59353 => -35,
    59354 => -35,
    59355 => -35,
    59356 => -35,
    59357 => -35,
    59358 => -35,
    59359 => -35,
    59360 => -35,
    59361 => -35,
    59362 => -35,
    59363 => -35,
    59364 => -35,
    59365 => -35,
    59366 => -35,
    59367 => -35,
    59368 => -35,
    59369 => -35,
    59370 => -35,
    59371 => -35,
    59372 => -35,
    59373 => -35,
    59374 => -35,
    59375 => -35,
    59376 => -35,
    59377 => -35,
    59378 => -35,
    59379 => -35,
    59380 => -35,
    59381 => -35,
    59382 => -35,
    59383 => -35,
    59384 => -35,
    59385 => -35,
    59386 => -35,
    59387 => -35,
    59388 => -35,
    59389 => -35,
    59390 => -35,
    59391 => -35,
    59392 => -35,
    59393 => -35,
    59394 => -35,
    59395 => -35,
    59396 => -35,
    59397 => -35,
    59398 => -35,
    59399 => -35,
    59400 => -35,
    59401 => -35,
    59402 => -35,
    59403 => -35,
    59404 => -35,
    59405 => -35,
    59406 => -35,
    59407 => -35,
    59408 => -35,
    59409 => -35,
    59410 => -35,
    59411 => -35,
    59412 => -35,
    59413 => -35,
    59414 => -35,
    59415 => -35,
    59416 => -35,
    59417 => -35,
    59418 => -35,
    59419 => -35,
    59420 => -35,
    59421 => -35,
    59422 => -35,
    59423 => -35,
    59424 => -35,
    59425 => -35,
    59426 => -35,
    59427 => -35,
    59428 => -35,
    59429 => -35,
    59430 => -35,
    59431 => -35,
    59432 => -35,
    59433 => -35,
    59434 => -35,
    59435 => -35,
    59436 => -35,
    59437 => -35,
    59438 => -35,
    59439 => -35,
    59440 => -35,
    59441 => -35,
    59442 => -35,
    59443 => -35,
    59444 => -35,
    59445 => -35,
    59446 => -35,
    59447 => -35,
    59448 => -35,
    59449 => -35,
    59450 => -35,
    59451 => -35,
    59452 => -35,
    59453 => -35,
    59454 => -35,
    59455 => -35,
    59456 => -35,
    59457 => -35,
    59458 => -35,
    59459 => -35,
    59460 => -35,
    59461 => -35,
    59462 => -35,
    59463 => -35,
    59464 => -35,
    59465 => -35,
    59466 => -35,
    59467 => -35,
    59468 => -35,
    59469 => -35,
    59470 => -35,
    59471 => -35,
    59472 => -35,
    59473 => -35,
    59474 => -35,
    59475 => -35,
    59476 => -35,
    59477 => -35,
    59478 => -35,
    59479 => -35,
    59480 => -35,
    59481 => -35,
    59482 => -35,
    59483 => -35,
    59484 => -35,
    59485 => -35,
    59486 => -35,
    59487 => -35,
    59488 => -35,
    59489 => -35,
    59490 => -35,
    59491 => -35,
    59492 => -34,
    59493 => -34,
    59494 => -34,
    59495 => -34,
    59496 => -34,
    59497 => -34,
    59498 => -34,
    59499 => -34,
    59500 => -34,
    59501 => -34,
    59502 => -34,
    59503 => -34,
    59504 => -34,
    59505 => -34,
    59506 => -34,
    59507 => -34,
    59508 => -34,
    59509 => -34,
    59510 => -34,
    59511 => -34,
    59512 => -34,
    59513 => -34,
    59514 => -34,
    59515 => -34,
    59516 => -34,
    59517 => -34,
    59518 => -34,
    59519 => -34,
    59520 => -34,
    59521 => -34,
    59522 => -34,
    59523 => -34,
    59524 => -34,
    59525 => -34,
    59526 => -34,
    59527 => -34,
    59528 => -34,
    59529 => -34,
    59530 => -34,
    59531 => -34,
    59532 => -34,
    59533 => -34,
    59534 => -34,
    59535 => -34,
    59536 => -34,
    59537 => -34,
    59538 => -34,
    59539 => -34,
    59540 => -34,
    59541 => -34,
    59542 => -34,
    59543 => -34,
    59544 => -34,
    59545 => -34,
    59546 => -34,
    59547 => -34,
    59548 => -34,
    59549 => -34,
    59550 => -34,
    59551 => -34,
    59552 => -34,
    59553 => -34,
    59554 => -34,
    59555 => -34,
    59556 => -34,
    59557 => -34,
    59558 => -34,
    59559 => -34,
    59560 => -34,
    59561 => -34,
    59562 => -34,
    59563 => -34,
    59564 => -34,
    59565 => -34,
    59566 => -34,
    59567 => -34,
    59568 => -34,
    59569 => -34,
    59570 => -34,
    59571 => -34,
    59572 => -34,
    59573 => -34,
    59574 => -34,
    59575 => -34,
    59576 => -34,
    59577 => -34,
    59578 => -34,
    59579 => -34,
    59580 => -34,
    59581 => -34,
    59582 => -34,
    59583 => -34,
    59584 => -34,
    59585 => -34,
    59586 => -34,
    59587 => -34,
    59588 => -34,
    59589 => -34,
    59590 => -34,
    59591 => -34,
    59592 => -34,
    59593 => -34,
    59594 => -34,
    59595 => -34,
    59596 => -34,
    59597 => -34,
    59598 => -34,
    59599 => -34,
    59600 => -34,
    59601 => -34,
    59602 => -34,
    59603 => -34,
    59604 => -34,
    59605 => -34,
    59606 => -34,
    59607 => -34,
    59608 => -34,
    59609 => -34,
    59610 => -34,
    59611 => -34,
    59612 => -34,
    59613 => -34,
    59614 => -34,
    59615 => -34,
    59616 => -34,
    59617 => -34,
    59618 => -34,
    59619 => -34,
    59620 => -34,
    59621 => -34,
    59622 => -34,
    59623 => -34,
    59624 => -34,
    59625 => -34,
    59626 => -34,
    59627 => -34,
    59628 => -34,
    59629 => -34,
    59630 => -34,
    59631 => -34,
    59632 => -34,
    59633 => -34,
    59634 => -34,
    59635 => -34,
    59636 => -34,
    59637 => -34,
    59638 => -34,
    59639 => -34,
    59640 => -34,
    59641 => -34,
    59642 => -34,
    59643 => -34,
    59644 => -34,
    59645 => -34,
    59646 => -34,
    59647 => -34,
    59648 => -34,
    59649 => -34,
    59650 => -34,
    59651 => -34,
    59652 => -34,
    59653 => -34,
    59654 => -34,
    59655 => -34,
    59656 => -34,
    59657 => -34,
    59658 => -34,
    59659 => -34,
    59660 => -34,
    59661 => -34,
    59662 => -34,
    59663 => -34,
    59664 => -34,
    59665 => -34,
    59666 => -34,
    59667 => -34,
    59668 => -34,
    59669 => -34,
    59670 => -34,
    59671 => -34,
    59672 => -34,
    59673 => -34,
    59674 => -34,
    59675 => -34,
    59676 => -34,
    59677 => -34,
    59678 => -34,
    59679 => -34,
    59680 => -34,
    59681 => -34,
    59682 => -34,
    59683 => -34,
    59684 => -34,
    59685 => -34,
    59686 => -34,
    59687 => -34,
    59688 => -34,
    59689 => -33,
    59690 => -33,
    59691 => -33,
    59692 => -33,
    59693 => -33,
    59694 => -33,
    59695 => -33,
    59696 => -33,
    59697 => -33,
    59698 => -33,
    59699 => -33,
    59700 => -33,
    59701 => -33,
    59702 => -33,
    59703 => -33,
    59704 => -33,
    59705 => -33,
    59706 => -33,
    59707 => -33,
    59708 => -33,
    59709 => -33,
    59710 => -33,
    59711 => -33,
    59712 => -33,
    59713 => -33,
    59714 => -33,
    59715 => -33,
    59716 => -33,
    59717 => -33,
    59718 => -33,
    59719 => -33,
    59720 => -33,
    59721 => -33,
    59722 => -33,
    59723 => -33,
    59724 => -33,
    59725 => -33,
    59726 => -33,
    59727 => -33,
    59728 => -33,
    59729 => -33,
    59730 => -33,
    59731 => -33,
    59732 => -33,
    59733 => -33,
    59734 => -33,
    59735 => -33,
    59736 => -33,
    59737 => -33,
    59738 => -33,
    59739 => -33,
    59740 => -33,
    59741 => -33,
    59742 => -33,
    59743 => -33,
    59744 => -33,
    59745 => -33,
    59746 => -33,
    59747 => -33,
    59748 => -33,
    59749 => -33,
    59750 => -33,
    59751 => -33,
    59752 => -33,
    59753 => -33,
    59754 => -33,
    59755 => -33,
    59756 => -33,
    59757 => -33,
    59758 => -33,
    59759 => -33,
    59760 => -33,
    59761 => -33,
    59762 => -33,
    59763 => -33,
    59764 => -33,
    59765 => -33,
    59766 => -33,
    59767 => -33,
    59768 => -33,
    59769 => -33,
    59770 => -33,
    59771 => -33,
    59772 => -33,
    59773 => -33,
    59774 => -33,
    59775 => -33,
    59776 => -33,
    59777 => -33,
    59778 => -33,
    59779 => -33,
    59780 => -33,
    59781 => -33,
    59782 => -33,
    59783 => -33,
    59784 => -33,
    59785 => -33,
    59786 => -33,
    59787 => -33,
    59788 => -33,
    59789 => -33,
    59790 => -33,
    59791 => -33,
    59792 => -33,
    59793 => -33,
    59794 => -33,
    59795 => -33,
    59796 => -33,
    59797 => -33,
    59798 => -33,
    59799 => -33,
    59800 => -33,
    59801 => -33,
    59802 => -33,
    59803 => -33,
    59804 => -33,
    59805 => -33,
    59806 => -33,
    59807 => -33,
    59808 => -33,
    59809 => -33,
    59810 => -33,
    59811 => -33,
    59812 => -33,
    59813 => -33,
    59814 => -33,
    59815 => -33,
    59816 => -33,
    59817 => -33,
    59818 => -33,
    59819 => -33,
    59820 => -33,
    59821 => -33,
    59822 => -33,
    59823 => -33,
    59824 => -33,
    59825 => -33,
    59826 => -33,
    59827 => -33,
    59828 => -33,
    59829 => -33,
    59830 => -33,
    59831 => -33,
    59832 => -33,
    59833 => -33,
    59834 => -33,
    59835 => -33,
    59836 => -33,
    59837 => -33,
    59838 => -33,
    59839 => -33,
    59840 => -33,
    59841 => -33,
    59842 => -33,
    59843 => -33,
    59844 => -33,
    59845 => -33,
    59846 => -33,
    59847 => -33,
    59848 => -33,
    59849 => -33,
    59850 => -33,
    59851 => -33,
    59852 => -33,
    59853 => -33,
    59854 => -33,
    59855 => -33,
    59856 => -33,
    59857 => -33,
    59858 => -33,
    59859 => -33,
    59860 => -33,
    59861 => -33,
    59862 => -33,
    59863 => -33,
    59864 => -33,
    59865 => -33,
    59866 => -33,
    59867 => -33,
    59868 => -33,
    59869 => -33,
    59870 => -33,
    59871 => -33,
    59872 => -33,
    59873 => -33,
    59874 => -33,
    59875 => -33,
    59876 => -33,
    59877 => -33,
    59878 => -33,
    59879 => -33,
    59880 => -33,
    59881 => -33,
    59882 => -33,
    59883 => -32,
    59884 => -32,
    59885 => -32,
    59886 => -32,
    59887 => -32,
    59888 => -32,
    59889 => -32,
    59890 => -32,
    59891 => -32,
    59892 => -32,
    59893 => -32,
    59894 => -32,
    59895 => -32,
    59896 => -32,
    59897 => -32,
    59898 => -32,
    59899 => -32,
    59900 => -32,
    59901 => -32,
    59902 => -32,
    59903 => -32,
    59904 => -32,
    59905 => -32,
    59906 => -32,
    59907 => -32,
    59908 => -32,
    59909 => -32,
    59910 => -32,
    59911 => -32,
    59912 => -32,
    59913 => -32,
    59914 => -32,
    59915 => -32,
    59916 => -32,
    59917 => -32,
    59918 => -32,
    59919 => -32,
    59920 => -32,
    59921 => -32,
    59922 => -32,
    59923 => -32,
    59924 => -32,
    59925 => -32,
    59926 => -32,
    59927 => -32,
    59928 => -32,
    59929 => -32,
    59930 => -32,
    59931 => -32,
    59932 => -32,
    59933 => -32,
    59934 => -32,
    59935 => -32,
    59936 => -32,
    59937 => -32,
    59938 => -32,
    59939 => -32,
    59940 => -32,
    59941 => -32,
    59942 => -32,
    59943 => -32,
    59944 => -32,
    59945 => -32,
    59946 => -32,
    59947 => -32,
    59948 => -32,
    59949 => -32,
    59950 => -32,
    59951 => -32,
    59952 => -32,
    59953 => -32,
    59954 => -32,
    59955 => -32,
    59956 => -32,
    59957 => -32,
    59958 => -32,
    59959 => -32,
    59960 => -32,
    59961 => -32,
    59962 => -32,
    59963 => -32,
    59964 => -32,
    59965 => -32,
    59966 => -32,
    59967 => -32,
    59968 => -32,
    59969 => -32,
    59970 => -32,
    59971 => -32,
    59972 => -32,
    59973 => -32,
    59974 => -32,
    59975 => -32,
    59976 => -32,
    59977 => -32,
    59978 => -32,
    59979 => -32,
    59980 => -32,
    59981 => -32,
    59982 => -32,
    59983 => -32,
    59984 => -32,
    59985 => -32,
    59986 => -32,
    59987 => -32,
    59988 => -32,
    59989 => -32,
    59990 => -32,
    59991 => -32,
    59992 => -32,
    59993 => -32,
    59994 => -32,
    59995 => -32,
    59996 => -32,
    59997 => -32,
    59998 => -32,
    59999 => -32,
    60000 => -32,
    60001 => -32,
    60002 => -32,
    60003 => -32,
    60004 => -32,
    60005 => -32,
    60006 => -32,
    60007 => -32,
    60008 => -32,
    60009 => -32,
    60010 => -32,
    60011 => -32,
    60012 => -32,
    60013 => -32,
    60014 => -32,
    60015 => -32,
    60016 => -32,
    60017 => -32,
    60018 => -32,
    60019 => -32,
    60020 => -32,
    60021 => -32,
    60022 => -32,
    60023 => -32,
    60024 => -32,
    60025 => -32,
    60026 => -32,
    60027 => -32,
    60028 => -32,
    60029 => -32,
    60030 => -32,
    60031 => -32,
    60032 => -32,
    60033 => -32,
    60034 => -32,
    60035 => -32,
    60036 => -32,
    60037 => -32,
    60038 => -32,
    60039 => -32,
    60040 => -32,
    60041 => -32,
    60042 => -32,
    60043 => -32,
    60044 => -32,
    60045 => -32,
    60046 => -32,
    60047 => -32,
    60048 => -32,
    60049 => -32,
    60050 => -32,
    60051 => -32,
    60052 => -32,
    60053 => -32,
    60054 => -32,
    60055 => -32,
    60056 => -32,
    60057 => -32,
    60058 => -32,
    60059 => -32,
    60060 => -32,
    60061 => -32,
    60062 => -32,
    60063 => -32,
    60064 => -32,
    60065 => -32,
    60066 => -32,
    60067 => -32,
    60068 => -32,
    60069 => -32,
    60070 => -32,
    60071 => -32,
    60072 => -32,
    60073 => -32,
    60074 => -32,
    60075 => -31,
    60076 => -31,
    60077 => -31,
    60078 => -31,
    60079 => -31,
    60080 => -31,
    60081 => -31,
    60082 => -31,
    60083 => -31,
    60084 => -31,
    60085 => -31,
    60086 => -31,
    60087 => -31,
    60088 => -31,
    60089 => -31,
    60090 => -31,
    60091 => -31,
    60092 => -31,
    60093 => -31,
    60094 => -31,
    60095 => -31,
    60096 => -31,
    60097 => -31,
    60098 => -31,
    60099 => -31,
    60100 => -31,
    60101 => -31,
    60102 => -31,
    60103 => -31,
    60104 => -31,
    60105 => -31,
    60106 => -31,
    60107 => -31,
    60108 => -31,
    60109 => -31,
    60110 => -31,
    60111 => -31,
    60112 => -31,
    60113 => -31,
    60114 => -31,
    60115 => -31,
    60116 => -31,
    60117 => -31,
    60118 => -31,
    60119 => -31,
    60120 => -31,
    60121 => -31,
    60122 => -31,
    60123 => -31,
    60124 => -31,
    60125 => -31,
    60126 => -31,
    60127 => -31,
    60128 => -31,
    60129 => -31,
    60130 => -31,
    60131 => -31,
    60132 => -31,
    60133 => -31,
    60134 => -31,
    60135 => -31,
    60136 => -31,
    60137 => -31,
    60138 => -31,
    60139 => -31,
    60140 => -31,
    60141 => -31,
    60142 => -31,
    60143 => -31,
    60144 => -31,
    60145 => -31,
    60146 => -31,
    60147 => -31,
    60148 => -31,
    60149 => -31,
    60150 => -31,
    60151 => -31,
    60152 => -31,
    60153 => -31,
    60154 => -31,
    60155 => -31,
    60156 => -31,
    60157 => -31,
    60158 => -31,
    60159 => -31,
    60160 => -31,
    60161 => -31,
    60162 => -31,
    60163 => -31,
    60164 => -31,
    60165 => -31,
    60166 => -31,
    60167 => -31,
    60168 => -31,
    60169 => -31,
    60170 => -31,
    60171 => -31,
    60172 => -31,
    60173 => -31,
    60174 => -31,
    60175 => -31,
    60176 => -31,
    60177 => -31,
    60178 => -31,
    60179 => -31,
    60180 => -31,
    60181 => -31,
    60182 => -31,
    60183 => -31,
    60184 => -31,
    60185 => -31,
    60186 => -31,
    60187 => -31,
    60188 => -31,
    60189 => -31,
    60190 => -31,
    60191 => -31,
    60192 => -31,
    60193 => -31,
    60194 => -31,
    60195 => -31,
    60196 => -31,
    60197 => -31,
    60198 => -31,
    60199 => -31,
    60200 => -31,
    60201 => -31,
    60202 => -31,
    60203 => -31,
    60204 => -31,
    60205 => -31,
    60206 => -31,
    60207 => -31,
    60208 => -31,
    60209 => -31,
    60210 => -31,
    60211 => -31,
    60212 => -31,
    60213 => -31,
    60214 => -31,
    60215 => -31,
    60216 => -31,
    60217 => -31,
    60218 => -31,
    60219 => -31,
    60220 => -31,
    60221 => -31,
    60222 => -31,
    60223 => -31,
    60224 => -31,
    60225 => -31,
    60226 => -31,
    60227 => -31,
    60228 => -31,
    60229 => -31,
    60230 => -31,
    60231 => -31,
    60232 => -31,
    60233 => -31,
    60234 => -31,
    60235 => -31,
    60236 => -31,
    60237 => -31,
    60238 => -31,
    60239 => -31,
    60240 => -31,
    60241 => -31,
    60242 => -31,
    60243 => -31,
    60244 => -31,
    60245 => -31,
    60246 => -31,
    60247 => -31,
    60248 => -31,
    60249 => -31,
    60250 => -31,
    60251 => -31,
    60252 => -31,
    60253 => -31,
    60254 => -31,
    60255 => -31,
    60256 => -31,
    60257 => -31,
    60258 => -31,
    60259 => -31,
    60260 => -31,
    60261 => -31,
    60262 => -31,
    60263 => -31,
    60264 => -31,
    60265 => -30,
    60266 => -30,
    60267 => -30,
    60268 => -30,
    60269 => -30,
    60270 => -30,
    60271 => -30,
    60272 => -30,
    60273 => -30,
    60274 => -30,
    60275 => -30,
    60276 => -30,
    60277 => -30,
    60278 => -30,
    60279 => -30,
    60280 => -30,
    60281 => -30,
    60282 => -30,
    60283 => -30,
    60284 => -30,
    60285 => -30,
    60286 => -30,
    60287 => -30,
    60288 => -30,
    60289 => -30,
    60290 => -30,
    60291 => -30,
    60292 => -30,
    60293 => -30,
    60294 => -30,
    60295 => -30,
    60296 => -30,
    60297 => -30,
    60298 => -30,
    60299 => -30,
    60300 => -30,
    60301 => -30,
    60302 => -30,
    60303 => -30,
    60304 => -30,
    60305 => -30,
    60306 => -30,
    60307 => -30,
    60308 => -30,
    60309 => -30,
    60310 => -30,
    60311 => -30,
    60312 => -30,
    60313 => -30,
    60314 => -30,
    60315 => -30,
    60316 => -30,
    60317 => -30,
    60318 => -30,
    60319 => -30,
    60320 => -30,
    60321 => -30,
    60322 => -30,
    60323 => -30,
    60324 => -30,
    60325 => -30,
    60326 => -30,
    60327 => -30,
    60328 => -30,
    60329 => -30,
    60330 => -30,
    60331 => -30,
    60332 => -30,
    60333 => -30,
    60334 => -30,
    60335 => -30,
    60336 => -30,
    60337 => -30,
    60338 => -30,
    60339 => -30,
    60340 => -30,
    60341 => -30,
    60342 => -30,
    60343 => -30,
    60344 => -30,
    60345 => -30,
    60346 => -30,
    60347 => -30,
    60348 => -30,
    60349 => -30,
    60350 => -30,
    60351 => -30,
    60352 => -30,
    60353 => -30,
    60354 => -30,
    60355 => -30,
    60356 => -30,
    60357 => -30,
    60358 => -30,
    60359 => -30,
    60360 => -30,
    60361 => -30,
    60362 => -30,
    60363 => -30,
    60364 => -30,
    60365 => -30,
    60366 => -30,
    60367 => -30,
    60368 => -30,
    60369 => -30,
    60370 => -30,
    60371 => -30,
    60372 => -30,
    60373 => -30,
    60374 => -30,
    60375 => -30,
    60376 => -30,
    60377 => -30,
    60378 => -30,
    60379 => -30,
    60380 => -30,
    60381 => -30,
    60382 => -30,
    60383 => -30,
    60384 => -30,
    60385 => -30,
    60386 => -30,
    60387 => -30,
    60388 => -30,
    60389 => -30,
    60390 => -30,
    60391 => -30,
    60392 => -30,
    60393 => -30,
    60394 => -30,
    60395 => -30,
    60396 => -30,
    60397 => -30,
    60398 => -30,
    60399 => -30,
    60400 => -30,
    60401 => -30,
    60402 => -30,
    60403 => -30,
    60404 => -30,
    60405 => -30,
    60406 => -30,
    60407 => -30,
    60408 => -30,
    60409 => -30,
    60410 => -30,
    60411 => -30,
    60412 => -30,
    60413 => -30,
    60414 => -30,
    60415 => -30,
    60416 => -30,
    60417 => -30,
    60418 => -30,
    60419 => -30,
    60420 => -30,
    60421 => -30,
    60422 => -30,
    60423 => -30,
    60424 => -30,
    60425 => -30,
    60426 => -30,
    60427 => -30,
    60428 => -30,
    60429 => -30,
    60430 => -30,
    60431 => -30,
    60432 => -30,
    60433 => -30,
    60434 => -30,
    60435 => -30,
    60436 => -30,
    60437 => -30,
    60438 => -30,
    60439 => -30,
    60440 => -30,
    60441 => -30,
    60442 => -30,
    60443 => -30,
    60444 => -30,
    60445 => -30,
    60446 => -30,
    60447 => -30,
    60448 => -30,
    60449 => -30,
    60450 => -30,
    60451 => -30,
    60452 => -30,
    60453 => -30,
    60454 => -29,
    60455 => -29,
    60456 => -29,
    60457 => -29,
    60458 => -29,
    60459 => -29,
    60460 => -29,
    60461 => -29,
    60462 => -29,
    60463 => -29,
    60464 => -29,
    60465 => -29,
    60466 => -29,
    60467 => -29,
    60468 => -29,
    60469 => -29,
    60470 => -29,
    60471 => -29,
    60472 => -29,
    60473 => -29,
    60474 => -29,
    60475 => -29,
    60476 => -29,
    60477 => -29,
    60478 => -29,
    60479 => -29,
    60480 => -29,
    60481 => -29,
    60482 => -29,
    60483 => -29,
    60484 => -29,
    60485 => -29,
    60486 => -29,
    60487 => -29,
    60488 => -29,
    60489 => -29,
    60490 => -29,
    60491 => -29,
    60492 => -29,
    60493 => -29,
    60494 => -29,
    60495 => -29,
    60496 => -29,
    60497 => -29,
    60498 => -29,
    60499 => -29,
    60500 => -29,
    60501 => -29,
    60502 => -29,
    60503 => -29,
    60504 => -29,
    60505 => -29,
    60506 => -29,
    60507 => -29,
    60508 => -29,
    60509 => -29,
    60510 => -29,
    60511 => -29,
    60512 => -29,
    60513 => -29,
    60514 => -29,
    60515 => -29,
    60516 => -29,
    60517 => -29,
    60518 => -29,
    60519 => -29,
    60520 => -29,
    60521 => -29,
    60522 => -29,
    60523 => -29,
    60524 => -29,
    60525 => -29,
    60526 => -29,
    60527 => -29,
    60528 => -29,
    60529 => -29,
    60530 => -29,
    60531 => -29,
    60532 => -29,
    60533 => -29,
    60534 => -29,
    60535 => -29,
    60536 => -29,
    60537 => -29,
    60538 => -29,
    60539 => -29,
    60540 => -29,
    60541 => -29,
    60542 => -29,
    60543 => -29,
    60544 => -29,
    60545 => -29,
    60546 => -29,
    60547 => -29,
    60548 => -29,
    60549 => -29,
    60550 => -29,
    60551 => -29,
    60552 => -29,
    60553 => -29,
    60554 => -29,
    60555 => -29,
    60556 => -29,
    60557 => -29,
    60558 => -29,
    60559 => -29,
    60560 => -29,
    60561 => -29,
    60562 => -29,
    60563 => -29,
    60564 => -29,
    60565 => -29,
    60566 => -29,
    60567 => -29,
    60568 => -29,
    60569 => -29,
    60570 => -29,
    60571 => -29,
    60572 => -29,
    60573 => -29,
    60574 => -29,
    60575 => -29,
    60576 => -29,
    60577 => -29,
    60578 => -29,
    60579 => -29,
    60580 => -29,
    60581 => -29,
    60582 => -29,
    60583 => -29,
    60584 => -29,
    60585 => -29,
    60586 => -29,
    60587 => -29,
    60588 => -29,
    60589 => -29,
    60590 => -29,
    60591 => -29,
    60592 => -29,
    60593 => -29,
    60594 => -29,
    60595 => -29,
    60596 => -29,
    60597 => -29,
    60598 => -29,
    60599 => -29,
    60600 => -29,
    60601 => -29,
    60602 => -29,
    60603 => -29,
    60604 => -29,
    60605 => -29,
    60606 => -29,
    60607 => -29,
    60608 => -29,
    60609 => -29,
    60610 => -29,
    60611 => -29,
    60612 => -29,
    60613 => -29,
    60614 => -29,
    60615 => -29,
    60616 => -29,
    60617 => -29,
    60618 => -29,
    60619 => -29,
    60620 => -29,
    60621 => -29,
    60622 => -29,
    60623 => -29,
    60624 => -29,
    60625 => -29,
    60626 => -29,
    60627 => -29,
    60628 => -29,
    60629 => -29,
    60630 => -29,
    60631 => -29,
    60632 => -29,
    60633 => -29,
    60634 => -29,
    60635 => -29,
    60636 => -29,
    60637 => -29,
    60638 => -29,
    60639 => -29,
    60640 => -28,
    60641 => -28,
    60642 => -28,
    60643 => -28,
    60644 => -28,
    60645 => -28,
    60646 => -28,
    60647 => -28,
    60648 => -28,
    60649 => -28,
    60650 => -28,
    60651 => -28,
    60652 => -28,
    60653 => -28,
    60654 => -28,
    60655 => -28,
    60656 => -28,
    60657 => -28,
    60658 => -28,
    60659 => -28,
    60660 => -28,
    60661 => -28,
    60662 => -28,
    60663 => -28,
    60664 => -28,
    60665 => -28,
    60666 => -28,
    60667 => -28,
    60668 => -28,
    60669 => -28,
    60670 => -28,
    60671 => -28,
    60672 => -28,
    60673 => -28,
    60674 => -28,
    60675 => -28,
    60676 => -28,
    60677 => -28,
    60678 => -28,
    60679 => -28,
    60680 => -28,
    60681 => -28,
    60682 => -28,
    60683 => -28,
    60684 => -28,
    60685 => -28,
    60686 => -28,
    60687 => -28,
    60688 => -28,
    60689 => -28,
    60690 => -28,
    60691 => -28,
    60692 => -28,
    60693 => -28,
    60694 => -28,
    60695 => -28,
    60696 => -28,
    60697 => -28,
    60698 => -28,
    60699 => -28,
    60700 => -28,
    60701 => -28,
    60702 => -28,
    60703 => -28,
    60704 => -28,
    60705 => -28,
    60706 => -28,
    60707 => -28,
    60708 => -28,
    60709 => -28,
    60710 => -28,
    60711 => -28,
    60712 => -28,
    60713 => -28,
    60714 => -28,
    60715 => -28,
    60716 => -28,
    60717 => -28,
    60718 => -28,
    60719 => -28,
    60720 => -28,
    60721 => -28,
    60722 => -28,
    60723 => -28,
    60724 => -28,
    60725 => -28,
    60726 => -28,
    60727 => -28,
    60728 => -28,
    60729 => -28,
    60730 => -28,
    60731 => -28,
    60732 => -28,
    60733 => -28,
    60734 => -28,
    60735 => -28,
    60736 => -28,
    60737 => -28,
    60738 => -28,
    60739 => -28,
    60740 => -28,
    60741 => -28,
    60742 => -28,
    60743 => -28,
    60744 => -28,
    60745 => -28,
    60746 => -28,
    60747 => -28,
    60748 => -28,
    60749 => -28,
    60750 => -28,
    60751 => -28,
    60752 => -28,
    60753 => -28,
    60754 => -28,
    60755 => -28,
    60756 => -28,
    60757 => -28,
    60758 => -28,
    60759 => -28,
    60760 => -28,
    60761 => -28,
    60762 => -28,
    60763 => -28,
    60764 => -28,
    60765 => -28,
    60766 => -28,
    60767 => -28,
    60768 => -28,
    60769 => -28,
    60770 => -28,
    60771 => -28,
    60772 => -28,
    60773 => -28,
    60774 => -28,
    60775 => -28,
    60776 => -28,
    60777 => -28,
    60778 => -28,
    60779 => -28,
    60780 => -28,
    60781 => -28,
    60782 => -28,
    60783 => -28,
    60784 => -28,
    60785 => -28,
    60786 => -28,
    60787 => -28,
    60788 => -28,
    60789 => -28,
    60790 => -28,
    60791 => -28,
    60792 => -28,
    60793 => -28,
    60794 => -28,
    60795 => -28,
    60796 => -28,
    60797 => -28,
    60798 => -28,
    60799 => -28,
    60800 => -28,
    60801 => -28,
    60802 => -28,
    60803 => -28,
    60804 => -28,
    60805 => -28,
    60806 => -28,
    60807 => -28,
    60808 => -28,
    60809 => -28,
    60810 => -28,
    60811 => -28,
    60812 => -28,
    60813 => -28,
    60814 => -28,
    60815 => -28,
    60816 => -28,
    60817 => -28,
    60818 => -28,
    60819 => -28,
    60820 => -28,
    60821 => -28,
    60822 => -28,
    60823 => -28,
    60824 => -28,
    60825 => -27,
    60826 => -27,
    60827 => -27,
    60828 => -27,
    60829 => -27,
    60830 => -27,
    60831 => -27,
    60832 => -27,
    60833 => -27,
    60834 => -27,
    60835 => -27,
    60836 => -27,
    60837 => -27,
    60838 => -27,
    60839 => -27,
    60840 => -27,
    60841 => -27,
    60842 => -27,
    60843 => -27,
    60844 => -27,
    60845 => -27,
    60846 => -27,
    60847 => -27,
    60848 => -27,
    60849 => -27,
    60850 => -27,
    60851 => -27,
    60852 => -27,
    60853 => -27,
    60854 => -27,
    60855 => -27,
    60856 => -27,
    60857 => -27,
    60858 => -27,
    60859 => -27,
    60860 => -27,
    60861 => -27,
    60862 => -27,
    60863 => -27,
    60864 => -27,
    60865 => -27,
    60866 => -27,
    60867 => -27,
    60868 => -27,
    60869 => -27,
    60870 => -27,
    60871 => -27,
    60872 => -27,
    60873 => -27,
    60874 => -27,
    60875 => -27,
    60876 => -27,
    60877 => -27,
    60878 => -27,
    60879 => -27,
    60880 => -27,
    60881 => -27,
    60882 => -27,
    60883 => -27,
    60884 => -27,
    60885 => -27,
    60886 => -27,
    60887 => -27,
    60888 => -27,
    60889 => -27,
    60890 => -27,
    60891 => -27,
    60892 => -27,
    60893 => -27,
    60894 => -27,
    60895 => -27,
    60896 => -27,
    60897 => -27,
    60898 => -27,
    60899 => -27,
    60900 => -27,
    60901 => -27,
    60902 => -27,
    60903 => -27,
    60904 => -27,
    60905 => -27,
    60906 => -27,
    60907 => -27,
    60908 => -27,
    60909 => -27,
    60910 => -27,
    60911 => -27,
    60912 => -27,
    60913 => -27,
    60914 => -27,
    60915 => -27,
    60916 => -27,
    60917 => -27,
    60918 => -27,
    60919 => -27,
    60920 => -27,
    60921 => -27,
    60922 => -27,
    60923 => -27,
    60924 => -27,
    60925 => -27,
    60926 => -27,
    60927 => -27,
    60928 => -27,
    60929 => -27,
    60930 => -27,
    60931 => -27,
    60932 => -27,
    60933 => -27,
    60934 => -27,
    60935 => -27,
    60936 => -27,
    60937 => -27,
    60938 => -27,
    60939 => -27,
    60940 => -27,
    60941 => -27,
    60942 => -27,
    60943 => -27,
    60944 => -27,
    60945 => -27,
    60946 => -27,
    60947 => -27,
    60948 => -27,
    60949 => -27,
    60950 => -27,
    60951 => -27,
    60952 => -27,
    60953 => -27,
    60954 => -27,
    60955 => -27,
    60956 => -27,
    60957 => -27,
    60958 => -27,
    60959 => -27,
    60960 => -27,
    60961 => -27,
    60962 => -27,
    60963 => -27,
    60964 => -27,
    60965 => -27,
    60966 => -27,
    60967 => -27,
    60968 => -27,
    60969 => -27,
    60970 => -27,
    60971 => -27,
    60972 => -27,
    60973 => -27,
    60974 => -27,
    60975 => -27,
    60976 => -27,
    60977 => -27,
    60978 => -27,
    60979 => -27,
    60980 => -27,
    60981 => -27,
    60982 => -27,
    60983 => -27,
    60984 => -27,
    60985 => -27,
    60986 => -27,
    60987 => -27,
    60988 => -27,
    60989 => -27,
    60990 => -27,
    60991 => -27,
    60992 => -27,
    60993 => -27,
    60994 => -27,
    60995 => -27,
    60996 => -27,
    60997 => -27,
    60998 => -27,
    60999 => -27,
    61000 => -27,
    61001 => -27,
    61002 => -27,
    61003 => -27,
    61004 => -27,
    61005 => -27,
    61006 => -27,
    61007 => -27,
    61008 => -26,
    61009 => -26,
    61010 => -26,
    61011 => -26,
    61012 => -26,
    61013 => -26,
    61014 => -26,
    61015 => -26,
    61016 => -26,
    61017 => -26,
    61018 => -26,
    61019 => -26,
    61020 => -26,
    61021 => -26,
    61022 => -26,
    61023 => -26,
    61024 => -26,
    61025 => -26,
    61026 => -26,
    61027 => -26,
    61028 => -26,
    61029 => -26,
    61030 => -26,
    61031 => -26,
    61032 => -26,
    61033 => -26,
    61034 => -26,
    61035 => -26,
    61036 => -26,
    61037 => -26,
    61038 => -26,
    61039 => -26,
    61040 => -26,
    61041 => -26,
    61042 => -26,
    61043 => -26,
    61044 => -26,
    61045 => -26,
    61046 => -26,
    61047 => -26,
    61048 => -26,
    61049 => -26,
    61050 => -26,
    61051 => -26,
    61052 => -26,
    61053 => -26,
    61054 => -26,
    61055 => -26,
    61056 => -26,
    61057 => -26,
    61058 => -26,
    61059 => -26,
    61060 => -26,
    61061 => -26,
    61062 => -26,
    61063 => -26,
    61064 => -26,
    61065 => -26,
    61066 => -26,
    61067 => -26,
    61068 => -26,
    61069 => -26,
    61070 => -26,
    61071 => -26,
    61072 => -26,
    61073 => -26,
    61074 => -26,
    61075 => -26,
    61076 => -26,
    61077 => -26,
    61078 => -26,
    61079 => -26,
    61080 => -26,
    61081 => -26,
    61082 => -26,
    61083 => -26,
    61084 => -26,
    61085 => -26,
    61086 => -26,
    61087 => -26,
    61088 => -26,
    61089 => -26,
    61090 => -26,
    61091 => -26,
    61092 => -26,
    61093 => -26,
    61094 => -26,
    61095 => -26,
    61096 => -26,
    61097 => -26,
    61098 => -26,
    61099 => -26,
    61100 => -26,
    61101 => -26,
    61102 => -26,
    61103 => -26,
    61104 => -26,
    61105 => -26,
    61106 => -26,
    61107 => -26,
    61108 => -26,
    61109 => -26,
    61110 => -26,
    61111 => -26,
    61112 => -26,
    61113 => -26,
    61114 => -26,
    61115 => -26,
    61116 => -26,
    61117 => -26,
    61118 => -26,
    61119 => -26,
    61120 => -26,
    61121 => -26,
    61122 => -26,
    61123 => -26,
    61124 => -26,
    61125 => -26,
    61126 => -26,
    61127 => -26,
    61128 => -26,
    61129 => -26,
    61130 => -26,
    61131 => -26,
    61132 => -26,
    61133 => -26,
    61134 => -26,
    61135 => -26,
    61136 => -26,
    61137 => -26,
    61138 => -26,
    61139 => -26,
    61140 => -26,
    61141 => -26,
    61142 => -26,
    61143 => -26,
    61144 => -26,
    61145 => -26,
    61146 => -26,
    61147 => -26,
    61148 => -26,
    61149 => -26,
    61150 => -26,
    61151 => -26,
    61152 => -26,
    61153 => -26,
    61154 => -26,
    61155 => -26,
    61156 => -26,
    61157 => -26,
    61158 => -26,
    61159 => -26,
    61160 => -26,
    61161 => -26,
    61162 => -26,
    61163 => -26,
    61164 => -26,
    61165 => -26,
    61166 => -26,
    61167 => -26,
    61168 => -26,
    61169 => -26,
    61170 => -26,
    61171 => -26,
    61172 => -26,
    61173 => -26,
    61174 => -26,
    61175 => -26,
    61176 => -26,
    61177 => -26,
    61178 => -26,
    61179 => -26,
    61180 => -26,
    61181 => -26,
    61182 => -26,
    61183 => -26,
    61184 => -26,
    61185 => -26,
    61186 => -26,
    61187 => -26,
    61188 => -26,
    61189 => -26,
    61190 => -25,
    61191 => -25,
    61192 => -25,
    61193 => -25,
    61194 => -25,
    61195 => -25,
    61196 => -25,
    61197 => -25,
    61198 => -25,
    61199 => -25,
    61200 => -25,
    61201 => -25,
    61202 => -25,
    61203 => -25,
    61204 => -25,
    61205 => -25,
    61206 => -25,
    61207 => -25,
    61208 => -25,
    61209 => -25,
    61210 => -25,
    61211 => -25,
    61212 => -25,
    61213 => -25,
    61214 => -25,
    61215 => -25,
    61216 => -25,
    61217 => -25,
    61218 => -25,
    61219 => -25,
    61220 => -25,
    61221 => -25,
    61222 => -25,
    61223 => -25,
    61224 => -25,
    61225 => -25,
    61226 => -25,
    61227 => -25,
    61228 => -25,
    61229 => -25,
    61230 => -25,
    61231 => -25,
    61232 => -25,
    61233 => -25,
    61234 => -25,
    61235 => -25,
    61236 => -25,
    61237 => -25,
    61238 => -25,
    61239 => -25,
    61240 => -25,
    61241 => -25,
    61242 => -25,
    61243 => -25,
    61244 => -25,
    61245 => -25,
    61246 => -25,
    61247 => -25,
    61248 => -25,
    61249 => -25,
    61250 => -25,
    61251 => -25,
    61252 => -25,
    61253 => -25,
    61254 => -25,
    61255 => -25,
    61256 => -25,
    61257 => -25,
    61258 => -25,
    61259 => -25,
    61260 => -25,
    61261 => -25,
    61262 => -25,
    61263 => -25,
    61264 => -25,
    61265 => -25,
    61266 => -25,
    61267 => -25,
    61268 => -25,
    61269 => -25,
    61270 => -25,
    61271 => -25,
    61272 => -25,
    61273 => -25,
    61274 => -25,
    61275 => -25,
    61276 => -25,
    61277 => -25,
    61278 => -25,
    61279 => -25,
    61280 => -25,
    61281 => -25,
    61282 => -25,
    61283 => -25,
    61284 => -25,
    61285 => -25,
    61286 => -25,
    61287 => -25,
    61288 => -25,
    61289 => -25,
    61290 => -25,
    61291 => -25,
    61292 => -25,
    61293 => -25,
    61294 => -25,
    61295 => -25,
    61296 => -25,
    61297 => -25,
    61298 => -25,
    61299 => -25,
    61300 => -25,
    61301 => -25,
    61302 => -25,
    61303 => -25,
    61304 => -25,
    61305 => -25,
    61306 => -25,
    61307 => -25,
    61308 => -25,
    61309 => -25,
    61310 => -25,
    61311 => -25,
    61312 => -25,
    61313 => -25,
    61314 => -25,
    61315 => -25,
    61316 => -25,
    61317 => -25,
    61318 => -25,
    61319 => -25,
    61320 => -25,
    61321 => -25,
    61322 => -25,
    61323 => -25,
    61324 => -25,
    61325 => -25,
    61326 => -25,
    61327 => -25,
    61328 => -25,
    61329 => -25,
    61330 => -25,
    61331 => -25,
    61332 => -25,
    61333 => -25,
    61334 => -25,
    61335 => -25,
    61336 => -25,
    61337 => -25,
    61338 => -25,
    61339 => -25,
    61340 => -25,
    61341 => -25,
    61342 => -25,
    61343 => -25,
    61344 => -25,
    61345 => -25,
    61346 => -25,
    61347 => -25,
    61348 => -25,
    61349 => -25,
    61350 => -25,
    61351 => -25,
    61352 => -25,
    61353 => -25,
    61354 => -25,
    61355 => -25,
    61356 => -25,
    61357 => -25,
    61358 => -25,
    61359 => -25,
    61360 => -25,
    61361 => -25,
    61362 => -25,
    61363 => -25,
    61364 => -25,
    61365 => -25,
    61366 => -25,
    61367 => -25,
    61368 => -25,
    61369 => -25,
    61370 => -24,
    61371 => -24,
    61372 => -24,
    61373 => -24,
    61374 => -24,
    61375 => -24,
    61376 => -24,
    61377 => -24,
    61378 => -24,
    61379 => -24,
    61380 => -24,
    61381 => -24,
    61382 => -24,
    61383 => -24,
    61384 => -24,
    61385 => -24,
    61386 => -24,
    61387 => -24,
    61388 => -24,
    61389 => -24,
    61390 => -24,
    61391 => -24,
    61392 => -24,
    61393 => -24,
    61394 => -24,
    61395 => -24,
    61396 => -24,
    61397 => -24,
    61398 => -24,
    61399 => -24,
    61400 => -24,
    61401 => -24,
    61402 => -24,
    61403 => -24,
    61404 => -24,
    61405 => -24,
    61406 => -24,
    61407 => -24,
    61408 => -24,
    61409 => -24,
    61410 => -24,
    61411 => -24,
    61412 => -24,
    61413 => -24,
    61414 => -24,
    61415 => -24,
    61416 => -24,
    61417 => -24,
    61418 => -24,
    61419 => -24,
    61420 => -24,
    61421 => -24,
    61422 => -24,
    61423 => -24,
    61424 => -24,
    61425 => -24,
    61426 => -24,
    61427 => -24,
    61428 => -24,
    61429 => -24,
    61430 => -24,
    61431 => -24,
    61432 => -24,
    61433 => -24,
    61434 => -24,
    61435 => -24,
    61436 => -24,
    61437 => -24,
    61438 => -24,
    61439 => -24,
    61440 => -24,
    61441 => -24,
    61442 => -24,
    61443 => -24,
    61444 => -24,
    61445 => -24,
    61446 => -24,
    61447 => -24,
    61448 => -24,
    61449 => -24,
    61450 => -24,
    61451 => -24,
    61452 => -24,
    61453 => -24,
    61454 => -24,
    61455 => -24,
    61456 => -24,
    61457 => -24,
    61458 => -24,
    61459 => -24,
    61460 => -24,
    61461 => -24,
    61462 => -24,
    61463 => -24,
    61464 => -24,
    61465 => -24,
    61466 => -24,
    61467 => -24,
    61468 => -24,
    61469 => -24,
    61470 => -24,
    61471 => -24,
    61472 => -24,
    61473 => -24,
    61474 => -24,
    61475 => -24,
    61476 => -24,
    61477 => -24,
    61478 => -24,
    61479 => -24,
    61480 => -24,
    61481 => -24,
    61482 => -24,
    61483 => -24,
    61484 => -24,
    61485 => -24,
    61486 => -24,
    61487 => -24,
    61488 => -24,
    61489 => -24,
    61490 => -24,
    61491 => -24,
    61492 => -24,
    61493 => -24,
    61494 => -24,
    61495 => -24,
    61496 => -24,
    61497 => -24,
    61498 => -24,
    61499 => -24,
    61500 => -24,
    61501 => -24,
    61502 => -24,
    61503 => -24,
    61504 => -24,
    61505 => -24,
    61506 => -24,
    61507 => -24,
    61508 => -24,
    61509 => -24,
    61510 => -24,
    61511 => -24,
    61512 => -24,
    61513 => -24,
    61514 => -24,
    61515 => -24,
    61516 => -24,
    61517 => -24,
    61518 => -24,
    61519 => -24,
    61520 => -24,
    61521 => -24,
    61522 => -24,
    61523 => -24,
    61524 => -24,
    61525 => -24,
    61526 => -24,
    61527 => -24,
    61528 => -24,
    61529 => -24,
    61530 => -24,
    61531 => -24,
    61532 => -24,
    61533 => -24,
    61534 => -24,
    61535 => -24,
    61536 => -24,
    61537 => -24,
    61538 => -24,
    61539 => -24,
    61540 => -24,
    61541 => -24,
    61542 => -24,
    61543 => -24,
    61544 => -24,
    61545 => -24,
    61546 => -24,
    61547 => -24,
    61548 => -24,
    61549 => -23,
    61550 => -23,
    61551 => -23,
    61552 => -23,
    61553 => -23,
    61554 => -23,
    61555 => -23,
    61556 => -23,
    61557 => -23,
    61558 => -23,
    61559 => -23,
    61560 => -23,
    61561 => -23,
    61562 => -23,
    61563 => -23,
    61564 => -23,
    61565 => -23,
    61566 => -23,
    61567 => -23,
    61568 => -23,
    61569 => -23,
    61570 => -23,
    61571 => -23,
    61572 => -23,
    61573 => -23,
    61574 => -23,
    61575 => -23,
    61576 => -23,
    61577 => -23,
    61578 => -23,
    61579 => -23,
    61580 => -23,
    61581 => -23,
    61582 => -23,
    61583 => -23,
    61584 => -23,
    61585 => -23,
    61586 => -23,
    61587 => -23,
    61588 => -23,
    61589 => -23,
    61590 => -23,
    61591 => -23,
    61592 => -23,
    61593 => -23,
    61594 => -23,
    61595 => -23,
    61596 => -23,
    61597 => -23,
    61598 => -23,
    61599 => -23,
    61600 => -23,
    61601 => -23,
    61602 => -23,
    61603 => -23,
    61604 => -23,
    61605 => -23,
    61606 => -23,
    61607 => -23,
    61608 => -23,
    61609 => -23,
    61610 => -23,
    61611 => -23,
    61612 => -23,
    61613 => -23,
    61614 => -23,
    61615 => -23,
    61616 => -23,
    61617 => -23,
    61618 => -23,
    61619 => -23,
    61620 => -23,
    61621 => -23,
    61622 => -23,
    61623 => -23,
    61624 => -23,
    61625 => -23,
    61626 => -23,
    61627 => -23,
    61628 => -23,
    61629 => -23,
    61630 => -23,
    61631 => -23,
    61632 => -23,
    61633 => -23,
    61634 => -23,
    61635 => -23,
    61636 => -23,
    61637 => -23,
    61638 => -23,
    61639 => -23,
    61640 => -23,
    61641 => -23,
    61642 => -23,
    61643 => -23,
    61644 => -23,
    61645 => -23,
    61646 => -23,
    61647 => -23,
    61648 => -23,
    61649 => -23,
    61650 => -23,
    61651 => -23,
    61652 => -23,
    61653 => -23,
    61654 => -23,
    61655 => -23,
    61656 => -23,
    61657 => -23,
    61658 => -23,
    61659 => -23,
    61660 => -23,
    61661 => -23,
    61662 => -23,
    61663 => -23,
    61664 => -23,
    61665 => -23,
    61666 => -23,
    61667 => -23,
    61668 => -23,
    61669 => -23,
    61670 => -23,
    61671 => -23,
    61672 => -23,
    61673 => -23,
    61674 => -23,
    61675 => -23,
    61676 => -23,
    61677 => -23,
    61678 => -23,
    61679 => -23,
    61680 => -23,
    61681 => -23,
    61682 => -23,
    61683 => -23,
    61684 => -23,
    61685 => -23,
    61686 => -23,
    61687 => -23,
    61688 => -23,
    61689 => -23,
    61690 => -23,
    61691 => -23,
    61692 => -23,
    61693 => -23,
    61694 => -23,
    61695 => -23,
    61696 => -23,
    61697 => -23,
    61698 => -23,
    61699 => -23,
    61700 => -23,
    61701 => -23,
    61702 => -23,
    61703 => -23,
    61704 => -23,
    61705 => -23,
    61706 => -23,
    61707 => -23,
    61708 => -23,
    61709 => -23,
    61710 => -23,
    61711 => -23,
    61712 => -23,
    61713 => -23,
    61714 => -23,
    61715 => -23,
    61716 => -23,
    61717 => -23,
    61718 => -23,
    61719 => -23,
    61720 => -23,
    61721 => -23,
    61722 => -23,
    61723 => -23,
    61724 => -23,
    61725 => -23,
    61726 => -23,
    61727 => -22,
    61728 => -22,
    61729 => -22,
    61730 => -22,
    61731 => -22,
    61732 => -22,
    61733 => -22,
    61734 => -22,
    61735 => -22,
    61736 => -22,
    61737 => -22,
    61738 => -22,
    61739 => -22,
    61740 => -22,
    61741 => -22,
    61742 => -22,
    61743 => -22,
    61744 => -22,
    61745 => -22,
    61746 => -22,
    61747 => -22,
    61748 => -22,
    61749 => -22,
    61750 => -22,
    61751 => -22,
    61752 => -22,
    61753 => -22,
    61754 => -22,
    61755 => -22,
    61756 => -22,
    61757 => -22,
    61758 => -22,
    61759 => -22,
    61760 => -22,
    61761 => -22,
    61762 => -22,
    61763 => -22,
    61764 => -22,
    61765 => -22,
    61766 => -22,
    61767 => -22,
    61768 => -22,
    61769 => -22,
    61770 => -22,
    61771 => -22,
    61772 => -22,
    61773 => -22,
    61774 => -22,
    61775 => -22,
    61776 => -22,
    61777 => -22,
    61778 => -22,
    61779 => -22,
    61780 => -22,
    61781 => -22,
    61782 => -22,
    61783 => -22,
    61784 => -22,
    61785 => -22,
    61786 => -22,
    61787 => -22,
    61788 => -22,
    61789 => -22,
    61790 => -22,
    61791 => -22,
    61792 => -22,
    61793 => -22,
    61794 => -22,
    61795 => -22,
    61796 => -22,
    61797 => -22,
    61798 => -22,
    61799 => -22,
    61800 => -22,
    61801 => -22,
    61802 => -22,
    61803 => -22,
    61804 => -22,
    61805 => -22,
    61806 => -22,
    61807 => -22,
    61808 => -22,
    61809 => -22,
    61810 => -22,
    61811 => -22,
    61812 => -22,
    61813 => -22,
    61814 => -22,
    61815 => -22,
    61816 => -22,
    61817 => -22,
    61818 => -22,
    61819 => -22,
    61820 => -22,
    61821 => -22,
    61822 => -22,
    61823 => -22,
    61824 => -22,
    61825 => -22,
    61826 => -22,
    61827 => -22,
    61828 => -22,
    61829 => -22,
    61830 => -22,
    61831 => -22,
    61832 => -22,
    61833 => -22,
    61834 => -22,
    61835 => -22,
    61836 => -22,
    61837 => -22,
    61838 => -22,
    61839 => -22,
    61840 => -22,
    61841 => -22,
    61842 => -22,
    61843 => -22,
    61844 => -22,
    61845 => -22,
    61846 => -22,
    61847 => -22,
    61848 => -22,
    61849 => -22,
    61850 => -22,
    61851 => -22,
    61852 => -22,
    61853 => -22,
    61854 => -22,
    61855 => -22,
    61856 => -22,
    61857 => -22,
    61858 => -22,
    61859 => -22,
    61860 => -22,
    61861 => -22,
    61862 => -22,
    61863 => -22,
    61864 => -22,
    61865 => -22,
    61866 => -22,
    61867 => -22,
    61868 => -22,
    61869 => -22,
    61870 => -22,
    61871 => -22,
    61872 => -22,
    61873 => -22,
    61874 => -22,
    61875 => -22,
    61876 => -22,
    61877 => -22,
    61878 => -22,
    61879 => -22,
    61880 => -22,
    61881 => -22,
    61882 => -22,
    61883 => -22,
    61884 => -22,
    61885 => -22,
    61886 => -22,
    61887 => -22,
    61888 => -22,
    61889 => -22,
    61890 => -22,
    61891 => -22,
    61892 => -22,
    61893 => -22,
    61894 => -22,
    61895 => -22,
    61896 => -22,
    61897 => -22,
    61898 => -22,
    61899 => -22,
    61900 => -22,
    61901 => -22,
    61902 => -22,
    61903 => -22,
    61904 => -21,
    61905 => -21,
    61906 => -21,
    61907 => -21,
    61908 => -21,
    61909 => -21,
    61910 => -21,
    61911 => -21,
    61912 => -21,
    61913 => -21,
    61914 => -21,
    61915 => -21,
    61916 => -21,
    61917 => -21,
    61918 => -21,
    61919 => -21,
    61920 => -21,
    61921 => -21,
    61922 => -21,
    61923 => -21,
    61924 => -21,
    61925 => -21,
    61926 => -21,
    61927 => -21,
    61928 => -21,
    61929 => -21,
    61930 => -21,
    61931 => -21,
    61932 => -21,
    61933 => -21,
    61934 => -21,
    61935 => -21,
    61936 => -21,
    61937 => -21,
    61938 => -21,
    61939 => -21,
    61940 => -21,
    61941 => -21,
    61942 => -21,
    61943 => -21,
    61944 => -21,
    61945 => -21,
    61946 => -21,
    61947 => -21,
    61948 => -21,
    61949 => -21,
    61950 => -21,
    61951 => -21,
    61952 => -21,
    61953 => -21,
    61954 => -21,
    61955 => -21,
    61956 => -21,
    61957 => -21,
    61958 => -21,
    61959 => -21,
    61960 => -21,
    61961 => -21,
    61962 => -21,
    61963 => -21,
    61964 => -21,
    61965 => -21,
    61966 => -21,
    61967 => -21,
    61968 => -21,
    61969 => -21,
    61970 => -21,
    61971 => -21,
    61972 => -21,
    61973 => -21,
    61974 => -21,
    61975 => -21,
    61976 => -21,
    61977 => -21,
    61978 => -21,
    61979 => -21,
    61980 => -21,
    61981 => -21,
    61982 => -21,
    61983 => -21,
    61984 => -21,
    61985 => -21,
    61986 => -21,
    61987 => -21,
    61988 => -21,
    61989 => -21,
    61990 => -21,
    61991 => -21,
    61992 => -21,
    61993 => -21,
    61994 => -21,
    61995 => -21,
    61996 => -21,
    61997 => -21,
    61998 => -21,
    61999 => -21,
    62000 => -21,
    62001 => -21,
    62002 => -21,
    62003 => -21,
    62004 => -21,
    62005 => -21,
    62006 => -21,
    62007 => -21,
    62008 => -21,
    62009 => -21,
    62010 => -21,
    62011 => -21,
    62012 => -21,
    62013 => -21,
    62014 => -21,
    62015 => -21,
    62016 => -21,
    62017 => -21,
    62018 => -21,
    62019 => -21,
    62020 => -21,
    62021 => -21,
    62022 => -21,
    62023 => -21,
    62024 => -21,
    62025 => -21,
    62026 => -21,
    62027 => -21,
    62028 => -21,
    62029 => -21,
    62030 => -21,
    62031 => -21,
    62032 => -21,
    62033 => -21,
    62034 => -21,
    62035 => -21,
    62036 => -21,
    62037 => -21,
    62038 => -21,
    62039 => -21,
    62040 => -21,
    62041 => -21,
    62042 => -21,
    62043 => -21,
    62044 => -21,
    62045 => -21,
    62046 => -21,
    62047 => -21,
    62048 => -21,
    62049 => -21,
    62050 => -21,
    62051 => -21,
    62052 => -21,
    62053 => -21,
    62054 => -21,
    62055 => -21,
    62056 => -21,
    62057 => -21,
    62058 => -21,
    62059 => -21,
    62060 => -21,
    62061 => -21,
    62062 => -21,
    62063 => -21,
    62064 => -21,
    62065 => -21,
    62066 => -21,
    62067 => -21,
    62068 => -21,
    62069 => -21,
    62070 => -21,
    62071 => -21,
    62072 => -21,
    62073 => -21,
    62074 => -21,
    62075 => -21,
    62076 => -21,
    62077 => -21,
    62078 => -21,
    62079 => -21,
    62080 => -20,
    62081 => -20,
    62082 => -20,
    62083 => -20,
    62084 => -20,
    62085 => -20,
    62086 => -20,
    62087 => -20,
    62088 => -20,
    62089 => -20,
    62090 => -20,
    62091 => -20,
    62092 => -20,
    62093 => -20,
    62094 => -20,
    62095 => -20,
    62096 => -20,
    62097 => -20,
    62098 => -20,
    62099 => -20,
    62100 => -20,
    62101 => -20,
    62102 => -20,
    62103 => -20,
    62104 => -20,
    62105 => -20,
    62106 => -20,
    62107 => -20,
    62108 => -20,
    62109 => -20,
    62110 => -20,
    62111 => -20,
    62112 => -20,
    62113 => -20,
    62114 => -20,
    62115 => -20,
    62116 => -20,
    62117 => -20,
    62118 => -20,
    62119 => -20,
    62120 => -20,
    62121 => -20,
    62122 => -20,
    62123 => -20,
    62124 => -20,
    62125 => -20,
    62126 => -20,
    62127 => -20,
    62128 => -20,
    62129 => -20,
    62130 => -20,
    62131 => -20,
    62132 => -20,
    62133 => -20,
    62134 => -20,
    62135 => -20,
    62136 => -20,
    62137 => -20,
    62138 => -20,
    62139 => -20,
    62140 => -20,
    62141 => -20,
    62142 => -20,
    62143 => -20,
    62144 => -20,
    62145 => -20,
    62146 => -20,
    62147 => -20,
    62148 => -20,
    62149 => -20,
    62150 => -20,
    62151 => -20,
    62152 => -20,
    62153 => -20,
    62154 => -20,
    62155 => -20,
    62156 => -20,
    62157 => -20,
    62158 => -20,
    62159 => -20,
    62160 => -20,
    62161 => -20,
    62162 => -20,
    62163 => -20,
    62164 => -20,
    62165 => -20,
    62166 => -20,
    62167 => -20,
    62168 => -20,
    62169 => -20,
    62170 => -20,
    62171 => -20,
    62172 => -20,
    62173 => -20,
    62174 => -20,
    62175 => -20,
    62176 => -20,
    62177 => -20,
    62178 => -20,
    62179 => -20,
    62180 => -20,
    62181 => -20,
    62182 => -20,
    62183 => -20,
    62184 => -20,
    62185 => -20,
    62186 => -20,
    62187 => -20,
    62188 => -20,
    62189 => -20,
    62190 => -20,
    62191 => -20,
    62192 => -20,
    62193 => -20,
    62194 => -20,
    62195 => -20,
    62196 => -20,
    62197 => -20,
    62198 => -20,
    62199 => -20,
    62200 => -20,
    62201 => -20,
    62202 => -20,
    62203 => -20,
    62204 => -20,
    62205 => -20,
    62206 => -20,
    62207 => -20,
    62208 => -20,
    62209 => -20,
    62210 => -20,
    62211 => -20,
    62212 => -20,
    62213 => -20,
    62214 => -20,
    62215 => -20,
    62216 => -20,
    62217 => -20,
    62218 => -20,
    62219 => -20,
    62220 => -20,
    62221 => -20,
    62222 => -20,
    62223 => -20,
    62224 => -20,
    62225 => -20,
    62226 => -20,
    62227 => -20,
    62228 => -20,
    62229 => -20,
    62230 => -20,
    62231 => -20,
    62232 => -20,
    62233 => -20,
    62234 => -20,
    62235 => -20,
    62236 => -20,
    62237 => -20,
    62238 => -20,
    62239 => -20,
    62240 => -20,
    62241 => -20,
    62242 => -20,
    62243 => -20,
    62244 => -20,
    62245 => -20,
    62246 => -20,
    62247 => -20,
    62248 => -20,
    62249 => -20,
    62250 => -20,
    62251 => -20,
    62252 => -20,
    62253 => -20,
    62254 => -19,
    62255 => -19,
    62256 => -19,
    62257 => -19,
    62258 => -19,
    62259 => -19,
    62260 => -19,
    62261 => -19,
    62262 => -19,
    62263 => -19,
    62264 => -19,
    62265 => -19,
    62266 => -19,
    62267 => -19,
    62268 => -19,
    62269 => -19,
    62270 => -19,
    62271 => -19,
    62272 => -19,
    62273 => -19,
    62274 => -19,
    62275 => -19,
    62276 => -19,
    62277 => -19,
    62278 => -19,
    62279 => -19,
    62280 => -19,
    62281 => -19,
    62282 => -19,
    62283 => -19,
    62284 => -19,
    62285 => -19,
    62286 => -19,
    62287 => -19,
    62288 => -19,
    62289 => -19,
    62290 => -19,
    62291 => -19,
    62292 => -19,
    62293 => -19,
    62294 => -19,
    62295 => -19,
    62296 => -19,
    62297 => -19,
    62298 => -19,
    62299 => -19,
    62300 => -19,
    62301 => -19,
    62302 => -19,
    62303 => -19,
    62304 => -19,
    62305 => -19,
    62306 => -19,
    62307 => -19,
    62308 => -19,
    62309 => -19,
    62310 => -19,
    62311 => -19,
    62312 => -19,
    62313 => -19,
    62314 => -19,
    62315 => -19,
    62316 => -19,
    62317 => -19,
    62318 => -19,
    62319 => -19,
    62320 => -19,
    62321 => -19,
    62322 => -19,
    62323 => -19,
    62324 => -19,
    62325 => -19,
    62326 => -19,
    62327 => -19,
    62328 => -19,
    62329 => -19,
    62330 => -19,
    62331 => -19,
    62332 => -19,
    62333 => -19,
    62334 => -19,
    62335 => -19,
    62336 => -19,
    62337 => -19,
    62338 => -19,
    62339 => -19,
    62340 => -19,
    62341 => -19,
    62342 => -19,
    62343 => -19,
    62344 => -19,
    62345 => -19,
    62346 => -19,
    62347 => -19,
    62348 => -19,
    62349 => -19,
    62350 => -19,
    62351 => -19,
    62352 => -19,
    62353 => -19,
    62354 => -19,
    62355 => -19,
    62356 => -19,
    62357 => -19,
    62358 => -19,
    62359 => -19,
    62360 => -19,
    62361 => -19,
    62362 => -19,
    62363 => -19,
    62364 => -19,
    62365 => -19,
    62366 => -19,
    62367 => -19,
    62368 => -19,
    62369 => -19,
    62370 => -19,
    62371 => -19,
    62372 => -19,
    62373 => -19,
    62374 => -19,
    62375 => -19,
    62376 => -19,
    62377 => -19,
    62378 => -19,
    62379 => -19,
    62380 => -19,
    62381 => -19,
    62382 => -19,
    62383 => -19,
    62384 => -19,
    62385 => -19,
    62386 => -19,
    62387 => -19,
    62388 => -19,
    62389 => -19,
    62390 => -19,
    62391 => -19,
    62392 => -19,
    62393 => -19,
    62394 => -19,
    62395 => -19,
    62396 => -19,
    62397 => -19,
    62398 => -19,
    62399 => -19,
    62400 => -19,
    62401 => -19,
    62402 => -19,
    62403 => -19,
    62404 => -19,
    62405 => -19,
    62406 => -19,
    62407 => -19,
    62408 => -19,
    62409 => -19,
    62410 => -19,
    62411 => -19,
    62412 => -19,
    62413 => -19,
    62414 => -19,
    62415 => -19,
    62416 => -19,
    62417 => -19,
    62418 => -19,
    62419 => -19,
    62420 => -19,
    62421 => -19,
    62422 => -19,
    62423 => -19,
    62424 => -19,
    62425 => -19,
    62426 => -19,
    62427 => -19,
    62428 => -18,
    62429 => -18,
    62430 => -18,
    62431 => -18,
    62432 => -18,
    62433 => -18,
    62434 => -18,
    62435 => -18,
    62436 => -18,
    62437 => -18,
    62438 => -18,
    62439 => -18,
    62440 => -18,
    62441 => -18,
    62442 => -18,
    62443 => -18,
    62444 => -18,
    62445 => -18,
    62446 => -18,
    62447 => -18,
    62448 => -18,
    62449 => -18,
    62450 => -18,
    62451 => -18,
    62452 => -18,
    62453 => -18,
    62454 => -18,
    62455 => -18,
    62456 => -18,
    62457 => -18,
    62458 => -18,
    62459 => -18,
    62460 => -18,
    62461 => -18,
    62462 => -18,
    62463 => -18,
    62464 => -18,
    62465 => -18,
    62466 => -18,
    62467 => -18,
    62468 => -18,
    62469 => -18,
    62470 => -18,
    62471 => -18,
    62472 => -18,
    62473 => -18,
    62474 => -18,
    62475 => -18,
    62476 => -18,
    62477 => -18,
    62478 => -18,
    62479 => -18,
    62480 => -18,
    62481 => -18,
    62482 => -18,
    62483 => -18,
    62484 => -18,
    62485 => -18,
    62486 => -18,
    62487 => -18,
    62488 => -18,
    62489 => -18,
    62490 => -18,
    62491 => -18,
    62492 => -18,
    62493 => -18,
    62494 => -18,
    62495 => -18,
    62496 => -18,
    62497 => -18,
    62498 => -18,
    62499 => -18,
    62500 => -18,
    62501 => -18,
    62502 => -18,
    62503 => -18,
    62504 => -18,
    62505 => -18,
    62506 => -18,
    62507 => -18,
    62508 => -18,
    62509 => -18,
    62510 => -18,
    62511 => -18,
    62512 => -18,
    62513 => -18,
    62514 => -18,
    62515 => -18,
    62516 => -18,
    62517 => -18,
    62518 => -18,
    62519 => -18,
    62520 => -18,
    62521 => -18,
    62522 => -18,
    62523 => -18,
    62524 => -18,
    62525 => -18,
    62526 => -18,
    62527 => -18,
    62528 => -18,
    62529 => -18,
    62530 => -18,
    62531 => -18,
    62532 => -18,
    62533 => -18,
    62534 => -18,
    62535 => -18,
    62536 => -18,
    62537 => -18,
    62538 => -18,
    62539 => -18,
    62540 => -18,
    62541 => -18,
    62542 => -18,
    62543 => -18,
    62544 => -18,
    62545 => -18,
    62546 => -18,
    62547 => -18,
    62548 => -18,
    62549 => -18,
    62550 => -18,
    62551 => -18,
    62552 => -18,
    62553 => -18,
    62554 => -18,
    62555 => -18,
    62556 => -18,
    62557 => -18,
    62558 => -18,
    62559 => -18,
    62560 => -18,
    62561 => -18,
    62562 => -18,
    62563 => -18,
    62564 => -18,
    62565 => -18,
    62566 => -18,
    62567 => -18,
    62568 => -18,
    62569 => -18,
    62570 => -18,
    62571 => -18,
    62572 => -18,
    62573 => -18,
    62574 => -18,
    62575 => -18,
    62576 => -18,
    62577 => -18,
    62578 => -18,
    62579 => -18,
    62580 => -18,
    62581 => -18,
    62582 => -18,
    62583 => -18,
    62584 => -18,
    62585 => -18,
    62586 => -18,
    62587 => -18,
    62588 => -18,
    62589 => -18,
    62590 => -18,
    62591 => -18,
    62592 => -18,
    62593 => -18,
    62594 => -18,
    62595 => -18,
    62596 => -18,
    62597 => -18,
    62598 => -18,
    62599 => -18,
    62600 => -18,
    62601 => -17,
    62602 => -17,
    62603 => -17,
    62604 => -17,
    62605 => -17,
    62606 => -17,
    62607 => -17,
    62608 => -17,
    62609 => -17,
    62610 => -17,
    62611 => -17,
    62612 => -17,
    62613 => -17,
    62614 => -17,
    62615 => -17,
    62616 => -17,
    62617 => -17,
    62618 => -17,
    62619 => -17,
    62620 => -17,
    62621 => -17,
    62622 => -17,
    62623 => -17,
    62624 => -17,
    62625 => -17,
    62626 => -17,
    62627 => -17,
    62628 => -17,
    62629 => -17,
    62630 => -17,
    62631 => -17,
    62632 => -17,
    62633 => -17,
    62634 => -17,
    62635 => -17,
    62636 => -17,
    62637 => -17,
    62638 => -17,
    62639 => -17,
    62640 => -17,
    62641 => -17,
    62642 => -17,
    62643 => -17,
    62644 => -17,
    62645 => -17,
    62646 => -17,
    62647 => -17,
    62648 => -17,
    62649 => -17,
    62650 => -17,
    62651 => -17,
    62652 => -17,
    62653 => -17,
    62654 => -17,
    62655 => -17,
    62656 => -17,
    62657 => -17,
    62658 => -17,
    62659 => -17,
    62660 => -17,
    62661 => -17,
    62662 => -17,
    62663 => -17,
    62664 => -17,
    62665 => -17,
    62666 => -17,
    62667 => -17,
    62668 => -17,
    62669 => -17,
    62670 => -17,
    62671 => -17,
    62672 => -17,
    62673 => -17,
    62674 => -17,
    62675 => -17,
    62676 => -17,
    62677 => -17,
    62678 => -17,
    62679 => -17,
    62680 => -17,
    62681 => -17,
    62682 => -17,
    62683 => -17,
    62684 => -17,
    62685 => -17,
    62686 => -17,
    62687 => -17,
    62688 => -17,
    62689 => -17,
    62690 => -17,
    62691 => -17,
    62692 => -17,
    62693 => -17,
    62694 => -17,
    62695 => -17,
    62696 => -17,
    62697 => -17,
    62698 => -17,
    62699 => -17,
    62700 => -17,
    62701 => -17,
    62702 => -17,
    62703 => -17,
    62704 => -17,
    62705 => -17,
    62706 => -17,
    62707 => -17,
    62708 => -17,
    62709 => -17,
    62710 => -17,
    62711 => -17,
    62712 => -17,
    62713 => -17,
    62714 => -17,
    62715 => -17,
    62716 => -17,
    62717 => -17,
    62718 => -17,
    62719 => -17,
    62720 => -17,
    62721 => -17,
    62722 => -17,
    62723 => -17,
    62724 => -17,
    62725 => -17,
    62726 => -17,
    62727 => -17,
    62728 => -17,
    62729 => -17,
    62730 => -17,
    62731 => -17,
    62732 => -17,
    62733 => -17,
    62734 => -17,
    62735 => -17,
    62736 => -17,
    62737 => -17,
    62738 => -17,
    62739 => -17,
    62740 => -17,
    62741 => -17,
    62742 => -17,
    62743 => -17,
    62744 => -17,
    62745 => -17,
    62746 => -17,
    62747 => -17,
    62748 => -17,
    62749 => -17,
    62750 => -17,
    62751 => -17,
    62752 => -17,
    62753 => -17,
    62754 => -17,
    62755 => -17,
    62756 => -17,
    62757 => -17,
    62758 => -17,
    62759 => -17,
    62760 => -17,
    62761 => -17,
    62762 => -17,
    62763 => -17,
    62764 => -17,
    62765 => -17,
    62766 => -17,
    62767 => -17,
    62768 => -17,
    62769 => -17,
    62770 => -17,
    62771 => -17,
    62772 => -16,
    62773 => -16,
    62774 => -16,
    62775 => -16,
    62776 => -16,
    62777 => -16,
    62778 => -16,
    62779 => -16,
    62780 => -16,
    62781 => -16,
    62782 => -16,
    62783 => -16,
    62784 => -16,
    62785 => -16,
    62786 => -16,
    62787 => -16,
    62788 => -16,
    62789 => -16,
    62790 => -16,
    62791 => -16,
    62792 => -16,
    62793 => -16,
    62794 => -16,
    62795 => -16,
    62796 => -16,
    62797 => -16,
    62798 => -16,
    62799 => -16,
    62800 => -16,
    62801 => -16,
    62802 => -16,
    62803 => -16,
    62804 => -16,
    62805 => -16,
    62806 => -16,
    62807 => -16,
    62808 => -16,
    62809 => -16,
    62810 => -16,
    62811 => -16,
    62812 => -16,
    62813 => -16,
    62814 => -16,
    62815 => -16,
    62816 => -16,
    62817 => -16,
    62818 => -16,
    62819 => -16,
    62820 => -16,
    62821 => -16,
    62822 => -16,
    62823 => -16,
    62824 => -16,
    62825 => -16,
    62826 => -16,
    62827 => -16,
    62828 => -16,
    62829 => -16,
    62830 => -16,
    62831 => -16,
    62832 => -16,
    62833 => -16,
    62834 => -16,
    62835 => -16,
    62836 => -16,
    62837 => -16,
    62838 => -16,
    62839 => -16,
    62840 => -16,
    62841 => -16,
    62842 => -16,
    62843 => -16,
    62844 => -16,
    62845 => -16,
    62846 => -16,
    62847 => -16,
    62848 => -16,
    62849 => -16,
    62850 => -16,
    62851 => -16,
    62852 => -16,
    62853 => -16,
    62854 => -16,
    62855 => -16,
    62856 => -16,
    62857 => -16,
    62858 => -16,
    62859 => -16,
    62860 => -16,
    62861 => -16,
    62862 => -16,
    62863 => -16,
    62864 => -16,
    62865 => -16,
    62866 => -16,
    62867 => -16,
    62868 => -16,
    62869 => -16,
    62870 => -16,
    62871 => -16,
    62872 => -16,
    62873 => -16,
    62874 => -16,
    62875 => -16,
    62876 => -16,
    62877 => -16,
    62878 => -16,
    62879 => -16,
    62880 => -16,
    62881 => -16,
    62882 => -16,
    62883 => -16,
    62884 => -16,
    62885 => -16,
    62886 => -16,
    62887 => -16,
    62888 => -16,
    62889 => -16,
    62890 => -16,
    62891 => -16,
    62892 => -16,
    62893 => -16,
    62894 => -16,
    62895 => -16,
    62896 => -16,
    62897 => -16,
    62898 => -16,
    62899 => -16,
    62900 => -16,
    62901 => -16,
    62902 => -16,
    62903 => -16,
    62904 => -16,
    62905 => -16,
    62906 => -16,
    62907 => -16,
    62908 => -16,
    62909 => -16,
    62910 => -16,
    62911 => -16,
    62912 => -16,
    62913 => -16,
    62914 => -16,
    62915 => -16,
    62916 => -16,
    62917 => -16,
    62918 => -16,
    62919 => -16,
    62920 => -16,
    62921 => -16,
    62922 => -16,
    62923 => -16,
    62924 => -16,
    62925 => -16,
    62926 => -16,
    62927 => -16,
    62928 => -16,
    62929 => -16,
    62930 => -16,
    62931 => -16,
    62932 => -16,
    62933 => -16,
    62934 => -16,
    62935 => -16,
    62936 => -16,
    62937 => -16,
    62938 => -16,
    62939 => -16,
    62940 => -16,
    62941 => -16,
    62942 => -16,
    62943 => -16,
    62944 => -15,
    62945 => -15,
    62946 => -15,
    62947 => -15,
    62948 => -15,
    62949 => -15,
    62950 => -15,
    62951 => -15,
    62952 => -15,
    62953 => -15,
    62954 => -15,
    62955 => -15,
    62956 => -15,
    62957 => -15,
    62958 => -15,
    62959 => -15,
    62960 => -15,
    62961 => -15,
    62962 => -15,
    62963 => -15,
    62964 => -15,
    62965 => -15,
    62966 => -15,
    62967 => -15,
    62968 => -15,
    62969 => -15,
    62970 => -15,
    62971 => -15,
    62972 => -15,
    62973 => -15,
    62974 => -15,
    62975 => -15,
    62976 => -15,
    62977 => -15,
    62978 => -15,
    62979 => -15,
    62980 => -15,
    62981 => -15,
    62982 => -15,
    62983 => -15,
    62984 => -15,
    62985 => -15,
    62986 => -15,
    62987 => -15,
    62988 => -15,
    62989 => -15,
    62990 => -15,
    62991 => -15,
    62992 => -15,
    62993 => -15,
    62994 => -15,
    62995 => -15,
    62996 => -15,
    62997 => -15,
    62998 => -15,
    62999 => -15,
    63000 => -15,
    63001 => -15,
    63002 => -15,
    63003 => -15,
    63004 => -15,
    63005 => -15,
    63006 => -15,
    63007 => -15,
    63008 => -15,
    63009 => -15,
    63010 => -15,
    63011 => -15,
    63012 => -15,
    63013 => -15,
    63014 => -15,
    63015 => -15,
    63016 => -15,
    63017 => -15,
    63018 => -15,
    63019 => -15,
    63020 => -15,
    63021 => -15,
    63022 => -15,
    63023 => -15,
    63024 => -15,
    63025 => -15,
    63026 => -15,
    63027 => -15,
    63028 => -15,
    63029 => -15,
    63030 => -15,
    63031 => -15,
    63032 => -15,
    63033 => -15,
    63034 => -15,
    63035 => -15,
    63036 => -15,
    63037 => -15,
    63038 => -15,
    63039 => -15,
    63040 => -15,
    63041 => -15,
    63042 => -15,
    63043 => -15,
    63044 => -15,
    63045 => -15,
    63046 => -15,
    63047 => -15,
    63048 => -15,
    63049 => -15,
    63050 => -15,
    63051 => -15,
    63052 => -15,
    63053 => -15,
    63054 => -15,
    63055 => -15,
    63056 => -15,
    63057 => -15,
    63058 => -15,
    63059 => -15,
    63060 => -15,
    63061 => -15,
    63062 => -15,
    63063 => -15,
    63064 => -15,
    63065 => -15,
    63066 => -15,
    63067 => -15,
    63068 => -15,
    63069 => -15,
    63070 => -15,
    63071 => -15,
    63072 => -15,
    63073 => -15,
    63074 => -15,
    63075 => -15,
    63076 => -15,
    63077 => -15,
    63078 => -15,
    63079 => -15,
    63080 => -15,
    63081 => -15,
    63082 => -15,
    63083 => -15,
    63084 => -15,
    63085 => -15,
    63086 => -15,
    63087 => -15,
    63088 => -15,
    63089 => -15,
    63090 => -15,
    63091 => -15,
    63092 => -15,
    63093 => -15,
    63094 => -15,
    63095 => -15,
    63096 => -15,
    63097 => -15,
    63098 => -15,
    63099 => -15,
    63100 => -15,
    63101 => -15,
    63102 => -15,
    63103 => -15,
    63104 => -15,
    63105 => -15,
    63106 => -15,
    63107 => -15,
    63108 => -15,
    63109 => -15,
    63110 => -15,
    63111 => -15,
    63112 => -15,
    63113 => -15,
    63114 => -14,
    63115 => -14,
    63116 => -14,
    63117 => -14,
    63118 => -14,
    63119 => -14,
    63120 => -14,
    63121 => -14,
    63122 => -14,
    63123 => -14,
    63124 => -14,
    63125 => -14,
    63126 => -14,
    63127 => -14,
    63128 => -14,
    63129 => -14,
    63130 => -14,
    63131 => -14,
    63132 => -14,
    63133 => -14,
    63134 => -14,
    63135 => -14,
    63136 => -14,
    63137 => -14,
    63138 => -14,
    63139 => -14,
    63140 => -14,
    63141 => -14,
    63142 => -14,
    63143 => -14,
    63144 => -14,
    63145 => -14,
    63146 => -14,
    63147 => -14,
    63148 => -14,
    63149 => -14,
    63150 => -14,
    63151 => -14,
    63152 => -14,
    63153 => -14,
    63154 => -14,
    63155 => -14,
    63156 => -14,
    63157 => -14,
    63158 => -14,
    63159 => -14,
    63160 => -14,
    63161 => -14,
    63162 => -14,
    63163 => -14,
    63164 => -14,
    63165 => -14,
    63166 => -14,
    63167 => -14,
    63168 => -14,
    63169 => -14,
    63170 => -14,
    63171 => -14,
    63172 => -14,
    63173 => -14,
    63174 => -14,
    63175 => -14,
    63176 => -14,
    63177 => -14,
    63178 => -14,
    63179 => -14,
    63180 => -14,
    63181 => -14,
    63182 => -14,
    63183 => -14,
    63184 => -14,
    63185 => -14,
    63186 => -14,
    63187 => -14,
    63188 => -14,
    63189 => -14,
    63190 => -14,
    63191 => -14,
    63192 => -14,
    63193 => -14,
    63194 => -14,
    63195 => -14,
    63196 => -14,
    63197 => -14,
    63198 => -14,
    63199 => -14,
    63200 => -14,
    63201 => -14,
    63202 => -14,
    63203 => -14,
    63204 => -14,
    63205 => -14,
    63206 => -14,
    63207 => -14,
    63208 => -14,
    63209 => -14,
    63210 => -14,
    63211 => -14,
    63212 => -14,
    63213 => -14,
    63214 => -14,
    63215 => -14,
    63216 => -14,
    63217 => -14,
    63218 => -14,
    63219 => -14,
    63220 => -14,
    63221 => -14,
    63222 => -14,
    63223 => -14,
    63224 => -14,
    63225 => -14,
    63226 => -14,
    63227 => -14,
    63228 => -14,
    63229 => -14,
    63230 => -14,
    63231 => -14,
    63232 => -14,
    63233 => -14,
    63234 => -14,
    63235 => -14,
    63236 => -14,
    63237 => -14,
    63238 => -14,
    63239 => -14,
    63240 => -14,
    63241 => -14,
    63242 => -14,
    63243 => -14,
    63244 => -14,
    63245 => -14,
    63246 => -14,
    63247 => -14,
    63248 => -14,
    63249 => -14,
    63250 => -14,
    63251 => -14,
    63252 => -14,
    63253 => -14,
    63254 => -14,
    63255 => -14,
    63256 => -14,
    63257 => -14,
    63258 => -14,
    63259 => -14,
    63260 => -14,
    63261 => -14,
    63262 => -14,
    63263 => -14,
    63264 => -14,
    63265 => -14,
    63266 => -14,
    63267 => -14,
    63268 => -14,
    63269 => -14,
    63270 => -14,
    63271 => -14,
    63272 => -14,
    63273 => -14,
    63274 => -14,
    63275 => -14,
    63276 => -14,
    63277 => -14,
    63278 => -14,
    63279 => -14,
    63280 => -14,
    63281 => -14,
    63282 => -14,
    63283 => -14,
    63284 => -13,
    63285 => -13,
    63286 => -13,
    63287 => -13,
    63288 => -13,
    63289 => -13,
    63290 => -13,
    63291 => -13,
    63292 => -13,
    63293 => -13,
    63294 => -13,
    63295 => -13,
    63296 => -13,
    63297 => -13,
    63298 => -13,
    63299 => -13,
    63300 => -13,
    63301 => -13,
    63302 => -13,
    63303 => -13,
    63304 => -13,
    63305 => -13,
    63306 => -13,
    63307 => -13,
    63308 => -13,
    63309 => -13,
    63310 => -13,
    63311 => -13,
    63312 => -13,
    63313 => -13,
    63314 => -13,
    63315 => -13,
    63316 => -13,
    63317 => -13,
    63318 => -13,
    63319 => -13,
    63320 => -13,
    63321 => -13,
    63322 => -13,
    63323 => -13,
    63324 => -13,
    63325 => -13,
    63326 => -13,
    63327 => -13,
    63328 => -13,
    63329 => -13,
    63330 => -13,
    63331 => -13,
    63332 => -13,
    63333 => -13,
    63334 => -13,
    63335 => -13,
    63336 => -13,
    63337 => -13,
    63338 => -13,
    63339 => -13,
    63340 => -13,
    63341 => -13,
    63342 => -13,
    63343 => -13,
    63344 => -13,
    63345 => -13,
    63346 => -13,
    63347 => -13,
    63348 => -13,
    63349 => -13,
    63350 => -13,
    63351 => -13,
    63352 => -13,
    63353 => -13,
    63354 => -13,
    63355 => -13,
    63356 => -13,
    63357 => -13,
    63358 => -13,
    63359 => -13,
    63360 => -13,
    63361 => -13,
    63362 => -13,
    63363 => -13,
    63364 => -13,
    63365 => -13,
    63366 => -13,
    63367 => -13,
    63368 => -13,
    63369 => -13,
    63370 => -13,
    63371 => -13,
    63372 => -13,
    63373 => -13,
    63374 => -13,
    63375 => -13,
    63376 => -13,
    63377 => -13,
    63378 => -13,
    63379 => -13,
    63380 => -13,
    63381 => -13,
    63382 => -13,
    63383 => -13,
    63384 => -13,
    63385 => -13,
    63386 => -13,
    63387 => -13,
    63388 => -13,
    63389 => -13,
    63390 => -13,
    63391 => -13,
    63392 => -13,
    63393 => -13,
    63394 => -13,
    63395 => -13,
    63396 => -13,
    63397 => -13,
    63398 => -13,
    63399 => -13,
    63400 => -13,
    63401 => -13,
    63402 => -13,
    63403 => -13,
    63404 => -13,
    63405 => -13,
    63406 => -13,
    63407 => -13,
    63408 => -13,
    63409 => -13,
    63410 => -13,
    63411 => -13,
    63412 => -13,
    63413 => -13,
    63414 => -13,
    63415 => -13,
    63416 => -13,
    63417 => -13,
    63418 => -13,
    63419 => -13,
    63420 => -13,
    63421 => -13,
    63422 => -13,
    63423 => -13,
    63424 => -13,
    63425 => -13,
    63426 => -13,
    63427 => -13,
    63428 => -13,
    63429 => -13,
    63430 => -13,
    63431 => -13,
    63432 => -13,
    63433 => -13,
    63434 => -13,
    63435 => -13,
    63436 => -13,
    63437 => -13,
    63438 => -13,
    63439 => -13,
    63440 => -13,
    63441 => -13,
    63442 => -13,
    63443 => -13,
    63444 => -13,
    63445 => -13,
    63446 => -13,
    63447 => -13,
    63448 => -13,
    63449 => -13,
    63450 => -13,
    63451 => -13,
    63452 => -13,
    63453 => -12,
    63454 => -12,
    63455 => -12,
    63456 => -12,
    63457 => -12,
    63458 => -12,
    63459 => -12,
    63460 => -12,
    63461 => -12,
    63462 => -12,
    63463 => -12,
    63464 => -12,
    63465 => -12,
    63466 => -12,
    63467 => -12,
    63468 => -12,
    63469 => -12,
    63470 => -12,
    63471 => -12,
    63472 => -12,
    63473 => -12,
    63474 => -12,
    63475 => -12,
    63476 => -12,
    63477 => -12,
    63478 => -12,
    63479 => -12,
    63480 => -12,
    63481 => -12,
    63482 => -12,
    63483 => -12,
    63484 => -12,
    63485 => -12,
    63486 => -12,
    63487 => -12,
    63488 => -12,
    63489 => -12,
    63490 => -12,
    63491 => -12,
    63492 => -12,
    63493 => -12,
    63494 => -12,
    63495 => -12,
    63496 => -12,
    63497 => -12,
    63498 => -12,
    63499 => -12,
    63500 => -12,
    63501 => -12,
    63502 => -12,
    63503 => -12,
    63504 => -12,
    63505 => -12,
    63506 => -12,
    63507 => -12,
    63508 => -12,
    63509 => -12,
    63510 => -12,
    63511 => -12,
    63512 => -12,
    63513 => -12,
    63514 => -12,
    63515 => -12,
    63516 => -12,
    63517 => -12,
    63518 => -12,
    63519 => -12,
    63520 => -12,
    63521 => -12,
    63522 => -12,
    63523 => -12,
    63524 => -12,
    63525 => -12,
    63526 => -12,
    63527 => -12,
    63528 => -12,
    63529 => -12,
    63530 => -12,
    63531 => -12,
    63532 => -12,
    63533 => -12,
    63534 => -12,
    63535 => -12,
    63536 => -12,
    63537 => -12,
    63538 => -12,
    63539 => -12,
    63540 => -12,
    63541 => -12,
    63542 => -12,
    63543 => -12,
    63544 => -12,
    63545 => -12,
    63546 => -12,
    63547 => -12,
    63548 => -12,
    63549 => -12,
    63550 => -12,
    63551 => -12,
    63552 => -12,
    63553 => -12,
    63554 => -12,
    63555 => -12,
    63556 => -12,
    63557 => -12,
    63558 => -12,
    63559 => -12,
    63560 => -12,
    63561 => -12,
    63562 => -12,
    63563 => -12,
    63564 => -12,
    63565 => -12,
    63566 => -12,
    63567 => -12,
    63568 => -12,
    63569 => -12,
    63570 => -12,
    63571 => -12,
    63572 => -12,
    63573 => -12,
    63574 => -12,
    63575 => -12,
    63576 => -12,
    63577 => -12,
    63578 => -12,
    63579 => -12,
    63580 => -12,
    63581 => -12,
    63582 => -12,
    63583 => -12,
    63584 => -12,
    63585 => -12,
    63586 => -12,
    63587 => -12,
    63588 => -12,
    63589 => -12,
    63590 => -12,
    63591 => -12,
    63592 => -12,
    63593 => -12,
    63594 => -12,
    63595 => -12,
    63596 => -12,
    63597 => -12,
    63598 => -12,
    63599 => -12,
    63600 => -12,
    63601 => -12,
    63602 => -12,
    63603 => -12,
    63604 => -12,
    63605 => -12,
    63606 => -12,
    63607 => -12,
    63608 => -12,
    63609 => -12,
    63610 => -12,
    63611 => -12,
    63612 => -12,
    63613 => -12,
    63614 => -12,
    63615 => -12,
    63616 => -12,
    63617 => -12,
    63618 => -12,
    63619 => -12,
    63620 => -12,
    63621 => -12,
    63622 => -11,
    63623 => -11,
    63624 => -11,
    63625 => -11,
    63626 => -11,
    63627 => -11,
    63628 => -11,
    63629 => -11,
    63630 => -11,
    63631 => -11,
    63632 => -11,
    63633 => -11,
    63634 => -11,
    63635 => -11,
    63636 => -11,
    63637 => -11,
    63638 => -11,
    63639 => -11,
    63640 => -11,
    63641 => -11,
    63642 => -11,
    63643 => -11,
    63644 => -11,
    63645 => -11,
    63646 => -11,
    63647 => -11,
    63648 => -11,
    63649 => -11,
    63650 => -11,
    63651 => -11,
    63652 => -11,
    63653 => -11,
    63654 => -11,
    63655 => -11,
    63656 => -11,
    63657 => -11,
    63658 => -11,
    63659 => -11,
    63660 => -11,
    63661 => -11,
    63662 => -11,
    63663 => -11,
    63664 => -11,
    63665 => -11,
    63666 => -11,
    63667 => -11,
    63668 => -11,
    63669 => -11,
    63670 => -11,
    63671 => -11,
    63672 => -11,
    63673 => -11,
    63674 => -11,
    63675 => -11,
    63676 => -11,
    63677 => -11,
    63678 => -11,
    63679 => -11,
    63680 => -11,
    63681 => -11,
    63682 => -11,
    63683 => -11,
    63684 => -11,
    63685 => -11,
    63686 => -11,
    63687 => -11,
    63688 => -11,
    63689 => -11,
    63690 => -11,
    63691 => -11,
    63692 => -11,
    63693 => -11,
    63694 => -11,
    63695 => -11,
    63696 => -11,
    63697 => -11,
    63698 => -11,
    63699 => -11,
    63700 => -11,
    63701 => -11,
    63702 => -11,
    63703 => -11,
    63704 => -11,
    63705 => -11,
    63706 => -11,
    63707 => -11,
    63708 => -11,
    63709 => -11,
    63710 => -11,
    63711 => -11,
    63712 => -11,
    63713 => -11,
    63714 => -11,
    63715 => -11,
    63716 => -11,
    63717 => -11,
    63718 => -11,
    63719 => -11,
    63720 => -11,
    63721 => -11,
    63722 => -11,
    63723 => -11,
    63724 => -11,
    63725 => -11,
    63726 => -11,
    63727 => -11,
    63728 => -11,
    63729 => -11,
    63730 => -11,
    63731 => -11,
    63732 => -11,
    63733 => -11,
    63734 => -11,
    63735 => -11,
    63736 => -11,
    63737 => -11,
    63738 => -11,
    63739 => -11,
    63740 => -11,
    63741 => -11,
    63742 => -11,
    63743 => -11,
    63744 => -11,
    63745 => -11,
    63746 => -11,
    63747 => -11,
    63748 => -11,
    63749 => -11,
    63750 => -11,
    63751 => -11,
    63752 => -11,
    63753 => -11,
    63754 => -11,
    63755 => -11,
    63756 => -11,
    63757 => -11,
    63758 => -11,
    63759 => -11,
    63760 => -11,
    63761 => -11,
    63762 => -11,
    63763 => -11,
    63764 => -11,
    63765 => -11,
    63766 => -11,
    63767 => -11,
    63768 => -11,
    63769 => -11,
    63770 => -11,
    63771 => -11,
    63772 => -11,
    63773 => -11,
    63774 => -11,
    63775 => -11,
    63776 => -11,
    63777 => -11,
    63778 => -11,
    63779 => -11,
    63780 => -11,
    63781 => -11,
    63782 => -11,
    63783 => -11,
    63784 => -11,
    63785 => -11,
    63786 => -11,
    63787 => -11,
    63788 => -11,
    63789 => -11,
    63790 => -10,
    63791 => -10,
    63792 => -10,
    63793 => -10,
    63794 => -10,
    63795 => -10,
    63796 => -10,
    63797 => -10,
    63798 => -10,
    63799 => -10,
    63800 => -10,
    63801 => -10,
    63802 => -10,
    63803 => -10,
    63804 => -10,
    63805 => -10,
    63806 => -10,
    63807 => -10,
    63808 => -10,
    63809 => -10,
    63810 => -10,
    63811 => -10,
    63812 => -10,
    63813 => -10,
    63814 => -10,
    63815 => -10,
    63816 => -10,
    63817 => -10,
    63818 => -10,
    63819 => -10,
    63820 => -10,
    63821 => -10,
    63822 => -10,
    63823 => -10,
    63824 => -10,
    63825 => -10,
    63826 => -10,
    63827 => -10,
    63828 => -10,
    63829 => -10,
    63830 => -10,
    63831 => -10,
    63832 => -10,
    63833 => -10,
    63834 => -10,
    63835 => -10,
    63836 => -10,
    63837 => -10,
    63838 => -10,
    63839 => -10,
    63840 => -10,
    63841 => -10,
    63842 => -10,
    63843 => -10,
    63844 => -10,
    63845 => -10,
    63846 => -10,
    63847 => -10,
    63848 => -10,
    63849 => -10,
    63850 => -10,
    63851 => -10,
    63852 => -10,
    63853 => -10,
    63854 => -10,
    63855 => -10,
    63856 => -10,
    63857 => -10,
    63858 => -10,
    63859 => -10,
    63860 => -10,
    63861 => -10,
    63862 => -10,
    63863 => -10,
    63864 => -10,
    63865 => -10,
    63866 => -10,
    63867 => -10,
    63868 => -10,
    63869 => -10,
    63870 => -10,
    63871 => -10,
    63872 => -10,
    63873 => -10,
    63874 => -10,
    63875 => -10,
    63876 => -10,
    63877 => -10,
    63878 => -10,
    63879 => -10,
    63880 => -10,
    63881 => -10,
    63882 => -10,
    63883 => -10,
    63884 => -10,
    63885 => -10,
    63886 => -10,
    63887 => -10,
    63888 => -10,
    63889 => -10,
    63890 => -10,
    63891 => -10,
    63892 => -10,
    63893 => -10,
    63894 => -10,
    63895 => -10,
    63896 => -10,
    63897 => -10,
    63898 => -10,
    63899 => -10,
    63900 => -10,
    63901 => -10,
    63902 => -10,
    63903 => -10,
    63904 => -10,
    63905 => -10,
    63906 => -10,
    63907 => -10,
    63908 => -10,
    63909 => -10,
    63910 => -10,
    63911 => -10,
    63912 => -10,
    63913 => -10,
    63914 => -10,
    63915 => -10,
    63916 => -10,
    63917 => -10,
    63918 => -10,
    63919 => -10,
    63920 => -10,
    63921 => -10,
    63922 => -10,
    63923 => -10,
    63924 => -10,
    63925 => -10,
    63926 => -10,
    63927 => -10,
    63928 => -10,
    63929 => -10,
    63930 => -10,
    63931 => -10,
    63932 => -10,
    63933 => -10,
    63934 => -10,
    63935 => -10,
    63936 => -10,
    63937 => -10,
    63938 => -10,
    63939 => -10,
    63940 => -10,
    63941 => -10,
    63942 => -10,
    63943 => -10,
    63944 => -10,
    63945 => -10,
    63946 => -10,
    63947 => -10,
    63948 => -10,
    63949 => -10,
    63950 => -10,
    63951 => -10,
    63952 => -10,
    63953 => -10,
    63954 => -10,
    63955 => -10,
    63956 => -10,
    63957 => -10,
    63958 => -9,
    63959 => -9,
    63960 => -9,
    63961 => -9,
    63962 => -9,
    63963 => -9,
    63964 => -9,
    63965 => -9,
    63966 => -9,
    63967 => -9,
    63968 => -9,
    63969 => -9,
    63970 => -9,
    63971 => -9,
    63972 => -9,
    63973 => -9,
    63974 => -9,
    63975 => -9,
    63976 => -9,
    63977 => -9,
    63978 => -9,
    63979 => -9,
    63980 => -9,
    63981 => -9,
    63982 => -9,
    63983 => -9,
    63984 => -9,
    63985 => -9,
    63986 => -9,
    63987 => -9,
    63988 => -9,
    63989 => -9,
    63990 => -9,
    63991 => -9,
    63992 => -9,
    63993 => -9,
    63994 => -9,
    63995 => -9,
    63996 => -9,
    63997 => -9,
    63998 => -9,
    63999 => -9,
    64000 => -9,
    64001 => -9,
    64002 => -9,
    64003 => -9,
    64004 => -9,
    64005 => -9,
    64006 => -9,
    64007 => -9,
    64008 => -9,
    64009 => -9,
    64010 => -9,
    64011 => -9,
    64012 => -9,
    64013 => -9,
    64014 => -9,
    64015 => -9,
    64016 => -9,
    64017 => -9,
    64018 => -9,
    64019 => -9,
    64020 => -9,
    64021 => -9,
    64022 => -9,
    64023 => -9,
    64024 => -9,
    64025 => -9,
    64026 => -9,
    64027 => -9,
    64028 => -9,
    64029 => -9,
    64030 => -9,
    64031 => -9,
    64032 => -9,
    64033 => -9,
    64034 => -9,
    64035 => -9,
    64036 => -9,
    64037 => -9,
    64038 => -9,
    64039 => -9,
    64040 => -9,
    64041 => -9,
    64042 => -9,
    64043 => -9,
    64044 => -9,
    64045 => -9,
    64046 => -9,
    64047 => -9,
    64048 => -9,
    64049 => -9,
    64050 => -9,
    64051 => -9,
    64052 => -9,
    64053 => -9,
    64054 => -9,
    64055 => -9,
    64056 => -9,
    64057 => -9,
    64058 => -9,
    64059 => -9,
    64060 => -9,
    64061 => -9,
    64062 => -9,
    64063 => -9,
    64064 => -9,
    64065 => -9,
    64066 => -9,
    64067 => -9,
    64068 => -9,
    64069 => -9,
    64070 => -9,
    64071 => -9,
    64072 => -9,
    64073 => -9,
    64074 => -9,
    64075 => -9,
    64076 => -9,
    64077 => -9,
    64078 => -9,
    64079 => -9,
    64080 => -9,
    64081 => -9,
    64082 => -9,
    64083 => -9,
    64084 => -9,
    64085 => -9,
    64086 => -9,
    64087 => -9,
    64088 => -9,
    64089 => -9,
    64090 => -9,
    64091 => -9,
    64092 => -9,
    64093 => -9,
    64094 => -9,
    64095 => -9,
    64096 => -9,
    64097 => -9,
    64098 => -9,
    64099 => -9,
    64100 => -9,
    64101 => -9,
    64102 => -9,
    64103 => -9,
    64104 => -9,
    64105 => -9,
    64106 => -9,
    64107 => -9,
    64108 => -9,
    64109 => -9,
    64110 => -9,
    64111 => -9,
    64112 => -9,
    64113 => -9,
    64114 => -9,
    64115 => -9,
    64116 => -9,
    64117 => -9,
    64118 => -9,
    64119 => -9,
    64120 => -9,
    64121 => -9,
    64122 => -9,
    64123 => -9,
    64124 => -9,
    64125 => -8,
    64126 => -8,
    64127 => -8,
    64128 => -8,
    64129 => -8,
    64130 => -8,
    64131 => -8,
    64132 => -8,
    64133 => -8,
    64134 => -8,
    64135 => -8,
    64136 => -8,
    64137 => -8,
    64138 => -8,
    64139 => -8,
    64140 => -8,
    64141 => -8,
    64142 => -8,
    64143 => -8,
    64144 => -8,
    64145 => -8,
    64146 => -8,
    64147 => -8,
    64148 => -8,
    64149 => -8,
    64150 => -8,
    64151 => -8,
    64152 => -8,
    64153 => -8,
    64154 => -8,
    64155 => -8,
    64156 => -8,
    64157 => -8,
    64158 => -8,
    64159 => -8,
    64160 => -8,
    64161 => -8,
    64162 => -8,
    64163 => -8,
    64164 => -8,
    64165 => -8,
    64166 => -8,
    64167 => -8,
    64168 => -8,
    64169 => -8,
    64170 => -8,
    64171 => -8,
    64172 => -8,
    64173 => -8,
    64174 => -8,
    64175 => -8,
    64176 => -8,
    64177 => -8,
    64178 => -8,
    64179 => -8,
    64180 => -8,
    64181 => -8,
    64182 => -8,
    64183 => -8,
    64184 => -8,
    64185 => -8,
    64186 => -8,
    64187 => -8,
    64188 => -8,
    64189 => -8,
    64190 => -8,
    64191 => -8,
    64192 => -8,
    64193 => -8,
    64194 => -8,
    64195 => -8,
    64196 => -8,
    64197 => -8,
    64198 => -8,
    64199 => -8,
    64200 => -8,
    64201 => -8,
    64202 => -8,
    64203 => -8,
    64204 => -8,
    64205 => -8,
    64206 => -8,
    64207 => -8,
    64208 => -8,
    64209 => -8,
    64210 => -8,
    64211 => -8,
    64212 => -8,
    64213 => -8,
    64214 => -8,
    64215 => -8,
    64216 => -8,
    64217 => -8,
    64218 => -8,
    64219 => -8,
    64220 => -8,
    64221 => -8,
    64222 => -8,
    64223 => -8,
    64224 => -8,
    64225 => -8,
    64226 => -8,
    64227 => -8,
    64228 => -8,
    64229 => -8,
    64230 => -8,
    64231 => -8,
    64232 => -8,
    64233 => -8,
    64234 => -8,
    64235 => -8,
    64236 => -8,
    64237 => -8,
    64238 => -8,
    64239 => -8,
    64240 => -8,
    64241 => -8,
    64242 => -8,
    64243 => -8,
    64244 => -8,
    64245 => -8,
    64246 => -8,
    64247 => -8,
    64248 => -8,
    64249 => -8,
    64250 => -8,
    64251 => -8,
    64252 => -8,
    64253 => -8,
    64254 => -8,
    64255 => -8,
    64256 => -8,
    64257 => -8,
    64258 => -8,
    64259 => -8,
    64260 => -8,
    64261 => -8,
    64262 => -8,
    64263 => -8,
    64264 => -8,
    64265 => -8,
    64266 => -8,
    64267 => -8,
    64268 => -8,
    64269 => -8,
    64270 => -8,
    64271 => -8,
    64272 => -8,
    64273 => -8,
    64274 => -8,
    64275 => -8,
    64276 => -8,
    64277 => -8,
    64278 => -8,
    64279 => -8,
    64280 => -8,
    64281 => -8,
    64282 => -8,
    64283 => -8,
    64284 => -8,
    64285 => -8,
    64286 => -8,
    64287 => -8,
    64288 => -8,
    64289 => -8,
    64290 => -8,
    64291 => -8,
    64292 => -7,
    64293 => -7,
    64294 => -7,
    64295 => -7,
    64296 => -7,
    64297 => -7,
    64298 => -7,
    64299 => -7,
    64300 => -7,
    64301 => -7,
    64302 => -7,
    64303 => -7,
    64304 => -7,
    64305 => -7,
    64306 => -7,
    64307 => -7,
    64308 => -7,
    64309 => -7,
    64310 => -7,
    64311 => -7,
    64312 => -7,
    64313 => -7,
    64314 => -7,
    64315 => -7,
    64316 => -7,
    64317 => -7,
    64318 => -7,
    64319 => -7,
    64320 => -7,
    64321 => -7,
    64322 => -7,
    64323 => -7,
    64324 => -7,
    64325 => -7,
    64326 => -7,
    64327 => -7,
    64328 => -7,
    64329 => -7,
    64330 => -7,
    64331 => -7,
    64332 => -7,
    64333 => -7,
    64334 => -7,
    64335 => -7,
    64336 => -7,
    64337 => -7,
    64338 => -7,
    64339 => -7,
    64340 => -7,
    64341 => -7,
    64342 => -7,
    64343 => -7,
    64344 => -7,
    64345 => -7,
    64346 => -7,
    64347 => -7,
    64348 => -7,
    64349 => -7,
    64350 => -7,
    64351 => -7,
    64352 => -7,
    64353 => -7,
    64354 => -7,
    64355 => -7,
    64356 => -7,
    64357 => -7,
    64358 => -7,
    64359 => -7,
    64360 => -7,
    64361 => -7,
    64362 => -7,
    64363 => -7,
    64364 => -7,
    64365 => -7,
    64366 => -7,
    64367 => -7,
    64368 => -7,
    64369 => -7,
    64370 => -7,
    64371 => -7,
    64372 => -7,
    64373 => -7,
    64374 => -7,
    64375 => -7,
    64376 => -7,
    64377 => -7,
    64378 => -7,
    64379 => -7,
    64380 => -7,
    64381 => -7,
    64382 => -7,
    64383 => -7,
    64384 => -7,
    64385 => -7,
    64386 => -7,
    64387 => -7,
    64388 => -7,
    64389 => -7,
    64390 => -7,
    64391 => -7,
    64392 => -7,
    64393 => -7,
    64394 => -7,
    64395 => -7,
    64396 => -7,
    64397 => -7,
    64398 => -7,
    64399 => -7,
    64400 => -7,
    64401 => -7,
    64402 => -7,
    64403 => -7,
    64404 => -7,
    64405 => -7,
    64406 => -7,
    64407 => -7,
    64408 => -7,
    64409 => -7,
    64410 => -7,
    64411 => -7,
    64412 => -7,
    64413 => -7,
    64414 => -7,
    64415 => -7,
    64416 => -7,
    64417 => -7,
    64418 => -7,
    64419 => -7,
    64420 => -7,
    64421 => -7,
    64422 => -7,
    64423 => -7,
    64424 => -7,
    64425 => -7,
    64426 => -7,
    64427 => -7,
    64428 => -7,
    64429 => -7,
    64430 => -7,
    64431 => -7,
    64432 => -7,
    64433 => -7,
    64434 => -7,
    64435 => -7,
    64436 => -7,
    64437 => -7,
    64438 => -7,
    64439 => -7,
    64440 => -7,
    64441 => -7,
    64442 => -7,
    64443 => -7,
    64444 => -7,
    64445 => -7,
    64446 => -7,
    64447 => -7,
    64448 => -7,
    64449 => -7,
    64450 => -7,
    64451 => -7,
    64452 => -7,
    64453 => -7,
    64454 => -7,
    64455 => -7,
    64456 => -7,
    64457 => -7,
    64458 => -6,
    64459 => -6,
    64460 => -6,
    64461 => -6,
    64462 => -6,
    64463 => -6,
    64464 => -6,
    64465 => -6,
    64466 => -6,
    64467 => -6,
    64468 => -6,
    64469 => -6,
    64470 => -6,
    64471 => -6,
    64472 => -6,
    64473 => -6,
    64474 => -6,
    64475 => -6,
    64476 => -6,
    64477 => -6,
    64478 => -6,
    64479 => -6,
    64480 => -6,
    64481 => -6,
    64482 => -6,
    64483 => -6,
    64484 => -6,
    64485 => -6,
    64486 => -6,
    64487 => -6,
    64488 => -6,
    64489 => -6,
    64490 => -6,
    64491 => -6,
    64492 => -6,
    64493 => -6,
    64494 => -6,
    64495 => -6,
    64496 => -6,
    64497 => -6,
    64498 => -6,
    64499 => -6,
    64500 => -6,
    64501 => -6,
    64502 => -6,
    64503 => -6,
    64504 => -6,
    64505 => -6,
    64506 => -6,
    64507 => -6,
    64508 => -6,
    64509 => -6,
    64510 => -6,
    64511 => -6,
    64512 => -6,
    64513 => -6,
    64514 => -6,
    64515 => -6,
    64516 => -6,
    64517 => -6,
    64518 => -6,
    64519 => -6,
    64520 => -6,
    64521 => -6,
    64522 => -6,
    64523 => -6,
    64524 => -6,
    64525 => -6,
    64526 => -6,
    64527 => -6,
    64528 => -6,
    64529 => -6,
    64530 => -6,
    64531 => -6,
    64532 => -6,
    64533 => -6,
    64534 => -6,
    64535 => -6,
    64536 => -6,
    64537 => -6,
    64538 => -6,
    64539 => -6,
    64540 => -6,
    64541 => -6,
    64542 => -6,
    64543 => -6,
    64544 => -6,
    64545 => -6,
    64546 => -6,
    64547 => -6,
    64548 => -6,
    64549 => -6,
    64550 => -6,
    64551 => -6,
    64552 => -6,
    64553 => -6,
    64554 => -6,
    64555 => -6,
    64556 => -6,
    64557 => -6,
    64558 => -6,
    64559 => -6,
    64560 => -6,
    64561 => -6,
    64562 => -6,
    64563 => -6,
    64564 => -6,
    64565 => -6,
    64566 => -6,
    64567 => -6,
    64568 => -6,
    64569 => -6,
    64570 => -6,
    64571 => -6,
    64572 => -6,
    64573 => -6,
    64574 => -6,
    64575 => -6,
    64576 => -6,
    64577 => -6,
    64578 => -6,
    64579 => -6,
    64580 => -6,
    64581 => -6,
    64582 => -6,
    64583 => -6,
    64584 => -6,
    64585 => -6,
    64586 => -6,
    64587 => -6,
    64588 => -6,
    64589 => -6,
    64590 => -6,
    64591 => -6,
    64592 => -6,
    64593 => -6,
    64594 => -6,
    64595 => -6,
    64596 => -6,
    64597 => -6,
    64598 => -6,
    64599 => -6,
    64600 => -6,
    64601 => -6,
    64602 => -6,
    64603 => -6,
    64604 => -6,
    64605 => -6,
    64606 => -6,
    64607 => -6,
    64608 => -6,
    64609 => -6,
    64610 => -6,
    64611 => -6,
    64612 => -6,
    64613 => -6,
    64614 => -6,
    64615 => -6,
    64616 => -6,
    64617 => -6,
    64618 => -6,
    64619 => -6,
    64620 => -6,
    64621 => -6,
    64622 => -6,
    64623 => -6,
    64624 => -6,
    64625 => -5,
    64626 => -5,
    64627 => -5,
    64628 => -5,
    64629 => -5,
    64630 => -5,
    64631 => -5,
    64632 => -5,
    64633 => -5,
    64634 => -5,
    64635 => -5,
    64636 => -5,
    64637 => -5,
    64638 => -5,
    64639 => -5,
    64640 => -5,
    64641 => -5,
    64642 => -5,
    64643 => -5,
    64644 => -5,
    64645 => -5,
    64646 => -5,
    64647 => -5,
    64648 => -5,
    64649 => -5,
    64650 => -5,
    64651 => -5,
    64652 => -5,
    64653 => -5,
    64654 => -5,
    64655 => -5,
    64656 => -5,
    64657 => -5,
    64658 => -5,
    64659 => -5,
    64660 => -5,
    64661 => -5,
    64662 => -5,
    64663 => -5,
    64664 => -5,
    64665 => -5,
    64666 => -5,
    64667 => -5,
    64668 => -5,
    64669 => -5,
    64670 => -5,
    64671 => -5,
    64672 => -5,
    64673 => -5,
    64674 => -5,
    64675 => -5,
    64676 => -5,
    64677 => -5,
    64678 => -5,
    64679 => -5,
    64680 => -5,
    64681 => -5,
    64682 => -5,
    64683 => -5,
    64684 => -5,
    64685 => -5,
    64686 => -5,
    64687 => -5,
    64688 => -5,
    64689 => -5,
    64690 => -5,
    64691 => -5,
    64692 => -5,
    64693 => -5,
    64694 => -5,
    64695 => -5,
    64696 => -5,
    64697 => -5,
    64698 => -5,
    64699 => -5,
    64700 => -5,
    64701 => -5,
    64702 => -5,
    64703 => -5,
    64704 => -5,
    64705 => -5,
    64706 => -5,
    64707 => -5,
    64708 => -5,
    64709 => -5,
    64710 => -5,
    64711 => -5,
    64712 => -5,
    64713 => -5,
    64714 => -5,
    64715 => -5,
    64716 => -5,
    64717 => -5,
    64718 => -5,
    64719 => -5,
    64720 => -5,
    64721 => -5,
    64722 => -5,
    64723 => -5,
    64724 => -5,
    64725 => -5,
    64726 => -5,
    64727 => -5,
    64728 => -5,
    64729 => -5,
    64730 => -5,
    64731 => -5,
    64732 => -5,
    64733 => -5,
    64734 => -5,
    64735 => -5,
    64736 => -5,
    64737 => -5,
    64738 => -5,
    64739 => -5,
    64740 => -5,
    64741 => -5,
    64742 => -5,
    64743 => -5,
    64744 => -5,
    64745 => -5,
    64746 => -5,
    64747 => -5,
    64748 => -5,
    64749 => -5,
    64750 => -5,
    64751 => -5,
    64752 => -5,
    64753 => -5,
    64754 => -5,
    64755 => -5,
    64756 => -5,
    64757 => -5,
    64758 => -5,
    64759 => -5,
    64760 => -5,
    64761 => -5,
    64762 => -5,
    64763 => -5,
    64764 => -5,
    64765 => -5,
    64766 => -5,
    64767 => -5,
    64768 => -5,
    64769 => -5,
    64770 => -5,
    64771 => -5,
    64772 => -5,
    64773 => -5,
    64774 => -5,
    64775 => -5,
    64776 => -5,
    64777 => -5,
    64778 => -5,
    64779 => -5,
    64780 => -5,
    64781 => -5,
    64782 => -5,
    64783 => -5,
    64784 => -5,
    64785 => -5,
    64786 => -5,
    64787 => -5,
    64788 => -5,
    64789 => -5,
    64790 => -5,
    64791 => -4,
    64792 => -4,
    64793 => -4,
    64794 => -4,
    64795 => -4,
    64796 => -4,
    64797 => -4,
    64798 => -4,
    64799 => -4,
    64800 => -4,
    64801 => -4,
    64802 => -4,
    64803 => -4,
    64804 => -4,
    64805 => -4,
    64806 => -4,
    64807 => -4,
    64808 => -4,
    64809 => -4,
    64810 => -4,
    64811 => -4,
    64812 => -4,
    64813 => -4,
    64814 => -4,
    64815 => -4,
    64816 => -4,
    64817 => -4,
    64818 => -4,
    64819 => -4,
    64820 => -4,
    64821 => -4,
    64822 => -4,
    64823 => -4,
    64824 => -4,
    64825 => -4,
    64826 => -4,
    64827 => -4,
    64828 => -4,
    64829 => -4,
    64830 => -4,
    64831 => -4,
    64832 => -4,
    64833 => -4,
    64834 => -4,
    64835 => -4,
    64836 => -4,
    64837 => -4,
    64838 => -4,
    64839 => -4,
    64840 => -4,
    64841 => -4,
    64842 => -4,
    64843 => -4,
    64844 => -4,
    64845 => -4,
    64846 => -4,
    64847 => -4,
    64848 => -4,
    64849 => -4,
    64850 => -4,
    64851 => -4,
    64852 => -4,
    64853 => -4,
    64854 => -4,
    64855 => -4,
    64856 => -4,
    64857 => -4,
    64858 => -4,
    64859 => -4,
    64860 => -4,
    64861 => -4,
    64862 => -4,
    64863 => -4,
    64864 => -4,
    64865 => -4,
    64866 => -4,
    64867 => -4,
    64868 => -4,
    64869 => -4,
    64870 => -4,
    64871 => -4,
    64872 => -4,
    64873 => -4,
    64874 => -4,
    64875 => -4,
    64876 => -4,
    64877 => -4,
    64878 => -4,
    64879 => -4,
    64880 => -4,
    64881 => -4,
    64882 => -4,
    64883 => -4,
    64884 => -4,
    64885 => -4,
    64886 => -4,
    64887 => -4,
    64888 => -4,
    64889 => -4,
    64890 => -4,
    64891 => -4,
    64892 => -4,
    64893 => -4,
    64894 => -4,
    64895 => -4,
    64896 => -4,
    64897 => -4,
    64898 => -4,
    64899 => -4,
    64900 => -4,
    64901 => -4,
    64902 => -4,
    64903 => -4,
    64904 => -4,
    64905 => -4,
    64906 => -4,
    64907 => -4,
    64908 => -4,
    64909 => -4,
    64910 => -4,
    64911 => -4,
    64912 => -4,
    64913 => -4,
    64914 => -4,
    64915 => -4,
    64916 => -4,
    64917 => -4,
    64918 => -4,
    64919 => -4,
    64920 => -4,
    64921 => -4,
    64922 => -4,
    64923 => -4,
    64924 => -4,
    64925 => -4,
    64926 => -4,
    64927 => -4,
    64928 => -4,
    64929 => -4,
    64930 => -4,
    64931 => -4,
    64932 => -4,
    64933 => -4,
    64934 => -4,
    64935 => -4,
    64936 => -4,
    64937 => -4,
    64938 => -4,
    64939 => -4,
    64940 => -4,
    64941 => -4,
    64942 => -4,
    64943 => -4,
    64944 => -4,
    64945 => -4,
    64946 => -4,
    64947 => -4,
    64948 => -4,
    64949 => -4,
    64950 => -4,
    64951 => -4,
    64952 => -4,
    64953 => -4,
    64954 => -4,
    64955 => -4,
    64956 => -4,
    64957 => -3,
    64958 => -3,
    64959 => -3,
    64960 => -3,
    64961 => -3,
    64962 => -3,
    64963 => -3,
    64964 => -3,
    64965 => -3,
    64966 => -3,
    64967 => -3,
    64968 => -3,
    64969 => -3,
    64970 => -3,
    64971 => -3,
    64972 => -3,
    64973 => -3,
    64974 => -3,
    64975 => -3,
    64976 => -3,
    64977 => -3,
    64978 => -3,
    64979 => -3,
    64980 => -3,
    64981 => -3,
    64982 => -3,
    64983 => -3,
    64984 => -3,
    64985 => -3,
    64986 => -3,
    64987 => -3,
    64988 => -3,
    64989 => -3,
    64990 => -3,
    64991 => -3,
    64992 => -3,
    64993 => -3,
    64994 => -3,
    64995 => -3,
    64996 => -3,
    64997 => -3,
    64998 => -3,
    64999 => -3,
    65000 => -3,
    65001 => -3,
    65002 => -3,
    65003 => -3,
    65004 => -3,
    65005 => -3,
    65006 => -3,
    65007 => -3,
    65008 => -3,
    65009 => -3,
    65010 => -3,
    65011 => -3,
    65012 => -3,
    65013 => -3,
    65014 => -3,
    65015 => -3,
    65016 => -3,
    65017 => -3,
    65018 => -3,
    65019 => -3,
    65020 => -3,
    65021 => -3,
    65022 => -3,
    65023 => -3,
    65024 => -3,
    65025 => -3,
    65026 => -3,
    65027 => -3,
    65028 => -3,
    65029 => -3,
    65030 => -3,
    65031 => -3,
    65032 => -3,
    65033 => -3,
    65034 => -3,
    65035 => -3,
    65036 => -3,
    65037 => -3,
    65038 => -3,
    65039 => -3,
    65040 => -3,
    65041 => -3,
    65042 => -3,
    65043 => -3,
    65044 => -3,
    65045 => -3,
    65046 => -3,
    65047 => -3,
    65048 => -3,
    65049 => -3,
    65050 => -3,
    65051 => -3,
    65052 => -3,
    65053 => -3,
    65054 => -3,
    65055 => -3,
    65056 => -3,
    65057 => -3,
    65058 => -3,
    65059 => -3,
    65060 => -3,
    65061 => -3,
    65062 => -3,
    65063 => -3,
    65064 => -3,
    65065 => -3,
    65066 => -3,
    65067 => -3,
    65068 => -3,
    65069 => -3,
    65070 => -3,
    65071 => -3,
    65072 => -3,
    65073 => -3,
    65074 => -3,
    65075 => -3,
    65076 => -3,
    65077 => -3,
    65078 => -3,
    65079 => -3,
    65080 => -3,
    65081 => -3,
    65082 => -3,
    65083 => -3,
    65084 => -3,
    65085 => -3,
    65086 => -3,
    65087 => -3,
    65088 => -3,
    65089 => -3,
    65090 => -3,
    65091 => -3,
    65092 => -3,
    65093 => -3,
    65094 => -3,
    65095 => -3,
    65096 => -3,
    65097 => -3,
    65098 => -3,
    65099 => -3,
    65100 => -3,
    65101 => -3,
    65102 => -3,
    65103 => -3,
    65104 => -3,
    65105 => -3,
    65106 => -3,
    65107 => -3,
    65108 => -3,
    65109 => -3,
    65110 => -3,
    65111 => -3,
    65112 => -3,
    65113 => -3,
    65114 => -3,
    65115 => -3,
    65116 => -3,
    65117 => -3,
    65118 => -3,
    65119 => -3,
    65120 => -3,
    65121 => -3,
    65122 => -2,
    65123 => -2,
    65124 => -2,
    65125 => -2,
    65126 => -2,
    65127 => -2,
    65128 => -2,
    65129 => -2,
    65130 => -2,
    65131 => -2,
    65132 => -2,
    65133 => -2,
    65134 => -2,
    65135 => -2,
    65136 => -2,
    65137 => -2,
    65138 => -2,
    65139 => -2,
    65140 => -2,
    65141 => -2,
    65142 => -2,
    65143 => -2,
    65144 => -2,
    65145 => -2,
    65146 => -2,
    65147 => -2,
    65148 => -2,
    65149 => -2,
    65150 => -2,
    65151 => -2,
    65152 => -2,
    65153 => -2,
    65154 => -2,
    65155 => -2,
    65156 => -2,
    65157 => -2,
    65158 => -2,
    65159 => -2,
    65160 => -2,
    65161 => -2,
    65162 => -2,
    65163 => -2,
    65164 => -2,
    65165 => -2,
    65166 => -2,
    65167 => -2,
    65168 => -2,
    65169 => -2,
    65170 => -2,
    65171 => -2,
    65172 => -2,
    65173 => -2,
    65174 => -2,
    65175 => -2,
    65176 => -2,
    65177 => -2,
    65178 => -2,
    65179 => -2,
    65180 => -2,
    65181 => -2,
    65182 => -2,
    65183 => -2,
    65184 => -2,
    65185 => -2,
    65186 => -2,
    65187 => -2,
    65188 => -2,
    65189 => -2,
    65190 => -2,
    65191 => -2,
    65192 => -2,
    65193 => -2,
    65194 => -2,
    65195 => -2,
    65196 => -2,
    65197 => -2,
    65198 => -2,
    65199 => -2,
    65200 => -2,
    65201 => -2,
    65202 => -2,
    65203 => -2,
    65204 => -2,
    65205 => -2,
    65206 => -2,
    65207 => -2,
    65208 => -2,
    65209 => -2,
    65210 => -2,
    65211 => -2,
    65212 => -2,
    65213 => -2,
    65214 => -2,
    65215 => -2,
    65216 => -2,
    65217 => -2,
    65218 => -2,
    65219 => -2,
    65220 => -2,
    65221 => -2,
    65222 => -2,
    65223 => -2,
    65224 => -2,
    65225 => -2,
    65226 => -2,
    65227 => -2,
    65228 => -2,
    65229 => -2,
    65230 => -2,
    65231 => -2,
    65232 => -2,
    65233 => -2,
    65234 => -2,
    65235 => -2,
    65236 => -2,
    65237 => -2,
    65238 => -2,
    65239 => -2,
    65240 => -2,
    65241 => -2,
    65242 => -2,
    65243 => -2,
    65244 => -2,
    65245 => -2,
    65246 => -2,
    65247 => -2,
    65248 => -2,
    65249 => -2,
    65250 => -2,
    65251 => -2,
    65252 => -2,
    65253 => -2,
    65254 => -2,
    65255 => -2,
    65256 => -2,
    65257 => -2,
    65258 => -2,
    65259 => -2,
    65260 => -2,
    65261 => -2,
    65262 => -2,
    65263 => -2,
    65264 => -2,
    65265 => -2,
    65266 => -2,
    65267 => -2,
    65268 => -2,
    65269 => -2,
    65270 => -2,
    65271 => -2,
    65272 => -2,
    65273 => -2,
    65274 => -2,
    65275 => -2,
    65276 => -2,
    65277 => -2,
    65278 => -2,
    65279 => -2,
    65280 => -2,
    65281 => -2,
    65282 => -2,
    65283 => -2,
    65284 => -2,
    65285 => -2,
    65286 => -2,
    65287 => -2,
    65288 => -1,
    65289 => -1,
    65290 => -1,
    65291 => -1,
    65292 => -1,
    65293 => -1,
    65294 => -1,
    65295 => -1,
    65296 => -1,
    65297 => -1,
    65298 => -1,
    65299 => -1,
    65300 => -1,
    65301 => -1,
    65302 => -1,
    65303 => -1,
    65304 => -1,
    65305 => -1,
    65306 => -1,
    65307 => -1,
    65308 => -1,
    65309 => -1,
    65310 => -1,
    65311 => -1,
    65312 => -1,
    65313 => -1,
    65314 => -1,
    65315 => -1,
    65316 => -1,
    65317 => -1,
    65318 => -1,
    65319 => -1,
    65320 => -1,
    65321 => -1,
    65322 => -1,
    65323 => -1,
    65324 => -1,
    65325 => -1,
    65326 => -1,
    65327 => -1,
    65328 => -1,
    65329 => -1,
    65330 => -1,
    65331 => -1,
    65332 => -1,
    65333 => -1,
    65334 => -1,
    65335 => -1,
    65336 => -1,
    65337 => -1,
    65338 => -1,
    65339 => -1,
    65340 => -1,
    65341 => -1,
    65342 => -1,
    65343 => -1,
    65344 => -1,
    65345 => -1,
    65346 => -1,
    65347 => -1,
    65348 => -1,
    65349 => -1,
    65350 => -1,
    65351 => -1,
    65352 => -1,
    65353 => -1,
    65354 => -1,
    65355 => -1,
    65356 => -1,
    65357 => -1,
    65358 => -1,
    65359 => -1,
    65360 => -1,
    65361 => -1,
    65362 => -1,
    65363 => -1,
    65364 => -1,
    65365 => -1,
    65366 => -1,
    65367 => -1,
    65368 => -1,
    65369 => -1,
    65370 => -1,
    65371 => -1,
    65372 => -1,
    65373 => -1,
    65374 => -1,
    65375 => -1,
    65376 => -1,
    65377 => -1,
    65378 => -1,
    65379 => -1,
    65380 => -1,
    65381 => -1,
    65382 => -1,
    65383 => -1,
    65384 => -1,
    65385 => -1,
    65386 => -1,
    65387 => -1,
    65388 => -1,
    65389 => -1,
    65390 => -1,
    65391 => -1,
    65392 => -1,
    65393 => -1,
    65394 => -1,
    65395 => -1,
    65396 => -1,
    65397 => -1,
    65398 => -1,
    65399 => -1,
    65400 => -1,
    65401 => -1,
    65402 => -1,
    65403 => -1,
    65404 => -1,
    65405 => -1,
    65406 => -1,
    65407 => -1,
    65408 => -1,
    65409 => -1,
    65410 => -1,
    65411 => -1,
    65412 => -1,
    65413 => -1,
    65414 => -1,
    65415 => -1,
    65416 => -1,
    65417 => -1,
    65418 => -1,
    65419 => -1,
    65420 => -1,
    65421 => -1,
    65422 => -1,
    65423 => -1,
    65424 => -1,
    65425 => -1,
    65426 => -1,
    65427 => -1,
    65428 => -1,
    65429 => -1,
    65430 => -1,
    65431 => -1,
    65432 => -1,
    65433 => -1,
    65434 => -1,
    65435 => -1,
    65436 => -1,
    65437 => -1,
    65438 => -1,
    65439 => -1,
    65440 => -1,
    65441 => -1,
    65442 => -1,
    65443 => -1,
    65444 => -1,
    65445 => -1,
    65446 => -1,
    65447 => -1,
    65448 => -1,
    65449 => -1,
    65450 => -1,
    65451 => -1,
    65452 => -1,
    65453 => -1,
    65454 => 0,
    65455 => 0,
    65456 => 0,
    65457 => 0,
    65458 => 0,
    65459 => 0,
    65460 => 0,
    65461 => 0,
    65462 => 0,
    65463 => 0,
    65464 => 0,
    65465 => 0,
    65466 => 0,
    65467 => 0,
    65468 => 0,
    65469 => 0,
    65470 => 0,
    65471 => 0,
    65472 => 0,
    65473 => 0,
    65474 => 0,
    65475 => 0,
    65476 => 0,
    65477 => 0,
    65478 => 0,
    65479 => 0,
    65480 => 0,
    65481 => 0,
    65482 => 0,
    65483 => 0,
    65484 => 0,
    65485 => 0,
    65486 => 0,
    65487 => 0,
    65488 => 0,
    65489 => 0,
    65490 => 0,
    65491 => 0,
    65492 => 0,
    65493 => 0,
    65494 => 0,
    65495 => 0,
    65496 => 0,
    65497 => 0,
    65498 => 0,
    65499 => 0,
    65500 => 0,
    65501 => 0,
    65502 => 0,
    65503 => 0,
    65504 => 0,
    65505 => 0,
    65506 => 0,
    65507 => 0,
    65508 => 0,
    65509 => 0,
    65510 => 0,
    65511 => 0,
    65512 => 0,
    65513 => 0,
    65514 => 0,
    65515 => 0,
    65516 => 0,
    65517 => 0,
    65518 => 0,
    65519 => 0,
    65520 => 0,
    65521 => 0,
    65522 => 0,
    65523 => 0,
    65524 => 0,
    65525 => 0,
    65526 => 0,
    65527 => 0,
    65528 => 0,
    65529 => 0,
    65530 => 0,
    65531 => 0,
    65532 => 0,
    65533 => 0,
    65534 => 0,
    65535 => 0
  );

begin
  lut_out <= std_logic_vector(to_signed(LUT(to_integer(unsigned(address))),P));
end architecture;
