library IEEE;
  use IEEE.std_logic_1164.all;
  use IEEE.numeric_std.all;

entity lut_table_16384_7bit is
  generic (
    N : integer := 14;
    P : integer := 7
  );
  port (
    address  : in  std_logic_vector(N-1 downto 0);
    lut_out : out std_logic_vector(P-1 downto 0)
  );
end entity;

architecture behavior of lut_table_16384_7bit is

  type LUT_t is array (natural range 0 to 16383) of integer;
  constant LUT: LUT_t := (
    0 => 0,
    1 => 0,
    2 => 0,
    3 => 0,
    4 => 0,
    5 => 0,
    6 => 0,
    7 => 0,
    8 => 0,
    9 => 0,
    10 => 0,
    11 => 0,
    12 => 0,
    13 => 0,
    14 => 0,
    15 => 0,
    16 => 0,
    17 => 0,
    18 => 0,
    19 => 0,
    20 => 0,
    21 => 1,
    22 => 1,
    23 => 1,
    24 => 1,
    25 => 1,
    26 => 1,
    27 => 1,
    28 => 1,
    29 => 1,
    30 => 1,
    31 => 1,
    32 => 1,
    33 => 1,
    34 => 1,
    35 => 1,
    36 => 1,
    37 => 1,
    38 => 1,
    39 => 1,
    40 => 1,
    41 => 1,
    42 => 1,
    43 => 1,
    44 => 1,
    45 => 1,
    46 => 1,
    47 => 1,
    48 => 1,
    49 => 1,
    50 => 1,
    51 => 1,
    52 => 1,
    53 => 1,
    54 => 1,
    55 => 1,
    56 => 1,
    57 => 1,
    58 => 1,
    59 => 1,
    60 => 1,
    61 => 1,
    62 => 1,
    63 => 2,
    64 => 2,
    65 => 2,
    66 => 2,
    67 => 2,
    68 => 2,
    69 => 2,
    70 => 2,
    71 => 2,
    72 => 2,
    73 => 2,
    74 => 2,
    75 => 2,
    76 => 2,
    77 => 2,
    78 => 2,
    79 => 2,
    80 => 2,
    81 => 2,
    82 => 2,
    83 => 2,
    84 => 2,
    85 => 2,
    86 => 2,
    87 => 2,
    88 => 2,
    89 => 2,
    90 => 2,
    91 => 2,
    92 => 2,
    93 => 2,
    94 => 2,
    95 => 2,
    96 => 2,
    97 => 2,
    98 => 2,
    99 => 2,
    100 => 2,
    101 => 2,
    102 => 2,
    103 => 2,
    104 => 3,
    105 => 3,
    106 => 3,
    107 => 3,
    108 => 3,
    109 => 3,
    110 => 3,
    111 => 3,
    112 => 3,
    113 => 3,
    114 => 3,
    115 => 3,
    116 => 3,
    117 => 3,
    118 => 3,
    119 => 3,
    120 => 3,
    121 => 3,
    122 => 3,
    123 => 3,
    124 => 3,
    125 => 3,
    126 => 3,
    127 => 3,
    128 => 3,
    129 => 3,
    130 => 3,
    131 => 3,
    132 => 3,
    133 => 3,
    134 => 3,
    135 => 3,
    136 => 3,
    137 => 3,
    138 => 3,
    139 => 3,
    140 => 3,
    141 => 3,
    142 => 3,
    143 => 3,
    144 => 3,
    145 => 4,
    146 => 4,
    147 => 4,
    148 => 4,
    149 => 4,
    150 => 4,
    151 => 4,
    152 => 4,
    153 => 4,
    154 => 4,
    155 => 4,
    156 => 4,
    157 => 4,
    158 => 4,
    159 => 4,
    160 => 4,
    161 => 4,
    162 => 4,
    163 => 4,
    164 => 4,
    165 => 4,
    166 => 4,
    167 => 4,
    168 => 4,
    169 => 4,
    170 => 4,
    171 => 4,
    172 => 4,
    173 => 4,
    174 => 4,
    175 => 4,
    176 => 4,
    177 => 4,
    178 => 4,
    179 => 4,
    180 => 4,
    181 => 4,
    182 => 4,
    183 => 4,
    184 => 4,
    185 => 4,
    186 => 4,
    187 => 5,
    188 => 5,
    189 => 5,
    190 => 5,
    191 => 5,
    192 => 5,
    193 => 5,
    194 => 5,
    195 => 5,
    196 => 5,
    197 => 5,
    198 => 5,
    199 => 5,
    200 => 5,
    201 => 5,
    202 => 5,
    203 => 5,
    204 => 5,
    205 => 5,
    206 => 5,
    207 => 5,
    208 => 5,
    209 => 5,
    210 => 5,
    211 => 5,
    212 => 5,
    213 => 5,
    214 => 5,
    215 => 5,
    216 => 5,
    217 => 5,
    218 => 5,
    219 => 5,
    220 => 5,
    221 => 5,
    222 => 5,
    223 => 5,
    224 => 5,
    225 => 5,
    226 => 5,
    227 => 5,
    228 => 6,
    229 => 6,
    230 => 6,
    231 => 6,
    232 => 6,
    233 => 6,
    234 => 6,
    235 => 6,
    236 => 6,
    237 => 6,
    238 => 6,
    239 => 6,
    240 => 6,
    241 => 6,
    242 => 6,
    243 => 6,
    244 => 6,
    245 => 6,
    246 => 6,
    247 => 6,
    248 => 6,
    249 => 6,
    250 => 6,
    251 => 6,
    252 => 6,
    253 => 6,
    254 => 6,
    255 => 6,
    256 => 6,
    257 => 6,
    258 => 6,
    259 => 6,
    260 => 6,
    261 => 6,
    262 => 6,
    263 => 6,
    264 => 6,
    265 => 6,
    266 => 6,
    267 => 6,
    268 => 6,
    269 => 6,
    270 => 7,
    271 => 7,
    272 => 7,
    273 => 7,
    274 => 7,
    275 => 7,
    276 => 7,
    277 => 7,
    278 => 7,
    279 => 7,
    280 => 7,
    281 => 7,
    282 => 7,
    283 => 7,
    284 => 7,
    285 => 7,
    286 => 7,
    287 => 7,
    288 => 7,
    289 => 7,
    290 => 7,
    291 => 7,
    292 => 7,
    293 => 7,
    294 => 7,
    295 => 7,
    296 => 7,
    297 => 7,
    298 => 7,
    299 => 7,
    300 => 7,
    301 => 7,
    302 => 7,
    303 => 7,
    304 => 7,
    305 => 7,
    306 => 7,
    307 => 7,
    308 => 7,
    309 => 7,
    310 => 7,
    311 => 7,
    312 => 8,
    313 => 8,
    314 => 8,
    315 => 8,
    316 => 8,
    317 => 8,
    318 => 8,
    319 => 8,
    320 => 8,
    321 => 8,
    322 => 8,
    323 => 8,
    324 => 8,
    325 => 8,
    326 => 8,
    327 => 8,
    328 => 8,
    329 => 8,
    330 => 8,
    331 => 8,
    332 => 8,
    333 => 8,
    334 => 8,
    335 => 8,
    336 => 8,
    337 => 8,
    338 => 8,
    339 => 8,
    340 => 8,
    341 => 8,
    342 => 8,
    343 => 8,
    344 => 8,
    345 => 8,
    346 => 8,
    347 => 8,
    348 => 8,
    349 => 8,
    350 => 8,
    351 => 8,
    352 => 8,
    353 => 9,
    354 => 9,
    355 => 9,
    356 => 9,
    357 => 9,
    358 => 9,
    359 => 9,
    360 => 9,
    361 => 9,
    362 => 9,
    363 => 9,
    364 => 9,
    365 => 9,
    366 => 9,
    367 => 9,
    368 => 9,
    369 => 9,
    370 => 9,
    371 => 9,
    372 => 9,
    373 => 9,
    374 => 9,
    375 => 9,
    376 => 9,
    377 => 9,
    378 => 9,
    379 => 9,
    380 => 9,
    381 => 9,
    382 => 9,
    383 => 9,
    384 => 9,
    385 => 9,
    386 => 9,
    387 => 9,
    388 => 9,
    389 => 9,
    390 => 9,
    391 => 9,
    392 => 9,
    393 => 9,
    394 => 9,
    395 => 10,
    396 => 10,
    397 => 10,
    398 => 10,
    399 => 10,
    400 => 10,
    401 => 10,
    402 => 10,
    403 => 10,
    404 => 10,
    405 => 10,
    406 => 10,
    407 => 10,
    408 => 10,
    409 => 10,
    410 => 10,
    411 => 10,
    412 => 10,
    413 => 10,
    414 => 10,
    415 => 10,
    416 => 10,
    417 => 10,
    418 => 10,
    419 => 10,
    420 => 10,
    421 => 10,
    422 => 10,
    423 => 10,
    424 => 10,
    425 => 10,
    426 => 10,
    427 => 10,
    428 => 10,
    429 => 10,
    430 => 10,
    431 => 10,
    432 => 10,
    433 => 10,
    434 => 10,
    435 => 10,
    436 => 10,
    437 => 11,
    438 => 11,
    439 => 11,
    440 => 11,
    441 => 11,
    442 => 11,
    443 => 11,
    444 => 11,
    445 => 11,
    446 => 11,
    447 => 11,
    448 => 11,
    449 => 11,
    450 => 11,
    451 => 11,
    452 => 11,
    453 => 11,
    454 => 11,
    455 => 11,
    456 => 11,
    457 => 11,
    458 => 11,
    459 => 11,
    460 => 11,
    461 => 11,
    462 => 11,
    463 => 11,
    464 => 11,
    465 => 11,
    466 => 11,
    467 => 11,
    468 => 11,
    469 => 11,
    470 => 11,
    471 => 11,
    472 => 11,
    473 => 11,
    474 => 11,
    475 => 11,
    476 => 11,
    477 => 11,
    478 => 11,
    479 => 12,
    480 => 12,
    481 => 12,
    482 => 12,
    483 => 12,
    484 => 12,
    485 => 12,
    486 => 12,
    487 => 12,
    488 => 12,
    489 => 12,
    490 => 12,
    491 => 12,
    492 => 12,
    493 => 12,
    494 => 12,
    495 => 12,
    496 => 12,
    497 => 12,
    498 => 12,
    499 => 12,
    500 => 12,
    501 => 12,
    502 => 12,
    503 => 12,
    504 => 12,
    505 => 12,
    506 => 12,
    507 => 12,
    508 => 12,
    509 => 12,
    510 => 12,
    511 => 12,
    512 => 12,
    513 => 12,
    514 => 12,
    515 => 12,
    516 => 12,
    517 => 12,
    518 => 12,
    519 => 12,
    520 => 12,
    521 => 13,
    522 => 13,
    523 => 13,
    524 => 13,
    525 => 13,
    526 => 13,
    527 => 13,
    528 => 13,
    529 => 13,
    530 => 13,
    531 => 13,
    532 => 13,
    533 => 13,
    534 => 13,
    535 => 13,
    536 => 13,
    537 => 13,
    538 => 13,
    539 => 13,
    540 => 13,
    541 => 13,
    542 => 13,
    543 => 13,
    544 => 13,
    545 => 13,
    546 => 13,
    547 => 13,
    548 => 13,
    549 => 13,
    550 => 13,
    551 => 13,
    552 => 13,
    553 => 13,
    554 => 13,
    555 => 13,
    556 => 13,
    557 => 13,
    558 => 13,
    559 => 13,
    560 => 13,
    561 => 13,
    562 => 13,
    563 => 13,
    564 => 14,
    565 => 14,
    566 => 14,
    567 => 14,
    568 => 14,
    569 => 14,
    570 => 14,
    571 => 14,
    572 => 14,
    573 => 14,
    574 => 14,
    575 => 14,
    576 => 14,
    577 => 14,
    578 => 14,
    579 => 14,
    580 => 14,
    581 => 14,
    582 => 14,
    583 => 14,
    584 => 14,
    585 => 14,
    586 => 14,
    587 => 14,
    588 => 14,
    589 => 14,
    590 => 14,
    591 => 14,
    592 => 14,
    593 => 14,
    594 => 14,
    595 => 14,
    596 => 14,
    597 => 14,
    598 => 14,
    599 => 14,
    600 => 14,
    601 => 14,
    602 => 14,
    603 => 14,
    604 => 14,
    605 => 14,
    606 => 15,
    607 => 15,
    608 => 15,
    609 => 15,
    610 => 15,
    611 => 15,
    612 => 15,
    613 => 15,
    614 => 15,
    615 => 15,
    616 => 15,
    617 => 15,
    618 => 15,
    619 => 15,
    620 => 15,
    621 => 15,
    622 => 15,
    623 => 15,
    624 => 15,
    625 => 15,
    626 => 15,
    627 => 15,
    628 => 15,
    629 => 15,
    630 => 15,
    631 => 15,
    632 => 15,
    633 => 15,
    634 => 15,
    635 => 15,
    636 => 15,
    637 => 15,
    638 => 15,
    639 => 15,
    640 => 15,
    641 => 15,
    642 => 15,
    643 => 15,
    644 => 15,
    645 => 15,
    646 => 15,
    647 => 15,
    648 => 15,
    649 => 16,
    650 => 16,
    651 => 16,
    652 => 16,
    653 => 16,
    654 => 16,
    655 => 16,
    656 => 16,
    657 => 16,
    658 => 16,
    659 => 16,
    660 => 16,
    661 => 16,
    662 => 16,
    663 => 16,
    664 => 16,
    665 => 16,
    666 => 16,
    667 => 16,
    668 => 16,
    669 => 16,
    670 => 16,
    671 => 16,
    672 => 16,
    673 => 16,
    674 => 16,
    675 => 16,
    676 => 16,
    677 => 16,
    678 => 16,
    679 => 16,
    680 => 16,
    681 => 16,
    682 => 16,
    683 => 16,
    684 => 16,
    685 => 16,
    686 => 16,
    687 => 16,
    688 => 16,
    689 => 16,
    690 => 16,
    691 => 16,
    692 => 17,
    693 => 17,
    694 => 17,
    695 => 17,
    696 => 17,
    697 => 17,
    698 => 17,
    699 => 17,
    700 => 17,
    701 => 17,
    702 => 17,
    703 => 17,
    704 => 17,
    705 => 17,
    706 => 17,
    707 => 17,
    708 => 17,
    709 => 17,
    710 => 17,
    711 => 17,
    712 => 17,
    713 => 17,
    714 => 17,
    715 => 17,
    716 => 17,
    717 => 17,
    718 => 17,
    719 => 17,
    720 => 17,
    721 => 17,
    722 => 17,
    723 => 17,
    724 => 17,
    725 => 17,
    726 => 17,
    727 => 17,
    728 => 17,
    729 => 17,
    730 => 17,
    731 => 17,
    732 => 17,
    733 => 17,
    734 => 18,
    735 => 18,
    736 => 18,
    737 => 18,
    738 => 18,
    739 => 18,
    740 => 18,
    741 => 18,
    742 => 18,
    743 => 18,
    744 => 18,
    745 => 18,
    746 => 18,
    747 => 18,
    748 => 18,
    749 => 18,
    750 => 18,
    751 => 18,
    752 => 18,
    753 => 18,
    754 => 18,
    755 => 18,
    756 => 18,
    757 => 18,
    758 => 18,
    759 => 18,
    760 => 18,
    761 => 18,
    762 => 18,
    763 => 18,
    764 => 18,
    765 => 18,
    766 => 18,
    767 => 18,
    768 => 18,
    769 => 18,
    770 => 18,
    771 => 18,
    772 => 18,
    773 => 18,
    774 => 18,
    775 => 18,
    776 => 18,
    777 => 18,
    778 => 19,
    779 => 19,
    780 => 19,
    781 => 19,
    782 => 19,
    783 => 19,
    784 => 19,
    785 => 19,
    786 => 19,
    787 => 19,
    788 => 19,
    789 => 19,
    790 => 19,
    791 => 19,
    792 => 19,
    793 => 19,
    794 => 19,
    795 => 19,
    796 => 19,
    797 => 19,
    798 => 19,
    799 => 19,
    800 => 19,
    801 => 19,
    802 => 19,
    803 => 19,
    804 => 19,
    805 => 19,
    806 => 19,
    807 => 19,
    808 => 19,
    809 => 19,
    810 => 19,
    811 => 19,
    812 => 19,
    813 => 19,
    814 => 19,
    815 => 19,
    816 => 19,
    817 => 19,
    818 => 19,
    819 => 19,
    820 => 19,
    821 => 20,
    822 => 20,
    823 => 20,
    824 => 20,
    825 => 20,
    826 => 20,
    827 => 20,
    828 => 20,
    829 => 20,
    830 => 20,
    831 => 20,
    832 => 20,
    833 => 20,
    834 => 20,
    835 => 20,
    836 => 20,
    837 => 20,
    838 => 20,
    839 => 20,
    840 => 20,
    841 => 20,
    842 => 20,
    843 => 20,
    844 => 20,
    845 => 20,
    846 => 20,
    847 => 20,
    848 => 20,
    849 => 20,
    850 => 20,
    851 => 20,
    852 => 20,
    853 => 20,
    854 => 20,
    855 => 20,
    856 => 20,
    857 => 20,
    858 => 20,
    859 => 20,
    860 => 20,
    861 => 20,
    862 => 20,
    863 => 20,
    864 => 20,
    865 => 21,
    866 => 21,
    867 => 21,
    868 => 21,
    869 => 21,
    870 => 21,
    871 => 21,
    872 => 21,
    873 => 21,
    874 => 21,
    875 => 21,
    876 => 21,
    877 => 21,
    878 => 21,
    879 => 21,
    880 => 21,
    881 => 21,
    882 => 21,
    883 => 21,
    884 => 21,
    885 => 21,
    886 => 21,
    887 => 21,
    888 => 21,
    889 => 21,
    890 => 21,
    891 => 21,
    892 => 21,
    893 => 21,
    894 => 21,
    895 => 21,
    896 => 21,
    897 => 21,
    898 => 21,
    899 => 21,
    900 => 21,
    901 => 21,
    902 => 21,
    903 => 21,
    904 => 21,
    905 => 21,
    906 => 21,
    907 => 21,
    908 => 21,
    909 => 22,
    910 => 22,
    911 => 22,
    912 => 22,
    913 => 22,
    914 => 22,
    915 => 22,
    916 => 22,
    917 => 22,
    918 => 22,
    919 => 22,
    920 => 22,
    921 => 22,
    922 => 22,
    923 => 22,
    924 => 22,
    925 => 22,
    926 => 22,
    927 => 22,
    928 => 22,
    929 => 22,
    930 => 22,
    931 => 22,
    932 => 22,
    933 => 22,
    934 => 22,
    935 => 22,
    936 => 22,
    937 => 22,
    938 => 22,
    939 => 22,
    940 => 22,
    941 => 22,
    942 => 22,
    943 => 22,
    944 => 22,
    945 => 22,
    946 => 22,
    947 => 22,
    948 => 22,
    949 => 22,
    950 => 22,
    951 => 22,
    952 => 22,
    953 => 23,
    954 => 23,
    955 => 23,
    956 => 23,
    957 => 23,
    958 => 23,
    959 => 23,
    960 => 23,
    961 => 23,
    962 => 23,
    963 => 23,
    964 => 23,
    965 => 23,
    966 => 23,
    967 => 23,
    968 => 23,
    969 => 23,
    970 => 23,
    971 => 23,
    972 => 23,
    973 => 23,
    974 => 23,
    975 => 23,
    976 => 23,
    977 => 23,
    978 => 23,
    979 => 23,
    980 => 23,
    981 => 23,
    982 => 23,
    983 => 23,
    984 => 23,
    985 => 23,
    986 => 23,
    987 => 23,
    988 => 23,
    989 => 23,
    990 => 23,
    991 => 23,
    992 => 23,
    993 => 23,
    994 => 23,
    995 => 23,
    996 => 23,
    997 => 24,
    998 => 24,
    999 => 24,
    1000 => 24,
    1001 => 24,
    1002 => 24,
    1003 => 24,
    1004 => 24,
    1005 => 24,
    1006 => 24,
    1007 => 24,
    1008 => 24,
    1009 => 24,
    1010 => 24,
    1011 => 24,
    1012 => 24,
    1013 => 24,
    1014 => 24,
    1015 => 24,
    1016 => 24,
    1017 => 24,
    1018 => 24,
    1019 => 24,
    1020 => 24,
    1021 => 24,
    1022 => 24,
    1023 => 24,
    1024 => 24,
    1025 => 24,
    1026 => 24,
    1027 => 24,
    1028 => 24,
    1029 => 24,
    1030 => 24,
    1031 => 24,
    1032 => 24,
    1033 => 24,
    1034 => 24,
    1035 => 24,
    1036 => 24,
    1037 => 24,
    1038 => 24,
    1039 => 24,
    1040 => 24,
    1041 => 24,
    1042 => 25,
    1043 => 25,
    1044 => 25,
    1045 => 25,
    1046 => 25,
    1047 => 25,
    1048 => 25,
    1049 => 25,
    1050 => 25,
    1051 => 25,
    1052 => 25,
    1053 => 25,
    1054 => 25,
    1055 => 25,
    1056 => 25,
    1057 => 25,
    1058 => 25,
    1059 => 25,
    1060 => 25,
    1061 => 25,
    1062 => 25,
    1063 => 25,
    1064 => 25,
    1065 => 25,
    1066 => 25,
    1067 => 25,
    1068 => 25,
    1069 => 25,
    1070 => 25,
    1071 => 25,
    1072 => 25,
    1073 => 25,
    1074 => 25,
    1075 => 25,
    1076 => 25,
    1077 => 25,
    1078 => 25,
    1079 => 25,
    1080 => 25,
    1081 => 25,
    1082 => 25,
    1083 => 25,
    1084 => 25,
    1085 => 25,
    1086 => 25,
    1087 => 26,
    1088 => 26,
    1089 => 26,
    1090 => 26,
    1091 => 26,
    1092 => 26,
    1093 => 26,
    1094 => 26,
    1095 => 26,
    1096 => 26,
    1097 => 26,
    1098 => 26,
    1099 => 26,
    1100 => 26,
    1101 => 26,
    1102 => 26,
    1103 => 26,
    1104 => 26,
    1105 => 26,
    1106 => 26,
    1107 => 26,
    1108 => 26,
    1109 => 26,
    1110 => 26,
    1111 => 26,
    1112 => 26,
    1113 => 26,
    1114 => 26,
    1115 => 26,
    1116 => 26,
    1117 => 26,
    1118 => 26,
    1119 => 26,
    1120 => 26,
    1121 => 26,
    1122 => 26,
    1123 => 26,
    1124 => 26,
    1125 => 26,
    1126 => 26,
    1127 => 26,
    1128 => 26,
    1129 => 26,
    1130 => 26,
    1131 => 26,
    1132 => 26,
    1133 => 27,
    1134 => 27,
    1135 => 27,
    1136 => 27,
    1137 => 27,
    1138 => 27,
    1139 => 27,
    1140 => 27,
    1141 => 27,
    1142 => 27,
    1143 => 27,
    1144 => 27,
    1145 => 27,
    1146 => 27,
    1147 => 27,
    1148 => 27,
    1149 => 27,
    1150 => 27,
    1151 => 27,
    1152 => 27,
    1153 => 27,
    1154 => 27,
    1155 => 27,
    1156 => 27,
    1157 => 27,
    1158 => 27,
    1159 => 27,
    1160 => 27,
    1161 => 27,
    1162 => 27,
    1163 => 27,
    1164 => 27,
    1165 => 27,
    1166 => 27,
    1167 => 27,
    1168 => 27,
    1169 => 27,
    1170 => 27,
    1171 => 27,
    1172 => 27,
    1173 => 27,
    1174 => 27,
    1175 => 27,
    1176 => 27,
    1177 => 27,
    1178 => 28,
    1179 => 28,
    1180 => 28,
    1181 => 28,
    1182 => 28,
    1183 => 28,
    1184 => 28,
    1185 => 28,
    1186 => 28,
    1187 => 28,
    1188 => 28,
    1189 => 28,
    1190 => 28,
    1191 => 28,
    1192 => 28,
    1193 => 28,
    1194 => 28,
    1195 => 28,
    1196 => 28,
    1197 => 28,
    1198 => 28,
    1199 => 28,
    1200 => 28,
    1201 => 28,
    1202 => 28,
    1203 => 28,
    1204 => 28,
    1205 => 28,
    1206 => 28,
    1207 => 28,
    1208 => 28,
    1209 => 28,
    1210 => 28,
    1211 => 28,
    1212 => 28,
    1213 => 28,
    1214 => 28,
    1215 => 28,
    1216 => 28,
    1217 => 28,
    1218 => 28,
    1219 => 28,
    1220 => 28,
    1221 => 28,
    1222 => 28,
    1223 => 28,
    1224 => 28,
    1225 => 29,
    1226 => 29,
    1227 => 29,
    1228 => 29,
    1229 => 29,
    1230 => 29,
    1231 => 29,
    1232 => 29,
    1233 => 29,
    1234 => 29,
    1235 => 29,
    1236 => 29,
    1237 => 29,
    1238 => 29,
    1239 => 29,
    1240 => 29,
    1241 => 29,
    1242 => 29,
    1243 => 29,
    1244 => 29,
    1245 => 29,
    1246 => 29,
    1247 => 29,
    1248 => 29,
    1249 => 29,
    1250 => 29,
    1251 => 29,
    1252 => 29,
    1253 => 29,
    1254 => 29,
    1255 => 29,
    1256 => 29,
    1257 => 29,
    1258 => 29,
    1259 => 29,
    1260 => 29,
    1261 => 29,
    1262 => 29,
    1263 => 29,
    1264 => 29,
    1265 => 29,
    1266 => 29,
    1267 => 29,
    1268 => 29,
    1269 => 29,
    1270 => 29,
    1271 => 30,
    1272 => 30,
    1273 => 30,
    1274 => 30,
    1275 => 30,
    1276 => 30,
    1277 => 30,
    1278 => 30,
    1279 => 30,
    1280 => 30,
    1281 => 30,
    1282 => 30,
    1283 => 30,
    1284 => 30,
    1285 => 30,
    1286 => 30,
    1287 => 30,
    1288 => 30,
    1289 => 30,
    1290 => 30,
    1291 => 30,
    1292 => 30,
    1293 => 30,
    1294 => 30,
    1295 => 30,
    1296 => 30,
    1297 => 30,
    1298 => 30,
    1299 => 30,
    1300 => 30,
    1301 => 30,
    1302 => 30,
    1303 => 30,
    1304 => 30,
    1305 => 30,
    1306 => 30,
    1307 => 30,
    1308 => 30,
    1309 => 30,
    1310 => 30,
    1311 => 30,
    1312 => 30,
    1313 => 30,
    1314 => 30,
    1315 => 30,
    1316 => 30,
    1317 => 30,
    1318 => 31,
    1319 => 31,
    1320 => 31,
    1321 => 31,
    1322 => 31,
    1323 => 31,
    1324 => 31,
    1325 => 31,
    1326 => 31,
    1327 => 31,
    1328 => 31,
    1329 => 31,
    1330 => 31,
    1331 => 31,
    1332 => 31,
    1333 => 31,
    1334 => 31,
    1335 => 31,
    1336 => 31,
    1337 => 31,
    1338 => 31,
    1339 => 31,
    1340 => 31,
    1341 => 31,
    1342 => 31,
    1343 => 31,
    1344 => 31,
    1345 => 31,
    1346 => 31,
    1347 => 31,
    1348 => 31,
    1349 => 31,
    1350 => 31,
    1351 => 31,
    1352 => 31,
    1353 => 31,
    1354 => 31,
    1355 => 31,
    1356 => 31,
    1357 => 31,
    1358 => 31,
    1359 => 31,
    1360 => 31,
    1361 => 31,
    1362 => 31,
    1363 => 31,
    1364 => 31,
    1365 => 31,
    1366 => 32,
    1367 => 32,
    1368 => 32,
    1369 => 32,
    1370 => 32,
    1371 => 32,
    1372 => 32,
    1373 => 32,
    1374 => 32,
    1375 => 32,
    1376 => 32,
    1377 => 32,
    1378 => 32,
    1379 => 32,
    1380 => 32,
    1381 => 32,
    1382 => 32,
    1383 => 32,
    1384 => 32,
    1385 => 32,
    1386 => 32,
    1387 => 32,
    1388 => 32,
    1389 => 32,
    1390 => 32,
    1391 => 32,
    1392 => 32,
    1393 => 32,
    1394 => 32,
    1395 => 32,
    1396 => 32,
    1397 => 32,
    1398 => 32,
    1399 => 32,
    1400 => 32,
    1401 => 32,
    1402 => 32,
    1403 => 32,
    1404 => 32,
    1405 => 32,
    1406 => 32,
    1407 => 32,
    1408 => 32,
    1409 => 32,
    1410 => 32,
    1411 => 32,
    1412 => 32,
    1413 => 32,
    1414 => 33,
    1415 => 33,
    1416 => 33,
    1417 => 33,
    1418 => 33,
    1419 => 33,
    1420 => 33,
    1421 => 33,
    1422 => 33,
    1423 => 33,
    1424 => 33,
    1425 => 33,
    1426 => 33,
    1427 => 33,
    1428 => 33,
    1429 => 33,
    1430 => 33,
    1431 => 33,
    1432 => 33,
    1433 => 33,
    1434 => 33,
    1435 => 33,
    1436 => 33,
    1437 => 33,
    1438 => 33,
    1439 => 33,
    1440 => 33,
    1441 => 33,
    1442 => 33,
    1443 => 33,
    1444 => 33,
    1445 => 33,
    1446 => 33,
    1447 => 33,
    1448 => 33,
    1449 => 33,
    1450 => 33,
    1451 => 33,
    1452 => 33,
    1453 => 33,
    1454 => 33,
    1455 => 33,
    1456 => 33,
    1457 => 33,
    1458 => 33,
    1459 => 33,
    1460 => 33,
    1461 => 33,
    1462 => 34,
    1463 => 34,
    1464 => 34,
    1465 => 34,
    1466 => 34,
    1467 => 34,
    1468 => 34,
    1469 => 34,
    1470 => 34,
    1471 => 34,
    1472 => 34,
    1473 => 34,
    1474 => 34,
    1475 => 34,
    1476 => 34,
    1477 => 34,
    1478 => 34,
    1479 => 34,
    1480 => 34,
    1481 => 34,
    1482 => 34,
    1483 => 34,
    1484 => 34,
    1485 => 34,
    1486 => 34,
    1487 => 34,
    1488 => 34,
    1489 => 34,
    1490 => 34,
    1491 => 34,
    1492 => 34,
    1493 => 34,
    1494 => 34,
    1495 => 34,
    1496 => 34,
    1497 => 34,
    1498 => 34,
    1499 => 34,
    1500 => 34,
    1501 => 34,
    1502 => 34,
    1503 => 34,
    1504 => 34,
    1505 => 34,
    1506 => 34,
    1507 => 34,
    1508 => 34,
    1509 => 34,
    1510 => 34,
    1511 => 34,
    1512 => 35,
    1513 => 35,
    1514 => 35,
    1515 => 35,
    1516 => 35,
    1517 => 35,
    1518 => 35,
    1519 => 35,
    1520 => 35,
    1521 => 35,
    1522 => 35,
    1523 => 35,
    1524 => 35,
    1525 => 35,
    1526 => 35,
    1527 => 35,
    1528 => 35,
    1529 => 35,
    1530 => 35,
    1531 => 35,
    1532 => 35,
    1533 => 35,
    1534 => 35,
    1535 => 35,
    1536 => 35,
    1537 => 35,
    1538 => 35,
    1539 => 35,
    1540 => 35,
    1541 => 35,
    1542 => 35,
    1543 => 35,
    1544 => 35,
    1545 => 35,
    1546 => 35,
    1547 => 35,
    1548 => 35,
    1549 => 35,
    1550 => 35,
    1551 => 35,
    1552 => 35,
    1553 => 35,
    1554 => 35,
    1555 => 35,
    1556 => 35,
    1557 => 35,
    1558 => 35,
    1559 => 35,
    1560 => 35,
    1561 => 36,
    1562 => 36,
    1563 => 36,
    1564 => 36,
    1565 => 36,
    1566 => 36,
    1567 => 36,
    1568 => 36,
    1569 => 36,
    1570 => 36,
    1571 => 36,
    1572 => 36,
    1573 => 36,
    1574 => 36,
    1575 => 36,
    1576 => 36,
    1577 => 36,
    1578 => 36,
    1579 => 36,
    1580 => 36,
    1581 => 36,
    1582 => 36,
    1583 => 36,
    1584 => 36,
    1585 => 36,
    1586 => 36,
    1587 => 36,
    1588 => 36,
    1589 => 36,
    1590 => 36,
    1591 => 36,
    1592 => 36,
    1593 => 36,
    1594 => 36,
    1595 => 36,
    1596 => 36,
    1597 => 36,
    1598 => 36,
    1599 => 36,
    1600 => 36,
    1601 => 36,
    1602 => 36,
    1603 => 36,
    1604 => 36,
    1605 => 36,
    1606 => 36,
    1607 => 36,
    1608 => 36,
    1609 => 36,
    1610 => 36,
    1611 => 36,
    1612 => 37,
    1613 => 37,
    1614 => 37,
    1615 => 37,
    1616 => 37,
    1617 => 37,
    1618 => 37,
    1619 => 37,
    1620 => 37,
    1621 => 37,
    1622 => 37,
    1623 => 37,
    1624 => 37,
    1625 => 37,
    1626 => 37,
    1627 => 37,
    1628 => 37,
    1629 => 37,
    1630 => 37,
    1631 => 37,
    1632 => 37,
    1633 => 37,
    1634 => 37,
    1635 => 37,
    1636 => 37,
    1637 => 37,
    1638 => 37,
    1639 => 37,
    1640 => 37,
    1641 => 37,
    1642 => 37,
    1643 => 37,
    1644 => 37,
    1645 => 37,
    1646 => 37,
    1647 => 37,
    1648 => 37,
    1649 => 37,
    1650 => 37,
    1651 => 37,
    1652 => 37,
    1653 => 37,
    1654 => 37,
    1655 => 37,
    1656 => 37,
    1657 => 37,
    1658 => 37,
    1659 => 37,
    1660 => 37,
    1661 => 37,
    1662 => 37,
    1663 => 38,
    1664 => 38,
    1665 => 38,
    1666 => 38,
    1667 => 38,
    1668 => 38,
    1669 => 38,
    1670 => 38,
    1671 => 38,
    1672 => 38,
    1673 => 38,
    1674 => 38,
    1675 => 38,
    1676 => 38,
    1677 => 38,
    1678 => 38,
    1679 => 38,
    1680 => 38,
    1681 => 38,
    1682 => 38,
    1683 => 38,
    1684 => 38,
    1685 => 38,
    1686 => 38,
    1687 => 38,
    1688 => 38,
    1689 => 38,
    1690 => 38,
    1691 => 38,
    1692 => 38,
    1693 => 38,
    1694 => 38,
    1695 => 38,
    1696 => 38,
    1697 => 38,
    1698 => 38,
    1699 => 38,
    1700 => 38,
    1701 => 38,
    1702 => 38,
    1703 => 38,
    1704 => 38,
    1705 => 38,
    1706 => 38,
    1707 => 38,
    1708 => 38,
    1709 => 38,
    1710 => 38,
    1711 => 38,
    1712 => 38,
    1713 => 38,
    1714 => 38,
    1715 => 39,
    1716 => 39,
    1717 => 39,
    1718 => 39,
    1719 => 39,
    1720 => 39,
    1721 => 39,
    1722 => 39,
    1723 => 39,
    1724 => 39,
    1725 => 39,
    1726 => 39,
    1727 => 39,
    1728 => 39,
    1729 => 39,
    1730 => 39,
    1731 => 39,
    1732 => 39,
    1733 => 39,
    1734 => 39,
    1735 => 39,
    1736 => 39,
    1737 => 39,
    1738 => 39,
    1739 => 39,
    1740 => 39,
    1741 => 39,
    1742 => 39,
    1743 => 39,
    1744 => 39,
    1745 => 39,
    1746 => 39,
    1747 => 39,
    1748 => 39,
    1749 => 39,
    1750 => 39,
    1751 => 39,
    1752 => 39,
    1753 => 39,
    1754 => 39,
    1755 => 39,
    1756 => 39,
    1757 => 39,
    1758 => 39,
    1759 => 39,
    1760 => 39,
    1761 => 39,
    1762 => 39,
    1763 => 39,
    1764 => 39,
    1765 => 39,
    1766 => 39,
    1767 => 39,
    1768 => 40,
    1769 => 40,
    1770 => 40,
    1771 => 40,
    1772 => 40,
    1773 => 40,
    1774 => 40,
    1775 => 40,
    1776 => 40,
    1777 => 40,
    1778 => 40,
    1779 => 40,
    1780 => 40,
    1781 => 40,
    1782 => 40,
    1783 => 40,
    1784 => 40,
    1785 => 40,
    1786 => 40,
    1787 => 40,
    1788 => 40,
    1789 => 40,
    1790 => 40,
    1791 => 40,
    1792 => 40,
    1793 => 40,
    1794 => 40,
    1795 => 40,
    1796 => 40,
    1797 => 40,
    1798 => 40,
    1799 => 40,
    1800 => 40,
    1801 => 40,
    1802 => 40,
    1803 => 40,
    1804 => 40,
    1805 => 40,
    1806 => 40,
    1807 => 40,
    1808 => 40,
    1809 => 40,
    1810 => 40,
    1811 => 40,
    1812 => 40,
    1813 => 40,
    1814 => 40,
    1815 => 40,
    1816 => 40,
    1817 => 40,
    1818 => 40,
    1819 => 40,
    1820 => 40,
    1821 => 41,
    1822 => 41,
    1823 => 41,
    1824 => 41,
    1825 => 41,
    1826 => 41,
    1827 => 41,
    1828 => 41,
    1829 => 41,
    1830 => 41,
    1831 => 41,
    1832 => 41,
    1833 => 41,
    1834 => 41,
    1835 => 41,
    1836 => 41,
    1837 => 41,
    1838 => 41,
    1839 => 41,
    1840 => 41,
    1841 => 41,
    1842 => 41,
    1843 => 41,
    1844 => 41,
    1845 => 41,
    1846 => 41,
    1847 => 41,
    1848 => 41,
    1849 => 41,
    1850 => 41,
    1851 => 41,
    1852 => 41,
    1853 => 41,
    1854 => 41,
    1855 => 41,
    1856 => 41,
    1857 => 41,
    1858 => 41,
    1859 => 41,
    1860 => 41,
    1861 => 41,
    1862 => 41,
    1863 => 41,
    1864 => 41,
    1865 => 41,
    1866 => 41,
    1867 => 41,
    1868 => 41,
    1869 => 41,
    1870 => 41,
    1871 => 41,
    1872 => 41,
    1873 => 41,
    1874 => 41,
    1875 => 41,
    1876 => 42,
    1877 => 42,
    1878 => 42,
    1879 => 42,
    1880 => 42,
    1881 => 42,
    1882 => 42,
    1883 => 42,
    1884 => 42,
    1885 => 42,
    1886 => 42,
    1887 => 42,
    1888 => 42,
    1889 => 42,
    1890 => 42,
    1891 => 42,
    1892 => 42,
    1893 => 42,
    1894 => 42,
    1895 => 42,
    1896 => 42,
    1897 => 42,
    1898 => 42,
    1899 => 42,
    1900 => 42,
    1901 => 42,
    1902 => 42,
    1903 => 42,
    1904 => 42,
    1905 => 42,
    1906 => 42,
    1907 => 42,
    1908 => 42,
    1909 => 42,
    1910 => 42,
    1911 => 42,
    1912 => 42,
    1913 => 42,
    1914 => 42,
    1915 => 42,
    1916 => 42,
    1917 => 42,
    1918 => 42,
    1919 => 42,
    1920 => 42,
    1921 => 42,
    1922 => 42,
    1923 => 42,
    1924 => 42,
    1925 => 42,
    1926 => 42,
    1927 => 42,
    1928 => 42,
    1929 => 42,
    1930 => 42,
    1931 => 43,
    1932 => 43,
    1933 => 43,
    1934 => 43,
    1935 => 43,
    1936 => 43,
    1937 => 43,
    1938 => 43,
    1939 => 43,
    1940 => 43,
    1941 => 43,
    1942 => 43,
    1943 => 43,
    1944 => 43,
    1945 => 43,
    1946 => 43,
    1947 => 43,
    1948 => 43,
    1949 => 43,
    1950 => 43,
    1951 => 43,
    1952 => 43,
    1953 => 43,
    1954 => 43,
    1955 => 43,
    1956 => 43,
    1957 => 43,
    1958 => 43,
    1959 => 43,
    1960 => 43,
    1961 => 43,
    1962 => 43,
    1963 => 43,
    1964 => 43,
    1965 => 43,
    1966 => 43,
    1967 => 43,
    1968 => 43,
    1969 => 43,
    1970 => 43,
    1971 => 43,
    1972 => 43,
    1973 => 43,
    1974 => 43,
    1975 => 43,
    1976 => 43,
    1977 => 43,
    1978 => 43,
    1979 => 43,
    1980 => 43,
    1981 => 43,
    1982 => 43,
    1983 => 43,
    1984 => 43,
    1985 => 43,
    1986 => 43,
    1987 => 43,
    1988 => 44,
    1989 => 44,
    1990 => 44,
    1991 => 44,
    1992 => 44,
    1993 => 44,
    1994 => 44,
    1995 => 44,
    1996 => 44,
    1997 => 44,
    1998 => 44,
    1999 => 44,
    2000 => 44,
    2001 => 44,
    2002 => 44,
    2003 => 44,
    2004 => 44,
    2005 => 44,
    2006 => 44,
    2007 => 44,
    2008 => 44,
    2009 => 44,
    2010 => 44,
    2011 => 44,
    2012 => 44,
    2013 => 44,
    2014 => 44,
    2015 => 44,
    2016 => 44,
    2017 => 44,
    2018 => 44,
    2019 => 44,
    2020 => 44,
    2021 => 44,
    2022 => 44,
    2023 => 44,
    2024 => 44,
    2025 => 44,
    2026 => 44,
    2027 => 44,
    2028 => 44,
    2029 => 44,
    2030 => 44,
    2031 => 44,
    2032 => 44,
    2033 => 44,
    2034 => 44,
    2035 => 44,
    2036 => 44,
    2037 => 44,
    2038 => 44,
    2039 => 44,
    2040 => 44,
    2041 => 44,
    2042 => 44,
    2043 => 44,
    2044 => 44,
    2045 => 44,
    2046 => 45,
    2047 => 45,
    2048 => 45,
    2049 => 45,
    2050 => 45,
    2051 => 45,
    2052 => 45,
    2053 => 45,
    2054 => 45,
    2055 => 45,
    2056 => 45,
    2057 => 45,
    2058 => 45,
    2059 => 45,
    2060 => 45,
    2061 => 45,
    2062 => 45,
    2063 => 45,
    2064 => 45,
    2065 => 45,
    2066 => 45,
    2067 => 45,
    2068 => 45,
    2069 => 45,
    2070 => 45,
    2071 => 45,
    2072 => 45,
    2073 => 45,
    2074 => 45,
    2075 => 45,
    2076 => 45,
    2077 => 45,
    2078 => 45,
    2079 => 45,
    2080 => 45,
    2081 => 45,
    2082 => 45,
    2083 => 45,
    2084 => 45,
    2085 => 45,
    2086 => 45,
    2087 => 45,
    2088 => 45,
    2089 => 45,
    2090 => 45,
    2091 => 45,
    2092 => 45,
    2093 => 45,
    2094 => 45,
    2095 => 45,
    2096 => 45,
    2097 => 45,
    2098 => 45,
    2099 => 45,
    2100 => 45,
    2101 => 45,
    2102 => 45,
    2103 => 45,
    2104 => 45,
    2105 => 46,
    2106 => 46,
    2107 => 46,
    2108 => 46,
    2109 => 46,
    2110 => 46,
    2111 => 46,
    2112 => 46,
    2113 => 46,
    2114 => 46,
    2115 => 46,
    2116 => 46,
    2117 => 46,
    2118 => 46,
    2119 => 46,
    2120 => 46,
    2121 => 46,
    2122 => 46,
    2123 => 46,
    2124 => 46,
    2125 => 46,
    2126 => 46,
    2127 => 46,
    2128 => 46,
    2129 => 46,
    2130 => 46,
    2131 => 46,
    2132 => 46,
    2133 => 46,
    2134 => 46,
    2135 => 46,
    2136 => 46,
    2137 => 46,
    2138 => 46,
    2139 => 46,
    2140 => 46,
    2141 => 46,
    2142 => 46,
    2143 => 46,
    2144 => 46,
    2145 => 46,
    2146 => 46,
    2147 => 46,
    2148 => 46,
    2149 => 46,
    2150 => 46,
    2151 => 46,
    2152 => 46,
    2153 => 46,
    2154 => 46,
    2155 => 46,
    2156 => 46,
    2157 => 46,
    2158 => 46,
    2159 => 46,
    2160 => 46,
    2161 => 46,
    2162 => 46,
    2163 => 46,
    2164 => 46,
    2165 => 47,
    2166 => 47,
    2167 => 47,
    2168 => 47,
    2169 => 47,
    2170 => 47,
    2171 => 47,
    2172 => 47,
    2173 => 47,
    2174 => 47,
    2175 => 47,
    2176 => 47,
    2177 => 47,
    2178 => 47,
    2179 => 47,
    2180 => 47,
    2181 => 47,
    2182 => 47,
    2183 => 47,
    2184 => 47,
    2185 => 47,
    2186 => 47,
    2187 => 47,
    2188 => 47,
    2189 => 47,
    2190 => 47,
    2191 => 47,
    2192 => 47,
    2193 => 47,
    2194 => 47,
    2195 => 47,
    2196 => 47,
    2197 => 47,
    2198 => 47,
    2199 => 47,
    2200 => 47,
    2201 => 47,
    2202 => 47,
    2203 => 47,
    2204 => 47,
    2205 => 47,
    2206 => 47,
    2207 => 47,
    2208 => 47,
    2209 => 47,
    2210 => 47,
    2211 => 47,
    2212 => 47,
    2213 => 47,
    2214 => 47,
    2215 => 47,
    2216 => 47,
    2217 => 47,
    2218 => 47,
    2219 => 47,
    2220 => 47,
    2221 => 47,
    2222 => 47,
    2223 => 47,
    2224 => 47,
    2225 => 47,
    2226 => 47,
    2227 => 47,
    2228 => 48,
    2229 => 48,
    2230 => 48,
    2231 => 48,
    2232 => 48,
    2233 => 48,
    2234 => 48,
    2235 => 48,
    2236 => 48,
    2237 => 48,
    2238 => 48,
    2239 => 48,
    2240 => 48,
    2241 => 48,
    2242 => 48,
    2243 => 48,
    2244 => 48,
    2245 => 48,
    2246 => 48,
    2247 => 48,
    2248 => 48,
    2249 => 48,
    2250 => 48,
    2251 => 48,
    2252 => 48,
    2253 => 48,
    2254 => 48,
    2255 => 48,
    2256 => 48,
    2257 => 48,
    2258 => 48,
    2259 => 48,
    2260 => 48,
    2261 => 48,
    2262 => 48,
    2263 => 48,
    2264 => 48,
    2265 => 48,
    2266 => 48,
    2267 => 48,
    2268 => 48,
    2269 => 48,
    2270 => 48,
    2271 => 48,
    2272 => 48,
    2273 => 48,
    2274 => 48,
    2275 => 48,
    2276 => 48,
    2277 => 48,
    2278 => 48,
    2279 => 48,
    2280 => 48,
    2281 => 48,
    2282 => 48,
    2283 => 48,
    2284 => 48,
    2285 => 48,
    2286 => 48,
    2287 => 48,
    2288 => 48,
    2289 => 48,
    2290 => 48,
    2291 => 48,
    2292 => 49,
    2293 => 49,
    2294 => 49,
    2295 => 49,
    2296 => 49,
    2297 => 49,
    2298 => 49,
    2299 => 49,
    2300 => 49,
    2301 => 49,
    2302 => 49,
    2303 => 49,
    2304 => 49,
    2305 => 49,
    2306 => 49,
    2307 => 49,
    2308 => 49,
    2309 => 49,
    2310 => 49,
    2311 => 49,
    2312 => 49,
    2313 => 49,
    2314 => 49,
    2315 => 49,
    2316 => 49,
    2317 => 49,
    2318 => 49,
    2319 => 49,
    2320 => 49,
    2321 => 49,
    2322 => 49,
    2323 => 49,
    2324 => 49,
    2325 => 49,
    2326 => 49,
    2327 => 49,
    2328 => 49,
    2329 => 49,
    2330 => 49,
    2331 => 49,
    2332 => 49,
    2333 => 49,
    2334 => 49,
    2335 => 49,
    2336 => 49,
    2337 => 49,
    2338 => 49,
    2339 => 49,
    2340 => 49,
    2341 => 49,
    2342 => 49,
    2343 => 49,
    2344 => 49,
    2345 => 49,
    2346 => 49,
    2347 => 49,
    2348 => 49,
    2349 => 49,
    2350 => 49,
    2351 => 49,
    2352 => 49,
    2353 => 49,
    2354 => 49,
    2355 => 49,
    2356 => 49,
    2357 => 50,
    2358 => 50,
    2359 => 50,
    2360 => 50,
    2361 => 50,
    2362 => 50,
    2363 => 50,
    2364 => 50,
    2365 => 50,
    2366 => 50,
    2367 => 50,
    2368 => 50,
    2369 => 50,
    2370 => 50,
    2371 => 50,
    2372 => 50,
    2373 => 50,
    2374 => 50,
    2375 => 50,
    2376 => 50,
    2377 => 50,
    2378 => 50,
    2379 => 50,
    2380 => 50,
    2381 => 50,
    2382 => 50,
    2383 => 50,
    2384 => 50,
    2385 => 50,
    2386 => 50,
    2387 => 50,
    2388 => 50,
    2389 => 50,
    2390 => 50,
    2391 => 50,
    2392 => 50,
    2393 => 50,
    2394 => 50,
    2395 => 50,
    2396 => 50,
    2397 => 50,
    2398 => 50,
    2399 => 50,
    2400 => 50,
    2401 => 50,
    2402 => 50,
    2403 => 50,
    2404 => 50,
    2405 => 50,
    2406 => 50,
    2407 => 50,
    2408 => 50,
    2409 => 50,
    2410 => 50,
    2411 => 50,
    2412 => 50,
    2413 => 50,
    2414 => 50,
    2415 => 50,
    2416 => 50,
    2417 => 50,
    2418 => 50,
    2419 => 50,
    2420 => 50,
    2421 => 50,
    2422 => 50,
    2423 => 50,
    2424 => 50,
    2425 => 51,
    2426 => 51,
    2427 => 51,
    2428 => 51,
    2429 => 51,
    2430 => 51,
    2431 => 51,
    2432 => 51,
    2433 => 51,
    2434 => 51,
    2435 => 51,
    2436 => 51,
    2437 => 51,
    2438 => 51,
    2439 => 51,
    2440 => 51,
    2441 => 51,
    2442 => 51,
    2443 => 51,
    2444 => 51,
    2445 => 51,
    2446 => 51,
    2447 => 51,
    2448 => 51,
    2449 => 51,
    2450 => 51,
    2451 => 51,
    2452 => 51,
    2453 => 51,
    2454 => 51,
    2455 => 51,
    2456 => 51,
    2457 => 51,
    2458 => 51,
    2459 => 51,
    2460 => 51,
    2461 => 51,
    2462 => 51,
    2463 => 51,
    2464 => 51,
    2465 => 51,
    2466 => 51,
    2467 => 51,
    2468 => 51,
    2469 => 51,
    2470 => 51,
    2471 => 51,
    2472 => 51,
    2473 => 51,
    2474 => 51,
    2475 => 51,
    2476 => 51,
    2477 => 51,
    2478 => 51,
    2479 => 51,
    2480 => 51,
    2481 => 51,
    2482 => 51,
    2483 => 51,
    2484 => 51,
    2485 => 51,
    2486 => 51,
    2487 => 51,
    2488 => 51,
    2489 => 51,
    2490 => 51,
    2491 => 51,
    2492 => 51,
    2493 => 51,
    2494 => 51,
    2495 => 51,
    2496 => 52,
    2497 => 52,
    2498 => 52,
    2499 => 52,
    2500 => 52,
    2501 => 52,
    2502 => 52,
    2503 => 52,
    2504 => 52,
    2505 => 52,
    2506 => 52,
    2507 => 52,
    2508 => 52,
    2509 => 52,
    2510 => 52,
    2511 => 52,
    2512 => 52,
    2513 => 52,
    2514 => 52,
    2515 => 52,
    2516 => 52,
    2517 => 52,
    2518 => 52,
    2519 => 52,
    2520 => 52,
    2521 => 52,
    2522 => 52,
    2523 => 52,
    2524 => 52,
    2525 => 52,
    2526 => 52,
    2527 => 52,
    2528 => 52,
    2529 => 52,
    2530 => 52,
    2531 => 52,
    2532 => 52,
    2533 => 52,
    2534 => 52,
    2535 => 52,
    2536 => 52,
    2537 => 52,
    2538 => 52,
    2539 => 52,
    2540 => 52,
    2541 => 52,
    2542 => 52,
    2543 => 52,
    2544 => 52,
    2545 => 52,
    2546 => 52,
    2547 => 52,
    2548 => 52,
    2549 => 52,
    2550 => 52,
    2551 => 52,
    2552 => 52,
    2553 => 52,
    2554 => 52,
    2555 => 52,
    2556 => 52,
    2557 => 52,
    2558 => 52,
    2559 => 52,
    2560 => 52,
    2561 => 52,
    2562 => 52,
    2563 => 52,
    2564 => 52,
    2565 => 52,
    2566 => 52,
    2567 => 52,
    2568 => 52,
    2569 => 53,
    2570 => 53,
    2571 => 53,
    2572 => 53,
    2573 => 53,
    2574 => 53,
    2575 => 53,
    2576 => 53,
    2577 => 53,
    2578 => 53,
    2579 => 53,
    2580 => 53,
    2581 => 53,
    2582 => 53,
    2583 => 53,
    2584 => 53,
    2585 => 53,
    2586 => 53,
    2587 => 53,
    2588 => 53,
    2589 => 53,
    2590 => 53,
    2591 => 53,
    2592 => 53,
    2593 => 53,
    2594 => 53,
    2595 => 53,
    2596 => 53,
    2597 => 53,
    2598 => 53,
    2599 => 53,
    2600 => 53,
    2601 => 53,
    2602 => 53,
    2603 => 53,
    2604 => 53,
    2605 => 53,
    2606 => 53,
    2607 => 53,
    2608 => 53,
    2609 => 53,
    2610 => 53,
    2611 => 53,
    2612 => 53,
    2613 => 53,
    2614 => 53,
    2615 => 53,
    2616 => 53,
    2617 => 53,
    2618 => 53,
    2619 => 53,
    2620 => 53,
    2621 => 53,
    2622 => 53,
    2623 => 53,
    2624 => 53,
    2625 => 53,
    2626 => 53,
    2627 => 53,
    2628 => 53,
    2629 => 53,
    2630 => 53,
    2631 => 53,
    2632 => 53,
    2633 => 53,
    2634 => 53,
    2635 => 53,
    2636 => 53,
    2637 => 53,
    2638 => 53,
    2639 => 53,
    2640 => 53,
    2641 => 53,
    2642 => 53,
    2643 => 53,
    2644 => 53,
    2645 => 53,
    2646 => 54,
    2647 => 54,
    2648 => 54,
    2649 => 54,
    2650 => 54,
    2651 => 54,
    2652 => 54,
    2653 => 54,
    2654 => 54,
    2655 => 54,
    2656 => 54,
    2657 => 54,
    2658 => 54,
    2659 => 54,
    2660 => 54,
    2661 => 54,
    2662 => 54,
    2663 => 54,
    2664 => 54,
    2665 => 54,
    2666 => 54,
    2667 => 54,
    2668 => 54,
    2669 => 54,
    2670 => 54,
    2671 => 54,
    2672 => 54,
    2673 => 54,
    2674 => 54,
    2675 => 54,
    2676 => 54,
    2677 => 54,
    2678 => 54,
    2679 => 54,
    2680 => 54,
    2681 => 54,
    2682 => 54,
    2683 => 54,
    2684 => 54,
    2685 => 54,
    2686 => 54,
    2687 => 54,
    2688 => 54,
    2689 => 54,
    2690 => 54,
    2691 => 54,
    2692 => 54,
    2693 => 54,
    2694 => 54,
    2695 => 54,
    2696 => 54,
    2697 => 54,
    2698 => 54,
    2699 => 54,
    2700 => 54,
    2701 => 54,
    2702 => 54,
    2703 => 54,
    2704 => 54,
    2705 => 54,
    2706 => 54,
    2707 => 54,
    2708 => 54,
    2709 => 54,
    2710 => 54,
    2711 => 54,
    2712 => 54,
    2713 => 54,
    2714 => 54,
    2715 => 54,
    2716 => 54,
    2717 => 54,
    2718 => 54,
    2719 => 54,
    2720 => 54,
    2721 => 54,
    2722 => 54,
    2723 => 54,
    2724 => 54,
    2725 => 54,
    2726 => 55,
    2727 => 55,
    2728 => 55,
    2729 => 55,
    2730 => 55,
    2731 => 55,
    2732 => 55,
    2733 => 55,
    2734 => 55,
    2735 => 55,
    2736 => 55,
    2737 => 55,
    2738 => 55,
    2739 => 55,
    2740 => 55,
    2741 => 55,
    2742 => 55,
    2743 => 55,
    2744 => 55,
    2745 => 55,
    2746 => 55,
    2747 => 55,
    2748 => 55,
    2749 => 55,
    2750 => 55,
    2751 => 55,
    2752 => 55,
    2753 => 55,
    2754 => 55,
    2755 => 55,
    2756 => 55,
    2757 => 55,
    2758 => 55,
    2759 => 55,
    2760 => 55,
    2761 => 55,
    2762 => 55,
    2763 => 55,
    2764 => 55,
    2765 => 55,
    2766 => 55,
    2767 => 55,
    2768 => 55,
    2769 => 55,
    2770 => 55,
    2771 => 55,
    2772 => 55,
    2773 => 55,
    2774 => 55,
    2775 => 55,
    2776 => 55,
    2777 => 55,
    2778 => 55,
    2779 => 55,
    2780 => 55,
    2781 => 55,
    2782 => 55,
    2783 => 55,
    2784 => 55,
    2785 => 55,
    2786 => 55,
    2787 => 55,
    2788 => 55,
    2789 => 55,
    2790 => 55,
    2791 => 55,
    2792 => 55,
    2793 => 55,
    2794 => 55,
    2795 => 55,
    2796 => 55,
    2797 => 55,
    2798 => 55,
    2799 => 55,
    2800 => 55,
    2801 => 55,
    2802 => 55,
    2803 => 55,
    2804 => 55,
    2805 => 55,
    2806 => 55,
    2807 => 55,
    2808 => 55,
    2809 => 55,
    2810 => 55,
    2811 => 56,
    2812 => 56,
    2813 => 56,
    2814 => 56,
    2815 => 56,
    2816 => 56,
    2817 => 56,
    2818 => 56,
    2819 => 56,
    2820 => 56,
    2821 => 56,
    2822 => 56,
    2823 => 56,
    2824 => 56,
    2825 => 56,
    2826 => 56,
    2827 => 56,
    2828 => 56,
    2829 => 56,
    2830 => 56,
    2831 => 56,
    2832 => 56,
    2833 => 56,
    2834 => 56,
    2835 => 56,
    2836 => 56,
    2837 => 56,
    2838 => 56,
    2839 => 56,
    2840 => 56,
    2841 => 56,
    2842 => 56,
    2843 => 56,
    2844 => 56,
    2845 => 56,
    2846 => 56,
    2847 => 56,
    2848 => 56,
    2849 => 56,
    2850 => 56,
    2851 => 56,
    2852 => 56,
    2853 => 56,
    2854 => 56,
    2855 => 56,
    2856 => 56,
    2857 => 56,
    2858 => 56,
    2859 => 56,
    2860 => 56,
    2861 => 56,
    2862 => 56,
    2863 => 56,
    2864 => 56,
    2865 => 56,
    2866 => 56,
    2867 => 56,
    2868 => 56,
    2869 => 56,
    2870 => 56,
    2871 => 56,
    2872 => 56,
    2873 => 56,
    2874 => 56,
    2875 => 56,
    2876 => 56,
    2877 => 56,
    2878 => 56,
    2879 => 56,
    2880 => 56,
    2881 => 56,
    2882 => 56,
    2883 => 56,
    2884 => 56,
    2885 => 56,
    2886 => 56,
    2887 => 56,
    2888 => 56,
    2889 => 56,
    2890 => 56,
    2891 => 56,
    2892 => 56,
    2893 => 56,
    2894 => 56,
    2895 => 56,
    2896 => 56,
    2897 => 56,
    2898 => 56,
    2899 => 56,
    2900 => 56,
    2901 => 56,
    2902 => 57,
    2903 => 57,
    2904 => 57,
    2905 => 57,
    2906 => 57,
    2907 => 57,
    2908 => 57,
    2909 => 57,
    2910 => 57,
    2911 => 57,
    2912 => 57,
    2913 => 57,
    2914 => 57,
    2915 => 57,
    2916 => 57,
    2917 => 57,
    2918 => 57,
    2919 => 57,
    2920 => 57,
    2921 => 57,
    2922 => 57,
    2923 => 57,
    2924 => 57,
    2925 => 57,
    2926 => 57,
    2927 => 57,
    2928 => 57,
    2929 => 57,
    2930 => 57,
    2931 => 57,
    2932 => 57,
    2933 => 57,
    2934 => 57,
    2935 => 57,
    2936 => 57,
    2937 => 57,
    2938 => 57,
    2939 => 57,
    2940 => 57,
    2941 => 57,
    2942 => 57,
    2943 => 57,
    2944 => 57,
    2945 => 57,
    2946 => 57,
    2947 => 57,
    2948 => 57,
    2949 => 57,
    2950 => 57,
    2951 => 57,
    2952 => 57,
    2953 => 57,
    2954 => 57,
    2955 => 57,
    2956 => 57,
    2957 => 57,
    2958 => 57,
    2959 => 57,
    2960 => 57,
    2961 => 57,
    2962 => 57,
    2963 => 57,
    2964 => 57,
    2965 => 57,
    2966 => 57,
    2967 => 57,
    2968 => 57,
    2969 => 57,
    2970 => 57,
    2971 => 57,
    2972 => 57,
    2973 => 57,
    2974 => 57,
    2975 => 57,
    2976 => 57,
    2977 => 57,
    2978 => 57,
    2979 => 57,
    2980 => 57,
    2981 => 57,
    2982 => 57,
    2983 => 57,
    2984 => 57,
    2985 => 57,
    2986 => 57,
    2987 => 57,
    2988 => 57,
    2989 => 57,
    2990 => 57,
    2991 => 57,
    2992 => 57,
    2993 => 57,
    2994 => 57,
    2995 => 57,
    2996 => 57,
    2997 => 57,
    2998 => 57,
    2999 => 58,
    3000 => 58,
    3001 => 58,
    3002 => 58,
    3003 => 58,
    3004 => 58,
    3005 => 58,
    3006 => 58,
    3007 => 58,
    3008 => 58,
    3009 => 58,
    3010 => 58,
    3011 => 58,
    3012 => 58,
    3013 => 58,
    3014 => 58,
    3015 => 58,
    3016 => 58,
    3017 => 58,
    3018 => 58,
    3019 => 58,
    3020 => 58,
    3021 => 58,
    3022 => 58,
    3023 => 58,
    3024 => 58,
    3025 => 58,
    3026 => 58,
    3027 => 58,
    3028 => 58,
    3029 => 58,
    3030 => 58,
    3031 => 58,
    3032 => 58,
    3033 => 58,
    3034 => 58,
    3035 => 58,
    3036 => 58,
    3037 => 58,
    3038 => 58,
    3039 => 58,
    3040 => 58,
    3041 => 58,
    3042 => 58,
    3043 => 58,
    3044 => 58,
    3045 => 58,
    3046 => 58,
    3047 => 58,
    3048 => 58,
    3049 => 58,
    3050 => 58,
    3051 => 58,
    3052 => 58,
    3053 => 58,
    3054 => 58,
    3055 => 58,
    3056 => 58,
    3057 => 58,
    3058 => 58,
    3059 => 58,
    3060 => 58,
    3061 => 58,
    3062 => 58,
    3063 => 58,
    3064 => 58,
    3065 => 58,
    3066 => 58,
    3067 => 58,
    3068 => 58,
    3069 => 58,
    3070 => 58,
    3071 => 58,
    3072 => 58,
    3073 => 58,
    3074 => 58,
    3075 => 58,
    3076 => 58,
    3077 => 58,
    3078 => 58,
    3079 => 58,
    3080 => 58,
    3081 => 58,
    3082 => 58,
    3083 => 58,
    3084 => 58,
    3085 => 58,
    3086 => 58,
    3087 => 58,
    3088 => 58,
    3089 => 58,
    3090 => 58,
    3091 => 58,
    3092 => 58,
    3093 => 58,
    3094 => 58,
    3095 => 58,
    3096 => 58,
    3097 => 58,
    3098 => 58,
    3099 => 58,
    3100 => 58,
    3101 => 58,
    3102 => 58,
    3103 => 58,
    3104 => 58,
    3105 => 59,
    3106 => 59,
    3107 => 59,
    3108 => 59,
    3109 => 59,
    3110 => 59,
    3111 => 59,
    3112 => 59,
    3113 => 59,
    3114 => 59,
    3115 => 59,
    3116 => 59,
    3117 => 59,
    3118 => 59,
    3119 => 59,
    3120 => 59,
    3121 => 59,
    3122 => 59,
    3123 => 59,
    3124 => 59,
    3125 => 59,
    3126 => 59,
    3127 => 59,
    3128 => 59,
    3129 => 59,
    3130 => 59,
    3131 => 59,
    3132 => 59,
    3133 => 59,
    3134 => 59,
    3135 => 59,
    3136 => 59,
    3137 => 59,
    3138 => 59,
    3139 => 59,
    3140 => 59,
    3141 => 59,
    3142 => 59,
    3143 => 59,
    3144 => 59,
    3145 => 59,
    3146 => 59,
    3147 => 59,
    3148 => 59,
    3149 => 59,
    3150 => 59,
    3151 => 59,
    3152 => 59,
    3153 => 59,
    3154 => 59,
    3155 => 59,
    3156 => 59,
    3157 => 59,
    3158 => 59,
    3159 => 59,
    3160 => 59,
    3161 => 59,
    3162 => 59,
    3163 => 59,
    3164 => 59,
    3165 => 59,
    3166 => 59,
    3167 => 59,
    3168 => 59,
    3169 => 59,
    3170 => 59,
    3171 => 59,
    3172 => 59,
    3173 => 59,
    3174 => 59,
    3175 => 59,
    3176 => 59,
    3177 => 59,
    3178 => 59,
    3179 => 59,
    3180 => 59,
    3181 => 59,
    3182 => 59,
    3183 => 59,
    3184 => 59,
    3185 => 59,
    3186 => 59,
    3187 => 59,
    3188 => 59,
    3189 => 59,
    3190 => 59,
    3191 => 59,
    3192 => 59,
    3193 => 59,
    3194 => 59,
    3195 => 59,
    3196 => 59,
    3197 => 59,
    3198 => 59,
    3199 => 59,
    3200 => 59,
    3201 => 59,
    3202 => 59,
    3203 => 59,
    3204 => 59,
    3205 => 59,
    3206 => 59,
    3207 => 59,
    3208 => 59,
    3209 => 59,
    3210 => 59,
    3211 => 59,
    3212 => 59,
    3213 => 59,
    3214 => 59,
    3215 => 59,
    3216 => 59,
    3217 => 59,
    3218 => 59,
    3219 => 59,
    3220 => 59,
    3221 => 59,
    3222 => 59,
    3223 => 60,
    3224 => 60,
    3225 => 60,
    3226 => 60,
    3227 => 60,
    3228 => 60,
    3229 => 60,
    3230 => 60,
    3231 => 60,
    3232 => 60,
    3233 => 60,
    3234 => 60,
    3235 => 60,
    3236 => 60,
    3237 => 60,
    3238 => 60,
    3239 => 60,
    3240 => 60,
    3241 => 60,
    3242 => 60,
    3243 => 60,
    3244 => 60,
    3245 => 60,
    3246 => 60,
    3247 => 60,
    3248 => 60,
    3249 => 60,
    3250 => 60,
    3251 => 60,
    3252 => 60,
    3253 => 60,
    3254 => 60,
    3255 => 60,
    3256 => 60,
    3257 => 60,
    3258 => 60,
    3259 => 60,
    3260 => 60,
    3261 => 60,
    3262 => 60,
    3263 => 60,
    3264 => 60,
    3265 => 60,
    3266 => 60,
    3267 => 60,
    3268 => 60,
    3269 => 60,
    3270 => 60,
    3271 => 60,
    3272 => 60,
    3273 => 60,
    3274 => 60,
    3275 => 60,
    3276 => 60,
    3277 => 60,
    3278 => 60,
    3279 => 60,
    3280 => 60,
    3281 => 60,
    3282 => 60,
    3283 => 60,
    3284 => 60,
    3285 => 60,
    3286 => 60,
    3287 => 60,
    3288 => 60,
    3289 => 60,
    3290 => 60,
    3291 => 60,
    3292 => 60,
    3293 => 60,
    3294 => 60,
    3295 => 60,
    3296 => 60,
    3297 => 60,
    3298 => 60,
    3299 => 60,
    3300 => 60,
    3301 => 60,
    3302 => 60,
    3303 => 60,
    3304 => 60,
    3305 => 60,
    3306 => 60,
    3307 => 60,
    3308 => 60,
    3309 => 60,
    3310 => 60,
    3311 => 60,
    3312 => 60,
    3313 => 60,
    3314 => 60,
    3315 => 60,
    3316 => 60,
    3317 => 60,
    3318 => 60,
    3319 => 60,
    3320 => 60,
    3321 => 60,
    3322 => 60,
    3323 => 60,
    3324 => 60,
    3325 => 60,
    3326 => 60,
    3327 => 60,
    3328 => 60,
    3329 => 60,
    3330 => 60,
    3331 => 60,
    3332 => 60,
    3333 => 60,
    3334 => 60,
    3335 => 60,
    3336 => 60,
    3337 => 60,
    3338 => 60,
    3339 => 60,
    3340 => 60,
    3341 => 60,
    3342 => 60,
    3343 => 60,
    3344 => 60,
    3345 => 60,
    3346 => 60,
    3347 => 60,
    3348 => 60,
    3349 => 60,
    3350 => 60,
    3351 => 60,
    3352 => 60,
    3353 => 60,
    3354 => 60,
    3355 => 60,
    3356 => 60,
    3357 => 60,
    3358 => 60,
    3359 => 61,
    3360 => 61,
    3361 => 61,
    3362 => 61,
    3363 => 61,
    3364 => 61,
    3365 => 61,
    3366 => 61,
    3367 => 61,
    3368 => 61,
    3369 => 61,
    3370 => 61,
    3371 => 61,
    3372 => 61,
    3373 => 61,
    3374 => 61,
    3375 => 61,
    3376 => 61,
    3377 => 61,
    3378 => 61,
    3379 => 61,
    3380 => 61,
    3381 => 61,
    3382 => 61,
    3383 => 61,
    3384 => 61,
    3385 => 61,
    3386 => 61,
    3387 => 61,
    3388 => 61,
    3389 => 61,
    3390 => 61,
    3391 => 61,
    3392 => 61,
    3393 => 61,
    3394 => 61,
    3395 => 61,
    3396 => 61,
    3397 => 61,
    3398 => 61,
    3399 => 61,
    3400 => 61,
    3401 => 61,
    3402 => 61,
    3403 => 61,
    3404 => 61,
    3405 => 61,
    3406 => 61,
    3407 => 61,
    3408 => 61,
    3409 => 61,
    3410 => 61,
    3411 => 61,
    3412 => 61,
    3413 => 61,
    3414 => 61,
    3415 => 61,
    3416 => 61,
    3417 => 61,
    3418 => 61,
    3419 => 61,
    3420 => 61,
    3421 => 61,
    3422 => 61,
    3423 => 61,
    3424 => 61,
    3425 => 61,
    3426 => 61,
    3427 => 61,
    3428 => 61,
    3429 => 61,
    3430 => 61,
    3431 => 61,
    3432 => 61,
    3433 => 61,
    3434 => 61,
    3435 => 61,
    3436 => 61,
    3437 => 61,
    3438 => 61,
    3439 => 61,
    3440 => 61,
    3441 => 61,
    3442 => 61,
    3443 => 61,
    3444 => 61,
    3445 => 61,
    3446 => 61,
    3447 => 61,
    3448 => 61,
    3449 => 61,
    3450 => 61,
    3451 => 61,
    3452 => 61,
    3453 => 61,
    3454 => 61,
    3455 => 61,
    3456 => 61,
    3457 => 61,
    3458 => 61,
    3459 => 61,
    3460 => 61,
    3461 => 61,
    3462 => 61,
    3463 => 61,
    3464 => 61,
    3465 => 61,
    3466 => 61,
    3467 => 61,
    3468 => 61,
    3469 => 61,
    3470 => 61,
    3471 => 61,
    3472 => 61,
    3473 => 61,
    3474 => 61,
    3475 => 61,
    3476 => 61,
    3477 => 61,
    3478 => 61,
    3479 => 61,
    3480 => 61,
    3481 => 61,
    3482 => 61,
    3483 => 61,
    3484 => 61,
    3485 => 61,
    3486 => 61,
    3487 => 61,
    3488 => 61,
    3489 => 61,
    3490 => 61,
    3491 => 61,
    3492 => 61,
    3493 => 61,
    3494 => 61,
    3495 => 61,
    3496 => 61,
    3497 => 61,
    3498 => 61,
    3499 => 61,
    3500 => 61,
    3501 => 61,
    3502 => 61,
    3503 => 61,
    3504 => 61,
    3505 => 61,
    3506 => 61,
    3507 => 61,
    3508 => 61,
    3509 => 61,
    3510 => 61,
    3511 => 61,
    3512 => 61,
    3513 => 61,
    3514 => 61,
    3515 => 61,
    3516 => 61,
    3517 => 61,
    3518 => 61,
    3519 => 61,
    3520 => 61,
    3521 => 61,
    3522 => 61,
    3523 => 61,
    3524 => 61,
    3525 => 61,
    3526 => 62,
    3527 => 62,
    3528 => 62,
    3529 => 62,
    3530 => 62,
    3531 => 62,
    3532 => 62,
    3533 => 62,
    3534 => 62,
    3535 => 62,
    3536 => 62,
    3537 => 62,
    3538 => 62,
    3539 => 62,
    3540 => 62,
    3541 => 62,
    3542 => 62,
    3543 => 62,
    3544 => 62,
    3545 => 62,
    3546 => 62,
    3547 => 62,
    3548 => 62,
    3549 => 62,
    3550 => 62,
    3551 => 62,
    3552 => 62,
    3553 => 62,
    3554 => 62,
    3555 => 62,
    3556 => 62,
    3557 => 62,
    3558 => 62,
    3559 => 62,
    3560 => 62,
    3561 => 62,
    3562 => 62,
    3563 => 62,
    3564 => 62,
    3565 => 62,
    3566 => 62,
    3567 => 62,
    3568 => 62,
    3569 => 62,
    3570 => 62,
    3571 => 62,
    3572 => 62,
    3573 => 62,
    3574 => 62,
    3575 => 62,
    3576 => 62,
    3577 => 62,
    3578 => 62,
    3579 => 62,
    3580 => 62,
    3581 => 62,
    3582 => 62,
    3583 => 62,
    3584 => 62,
    3585 => 62,
    3586 => 62,
    3587 => 62,
    3588 => 62,
    3589 => 62,
    3590 => 62,
    3591 => 62,
    3592 => 62,
    3593 => 62,
    3594 => 62,
    3595 => 62,
    3596 => 62,
    3597 => 62,
    3598 => 62,
    3599 => 62,
    3600 => 62,
    3601 => 62,
    3602 => 62,
    3603 => 62,
    3604 => 62,
    3605 => 62,
    3606 => 62,
    3607 => 62,
    3608 => 62,
    3609 => 62,
    3610 => 62,
    3611 => 62,
    3612 => 62,
    3613 => 62,
    3614 => 62,
    3615 => 62,
    3616 => 62,
    3617 => 62,
    3618 => 62,
    3619 => 62,
    3620 => 62,
    3621 => 62,
    3622 => 62,
    3623 => 62,
    3624 => 62,
    3625 => 62,
    3626 => 62,
    3627 => 62,
    3628 => 62,
    3629 => 62,
    3630 => 62,
    3631 => 62,
    3632 => 62,
    3633 => 62,
    3634 => 62,
    3635 => 62,
    3636 => 62,
    3637 => 62,
    3638 => 62,
    3639 => 62,
    3640 => 62,
    3641 => 62,
    3642 => 62,
    3643 => 62,
    3644 => 62,
    3645 => 62,
    3646 => 62,
    3647 => 62,
    3648 => 62,
    3649 => 62,
    3650 => 62,
    3651 => 62,
    3652 => 62,
    3653 => 62,
    3654 => 62,
    3655 => 62,
    3656 => 62,
    3657 => 62,
    3658 => 62,
    3659 => 62,
    3660 => 62,
    3661 => 62,
    3662 => 62,
    3663 => 62,
    3664 => 62,
    3665 => 62,
    3666 => 62,
    3667 => 62,
    3668 => 62,
    3669 => 62,
    3670 => 62,
    3671 => 62,
    3672 => 62,
    3673 => 62,
    3674 => 62,
    3675 => 62,
    3676 => 62,
    3677 => 62,
    3678 => 62,
    3679 => 62,
    3680 => 62,
    3681 => 62,
    3682 => 62,
    3683 => 62,
    3684 => 62,
    3685 => 62,
    3686 => 62,
    3687 => 62,
    3688 => 62,
    3689 => 62,
    3690 => 62,
    3691 => 62,
    3692 => 62,
    3693 => 62,
    3694 => 62,
    3695 => 62,
    3696 => 62,
    3697 => 62,
    3698 => 62,
    3699 => 62,
    3700 => 62,
    3701 => 62,
    3702 => 62,
    3703 => 62,
    3704 => 62,
    3705 => 62,
    3706 => 62,
    3707 => 62,
    3708 => 62,
    3709 => 62,
    3710 => 62,
    3711 => 62,
    3712 => 62,
    3713 => 62,
    3714 => 62,
    3715 => 62,
    3716 => 62,
    3717 => 62,
    3718 => 62,
    3719 => 62,
    3720 => 62,
    3721 => 62,
    3722 => 62,
    3723 => 62,
    3724 => 62,
    3725 => 62,
    3726 => 62,
    3727 => 62,
    3728 => 62,
    3729 => 62,
    3730 => 62,
    3731 => 62,
    3732 => 62,
    3733 => 62,
    3734 => 62,
    3735 => 62,
    3736 => 62,
    3737 => 62,
    3738 => 62,
    3739 => 62,
    3740 => 62,
    3741 => 62,
    3742 => 62,
    3743 => 62,
    3744 => 62,
    3745 => 62,
    3746 => 62,
    3747 => 62,
    3748 => 62,
    3749 => 62,
    3750 => 62,
    3751 => 62,
    3752 => 62,
    3753 => 62,
    3754 => 62,
    3755 => 62,
    3756 => 62,
    3757 => 62,
    3758 => 62,
    3759 => 62,
    3760 => 62,
    3761 => 62,
    3762 => 62,
    3763 => 62,
    3764 => 62,
    3765 => 62,
    3766 => 62,
    3767 => 62,
    3768 => 63,
    3769 => 63,
    3770 => 63,
    3771 => 63,
    3772 => 63,
    3773 => 63,
    3774 => 63,
    3775 => 63,
    3776 => 63,
    3777 => 63,
    3778 => 63,
    3779 => 63,
    3780 => 63,
    3781 => 63,
    3782 => 63,
    3783 => 63,
    3784 => 63,
    3785 => 63,
    3786 => 63,
    3787 => 63,
    3788 => 63,
    3789 => 63,
    3790 => 63,
    3791 => 63,
    3792 => 63,
    3793 => 63,
    3794 => 63,
    3795 => 63,
    3796 => 63,
    3797 => 63,
    3798 => 63,
    3799 => 63,
    3800 => 63,
    3801 => 63,
    3802 => 63,
    3803 => 63,
    3804 => 63,
    3805 => 63,
    3806 => 63,
    3807 => 63,
    3808 => 63,
    3809 => 63,
    3810 => 63,
    3811 => 63,
    3812 => 63,
    3813 => 63,
    3814 => 63,
    3815 => 63,
    3816 => 63,
    3817 => 63,
    3818 => 63,
    3819 => 63,
    3820 => 63,
    3821 => 63,
    3822 => 63,
    3823 => 63,
    3824 => 63,
    3825 => 63,
    3826 => 63,
    3827 => 63,
    3828 => 63,
    3829 => 63,
    3830 => 63,
    3831 => 63,
    3832 => 63,
    3833 => 63,
    3834 => 63,
    3835 => 63,
    3836 => 63,
    3837 => 63,
    3838 => 63,
    3839 => 63,
    3840 => 63,
    3841 => 63,
    3842 => 63,
    3843 => 63,
    3844 => 63,
    3845 => 63,
    3846 => 63,
    3847 => 63,
    3848 => 63,
    3849 => 63,
    3850 => 63,
    3851 => 63,
    3852 => 63,
    3853 => 63,
    3854 => 63,
    3855 => 63,
    3856 => 63,
    3857 => 63,
    3858 => 63,
    3859 => 63,
    3860 => 63,
    3861 => 63,
    3862 => 63,
    3863 => 63,
    3864 => 63,
    3865 => 63,
    3866 => 63,
    3867 => 63,
    3868 => 63,
    3869 => 63,
    3870 => 63,
    3871 => 63,
    3872 => 63,
    3873 => 63,
    3874 => 63,
    3875 => 63,
    3876 => 63,
    3877 => 63,
    3878 => 63,
    3879 => 63,
    3880 => 63,
    3881 => 63,
    3882 => 63,
    3883 => 63,
    3884 => 63,
    3885 => 63,
    3886 => 63,
    3887 => 63,
    3888 => 63,
    3889 => 63,
    3890 => 63,
    3891 => 63,
    3892 => 63,
    3893 => 63,
    3894 => 63,
    3895 => 63,
    3896 => 63,
    3897 => 63,
    3898 => 63,
    3899 => 63,
    3900 => 63,
    3901 => 63,
    3902 => 63,
    3903 => 63,
    3904 => 63,
    3905 => 63,
    3906 => 63,
    3907 => 63,
    3908 => 63,
    3909 => 63,
    3910 => 63,
    3911 => 63,
    3912 => 63,
    3913 => 63,
    3914 => 63,
    3915 => 63,
    3916 => 63,
    3917 => 63,
    3918 => 63,
    3919 => 63,
    3920 => 63,
    3921 => 63,
    3922 => 63,
    3923 => 63,
    3924 => 63,
    3925 => 63,
    3926 => 63,
    3927 => 63,
    3928 => 63,
    3929 => 63,
    3930 => 63,
    3931 => 63,
    3932 => 63,
    3933 => 63,
    3934 => 63,
    3935 => 63,
    3936 => 63,
    3937 => 63,
    3938 => 63,
    3939 => 63,
    3940 => 63,
    3941 => 63,
    3942 => 63,
    3943 => 63,
    3944 => 63,
    3945 => 63,
    3946 => 63,
    3947 => 63,
    3948 => 63,
    3949 => 63,
    3950 => 63,
    3951 => 63,
    3952 => 63,
    3953 => 63,
    3954 => 63,
    3955 => 63,
    3956 => 63,
    3957 => 63,
    3958 => 63,
    3959 => 63,
    3960 => 63,
    3961 => 63,
    3962 => 63,
    3963 => 63,
    3964 => 63,
    3965 => 63,
    3966 => 63,
    3967 => 63,
    3968 => 63,
    3969 => 63,
    3970 => 63,
    3971 => 63,
    3972 => 63,
    3973 => 63,
    3974 => 63,
    3975 => 63,
    3976 => 63,
    3977 => 63,
    3978 => 63,
    3979 => 63,
    3980 => 63,
    3981 => 63,
    3982 => 63,
    3983 => 63,
    3984 => 63,
    3985 => 63,
    3986 => 63,
    3987 => 63,
    3988 => 63,
    3989 => 63,
    3990 => 63,
    3991 => 63,
    3992 => 63,
    3993 => 63,
    3994 => 63,
    3995 => 63,
    3996 => 63,
    3997 => 63,
    3998 => 63,
    3999 => 63,
    4000 => 63,
    4001 => 63,
    4002 => 63,
    4003 => 63,
    4004 => 63,
    4005 => 63,
    4006 => 63,
    4007 => 63,
    4008 => 63,
    4009 => 63,
    4010 => 63,
    4011 => 63,
    4012 => 63,
    4013 => 63,
    4014 => 63,
    4015 => 63,
    4016 => 63,
    4017 => 63,
    4018 => 63,
    4019 => 63,
    4020 => 63,
    4021 => 63,
    4022 => 63,
    4023 => 63,
    4024 => 63,
    4025 => 63,
    4026 => 63,
    4027 => 63,
    4028 => 63,
    4029 => 63,
    4030 => 63,
    4031 => 63,
    4032 => 63,
    4033 => 63,
    4034 => 63,
    4035 => 63,
    4036 => 63,
    4037 => 63,
    4038 => 63,
    4039 => 63,
    4040 => 63,
    4041 => 63,
    4042 => 63,
    4043 => 63,
    4044 => 63,
    4045 => 63,
    4046 => 63,
    4047 => 63,
    4048 => 63,
    4049 => 63,
    4050 => 63,
    4051 => 63,
    4052 => 63,
    4053 => 63,
    4054 => 63,
    4055 => 63,
    4056 => 63,
    4057 => 63,
    4058 => 63,
    4059 => 63,
    4060 => 63,
    4061 => 63,
    4062 => 63,
    4063 => 63,
    4064 => 63,
    4065 => 63,
    4066 => 63,
    4067 => 63,
    4068 => 63,
    4069 => 63,
    4070 => 63,
    4071 => 63,
    4072 => 63,
    4073 => 63,
    4074 => 63,
    4075 => 63,
    4076 => 63,
    4077 => 63,
    4078 => 63,
    4079 => 63,
    4080 => 63,
    4081 => 63,
    4082 => 63,
    4083 => 63,
    4084 => 63,
    4085 => 63,
    4086 => 63,
    4087 => 63,
    4088 => 63,
    4089 => 63,
    4090 => 63,
    4091 => 63,
    4092 => 63,
    4093 => 63,
    4094 => 63,
    4095 => 63,
    4096 => 63,
    4097 => 63,
    4098 => 63,
    4099 => 63,
    4100 => 63,
    4101 => 63,
    4102 => 63,
    4103 => 63,
    4104 => 63,
    4105 => 63,
    4106 => 63,
    4107 => 63,
    4108 => 63,
    4109 => 63,
    4110 => 63,
    4111 => 63,
    4112 => 63,
    4113 => 63,
    4114 => 63,
    4115 => 63,
    4116 => 63,
    4117 => 63,
    4118 => 63,
    4119 => 63,
    4120 => 63,
    4121 => 63,
    4122 => 63,
    4123 => 63,
    4124 => 63,
    4125 => 63,
    4126 => 63,
    4127 => 63,
    4128 => 63,
    4129 => 63,
    4130 => 63,
    4131 => 63,
    4132 => 63,
    4133 => 63,
    4134 => 63,
    4135 => 63,
    4136 => 63,
    4137 => 63,
    4138 => 63,
    4139 => 63,
    4140 => 63,
    4141 => 63,
    4142 => 63,
    4143 => 63,
    4144 => 63,
    4145 => 63,
    4146 => 63,
    4147 => 63,
    4148 => 63,
    4149 => 63,
    4150 => 63,
    4151 => 63,
    4152 => 63,
    4153 => 63,
    4154 => 63,
    4155 => 63,
    4156 => 63,
    4157 => 63,
    4158 => 63,
    4159 => 63,
    4160 => 63,
    4161 => 63,
    4162 => 63,
    4163 => 63,
    4164 => 63,
    4165 => 63,
    4166 => 63,
    4167 => 63,
    4168 => 63,
    4169 => 63,
    4170 => 63,
    4171 => 63,
    4172 => 63,
    4173 => 63,
    4174 => 63,
    4175 => 63,
    4176 => 63,
    4177 => 63,
    4178 => 63,
    4179 => 63,
    4180 => 63,
    4181 => 63,
    4182 => 63,
    4183 => 63,
    4184 => 63,
    4185 => 63,
    4186 => 63,
    4187 => 63,
    4188 => 63,
    4189 => 63,
    4190 => 63,
    4191 => 63,
    4192 => 63,
    4193 => 63,
    4194 => 63,
    4195 => 63,
    4196 => 63,
    4197 => 63,
    4198 => 63,
    4199 => 63,
    4200 => 63,
    4201 => 63,
    4202 => 63,
    4203 => 63,
    4204 => 63,
    4205 => 63,
    4206 => 63,
    4207 => 63,
    4208 => 63,
    4209 => 63,
    4210 => 63,
    4211 => 63,
    4212 => 63,
    4213 => 63,
    4214 => 63,
    4215 => 63,
    4216 => 63,
    4217 => 63,
    4218 => 63,
    4219 => 63,
    4220 => 63,
    4221 => 63,
    4222 => 63,
    4223 => 63,
    4224 => 63,
    4225 => 63,
    4226 => 63,
    4227 => 63,
    4228 => 63,
    4229 => 63,
    4230 => 63,
    4231 => 63,
    4232 => 63,
    4233 => 63,
    4234 => 63,
    4235 => 63,
    4236 => 63,
    4237 => 63,
    4238 => 63,
    4239 => 63,
    4240 => 63,
    4241 => 63,
    4242 => 63,
    4243 => 63,
    4244 => 63,
    4245 => 63,
    4246 => 63,
    4247 => 63,
    4248 => 63,
    4249 => 63,
    4250 => 63,
    4251 => 63,
    4252 => 63,
    4253 => 63,
    4254 => 63,
    4255 => 63,
    4256 => 63,
    4257 => 63,
    4258 => 63,
    4259 => 63,
    4260 => 63,
    4261 => 63,
    4262 => 63,
    4263 => 63,
    4264 => 63,
    4265 => 63,
    4266 => 63,
    4267 => 63,
    4268 => 63,
    4269 => 63,
    4270 => 63,
    4271 => 63,
    4272 => 63,
    4273 => 63,
    4274 => 63,
    4275 => 63,
    4276 => 63,
    4277 => 63,
    4278 => 63,
    4279 => 63,
    4280 => 63,
    4281 => 63,
    4282 => 63,
    4283 => 63,
    4284 => 63,
    4285 => 63,
    4286 => 63,
    4287 => 63,
    4288 => 63,
    4289 => 63,
    4290 => 63,
    4291 => 63,
    4292 => 63,
    4293 => 63,
    4294 => 63,
    4295 => 63,
    4296 => 63,
    4297 => 63,
    4298 => 63,
    4299 => 63,
    4300 => 63,
    4301 => 63,
    4302 => 63,
    4303 => 63,
    4304 => 63,
    4305 => 63,
    4306 => 63,
    4307 => 63,
    4308 => 63,
    4309 => 63,
    4310 => 63,
    4311 => 63,
    4312 => 63,
    4313 => 63,
    4314 => 63,
    4315 => 63,
    4316 => 63,
    4317 => 63,
    4318 => 63,
    4319 => 63,
    4320 => 63,
    4321 => 63,
    4322 => 63,
    4323 => 63,
    4324 => 63,
    4325 => 63,
    4326 => 63,
    4327 => 63,
    4328 => 63,
    4329 => 63,
    4330 => 63,
    4331 => 63,
    4332 => 63,
    4333 => 63,
    4334 => 63,
    4335 => 63,
    4336 => 63,
    4337 => 63,
    4338 => 63,
    4339 => 63,
    4340 => 63,
    4341 => 63,
    4342 => 63,
    4343 => 63,
    4344 => 63,
    4345 => 63,
    4346 => 63,
    4347 => 63,
    4348 => 63,
    4349 => 63,
    4350 => 63,
    4351 => 63,
    4352 => 63,
    4353 => 63,
    4354 => 63,
    4355 => 63,
    4356 => 63,
    4357 => 63,
    4358 => 63,
    4359 => 63,
    4360 => 63,
    4361 => 63,
    4362 => 63,
    4363 => 63,
    4364 => 63,
    4365 => 63,
    4366 => 63,
    4367 => 63,
    4368 => 63,
    4369 => 63,
    4370 => 63,
    4371 => 63,
    4372 => 63,
    4373 => 63,
    4374 => 63,
    4375 => 63,
    4376 => 63,
    4377 => 63,
    4378 => 63,
    4379 => 63,
    4380 => 63,
    4381 => 63,
    4382 => 63,
    4383 => 63,
    4384 => 63,
    4385 => 63,
    4386 => 63,
    4387 => 63,
    4388 => 63,
    4389 => 63,
    4390 => 63,
    4391 => 63,
    4392 => 63,
    4393 => 63,
    4394 => 63,
    4395 => 63,
    4396 => 63,
    4397 => 63,
    4398 => 63,
    4399 => 63,
    4400 => 63,
    4401 => 63,
    4402 => 63,
    4403 => 63,
    4404 => 63,
    4405 => 63,
    4406 => 63,
    4407 => 63,
    4408 => 63,
    4409 => 63,
    4410 => 63,
    4411 => 63,
    4412 => 63,
    4413 => 63,
    4414 => 63,
    4415 => 63,
    4416 => 63,
    4417 => 63,
    4418 => 63,
    4419 => 63,
    4420 => 63,
    4421 => 63,
    4422 => 63,
    4423 => 63,
    4424 => 63,
    4425 => 62,
    4426 => 62,
    4427 => 62,
    4428 => 62,
    4429 => 62,
    4430 => 62,
    4431 => 62,
    4432 => 62,
    4433 => 62,
    4434 => 62,
    4435 => 62,
    4436 => 62,
    4437 => 62,
    4438 => 62,
    4439 => 62,
    4440 => 62,
    4441 => 62,
    4442 => 62,
    4443 => 62,
    4444 => 62,
    4445 => 62,
    4446 => 62,
    4447 => 62,
    4448 => 62,
    4449 => 62,
    4450 => 62,
    4451 => 62,
    4452 => 62,
    4453 => 62,
    4454 => 62,
    4455 => 62,
    4456 => 62,
    4457 => 62,
    4458 => 62,
    4459 => 62,
    4460 => 62,
    4461 => 62,
    4462 => 62,
    4463 => 62,
    4464 => 62,
    4465 => 62,
    4466 => 62,
    4467 => 62,
    4468 => 62,
    4469 => 62,
    4470 => 62,
    4471 => 62,
    4472 => 62,
    4473 => 62,
    4474 => 62,
    4475 => 62,
    4476 => 62,
    4477 => 62,
    4478 => 62,
    4479 => 62,
    4480 => 62,
    4481 => 62,
    4482 => 62,
    4483 => 62,
    4484 => 62,
    4485 => 62,
    4486 => 62,
    4487 => 62,
    4488 => 62,
    4489 => 62,
    4490 => 62,
    4491 => 62,
    4492 => 62,
    4493 => 62,
    4494 => 62,
    4495 => 62,
    4496 => 62,
    4497 => 62,
    4498 => 62,
    4499 => 62,
    4500 => 62,
    4501 => 62,
    4502 => 62,
    4503 => 62,
    4504 => 62,
    4505 => 62,
    4506 => 62,
    4507 => 62,
    4508 => 62,
    4509 => 62,
    4510 => 62,
    4511 => 62,
    4512 => 62,
    4513 => 62,
    4514 => 62,
    4515 => 62,
    4516 => 62,
    4517 => 62,
    4518 => 62,
    4519 => 62,
    4520 => 62,
    4521 => 62,
    4522 => 62,
    4523 => 62,
    4524 => 62,
    4525 => 62,
    4526 => 62,
    4527 => 62,
    4528 => 62,
    4529 => 62,
    4530 => 62,
    4531 => 62,
    4532 => 62,
    4533 => 62,
    4534 => 62,
    4535 => 62,
    4536 => 62,
    4537 => 62,
    4538 => 62,
    4539 => 62,
    4540 => 62,
    4541 => 62,
    4542 => 62,
    4543 => 62,
    4544 => 62,
    4545 => 62,
    4546 => 62,
    4547 => 62,
    4548 => 62,
    4549 => 62,
    4550 => 62,
    4551 => 62,
    4552 => 62,
    4553 => 62,
    4554 => 62,
    4555 => 62,
    4556 => 62,
    4557 => 62,
    4558 => 62,
    4559 => 62,
    4560 => 62,
    4561 => 62,
    4562 => 62,
    4563 => 62,
    4564 => 62,
    4565 => 62,
    4566 => 62,
    4567 => 62,
    4568 => 62,
    4569 => 62,
    4570 => 62,
    4571 => 62,
    4572 => 62,
    4573 => 62,
    4574 => 62,
    4575 => 62,
    4576 => 62,
    4577 => 62,
    4578 => 62,
    4579 => 62,
    4580 => 62,
    4581 => 62,
    4582 => 62,
    4583 => 62,
    4584 => 62,
    4585 => 62,
    4586 => 62,
    4587 => 62,
    4588 => 62,
    4589 => 62,
    4590 => 62,
    4591 => 62,
    4592 => 62,
    4593 => 62,
    4594 => 62,
    4595 => 62,
    4596 => 62,
    4597 => 62,
    4598 => 62,
    4599 => 62,
    4600 => 62,
    4601 => 62,
    4602 => 62,
    4603 => 62,
    4604 => 62,
    4605 => 62,
    4606 => 62,
    4607 => 62,
    4608 => 62,
    4609 => 62,
    4610 => 62,
    4611 => 62,
    4612 => 62,
    4613 => 62,
    4614 => 62,
    4615 => 62,
    4616 => 62,
    4617 => 62,
    4618 => 62,
    4619 => 62,
    4620 => 62,
    4621 => 62,
    4622 => 62,
    4623 => 62,
    4624 => 62,
    4625 => 62,
    4626 => 62,
    4627 => 62,
    4628 => 62,
    4629 => 62,
    4630 => 62,
    4631 => 62,
    4632 => 62,
    4633 => 62,
    4634 => 62,
    4635 => 62,
    4636 => 62,
    4637 => 62,
    4638 => 62,
    4639 => 62,
    4640 => 62,
    4641 => 62,
    4642 => 62,
    4643 => 62,
    4644 => 62,
    4645 => 62,
    4646 => 62,
    4647 => 62,
    4648 => 62,
    4649 => 62,
    4650 => 62,
    4651 => 62,
    4652 => 62,
    4653 => 62,
    4654 => 62,
    4655 => 62,
    4656 => 62,
    4657 => 62,
    4658 => 62,
    4659 => 62,
    4660 => 62,
    4661 => 62,
    4662 => 62,
    4663 => 62,
    4664 => 62,
    4665 => 62,
    4666 => 62,
    4667 => 61,
    4668 => 61,
    4669 => 61,
    4670 => 61,
    4671 => 61,
    4672 => 61,
    4673 => 61,
    4674 => 61,
    4675 => 61,
    4676 => 61,
    4677 => 61,
    4678 => 61,
    4679 => 61,
    4680 => 61,
    4681 => 61,
    4682 => 61,
    4683 => 61,
    4684 => 61,
    4685 => 61,
    4686 => 61,
    4687 => 61,
    4688 => 61,
    4689 => 61,
    4690 => 61,
    4691 => 61,
    4692 => 61,
    4693 => 61,
    4694 => 61,
    4695 => 61,
    4696 => 61,
    4697 => 61,
    4698 => 61,
    4699 => 61,
    4700 => 61,
    4701 => 61,
    4702 => 61,
    4703 => 61,
    4704 => 61,
    4705 => 61,
    4706 => 61,
    4707 => 61,
    4708 => 61,
    4709 => 61,
    4710 => 61,
    4711 => 61,
    4712 => 61,
    4713 => 61,
    4714 => 61,
    4715 => 61,
    4716 => 61,
    4717 => 61,
    4718 => 61,
    4719 => 61,
    4720 => 61,
    4721 => 61,
    4722 => 61,
    4723 => 61,
    4724 => 61,
    4725 => 61,
    4726 => 61,
    4727 => 61,
    4728 => 61,
    4729 => 61,
    4730 => 61,
    4731 => 61,
    4732 => 61,
    4733 => 61,
    4734 => 61,
    4735 => 61,
    4736 => 61,
    4737 => 61,
    4738 => 61,
    4739 => 61,
    4740 => 61,
    4741 => 61,
    4742 => 61,
    4743 => 61,
    4744 => 61,
    4745 => 61,
    4746 => 61,
    4747 => 61,
    4748 => 61,
    4749 => 61,
    4750 => 61,
    4751 => 61,
    4752 => 61,
    4753 => 61,
    4754 => 61,
    4755 => 61,
    4756 => 61,
    4757 => 61,
    4758 => 61,
    4759 => 61,
    4760 => 61,
    4761 => 61,
    4762 => 61,
    4763 => 61,
    4764 => 61,
    4765 => 61,
    4766 => 61,
    4767 => 61,
    4768 => 61,
    4769 => 61,
    4770 => 61,
    4771 => 61,
    4772 => 61,
    4773 => 61,
    4774 => 61,
    4775 => 61,
    4776 => 61,
    4777 => 61,
    4778 => 61,
    4779 => 61,
    4780 => 61,
    4781 => 61,
    4782 => 61,
    4783 => 61,
    4784 => 61,
    4785 => 61,
    4786 => 61,
    4787 => 61,
    4788 => 61,
    4789 => 61,
    4790 => 61,
    4791 => 61,
    4792 => 61,
    4793 => 61,
    4794 => 61,
    4795 => 61,
    4796 => 61,
    4797 => 61,
    4798 => 61,
    4799 => 61,
    4800 => 61,
    4801 => 61,
    4802 => 61,
    4803 => 61,
    4804 => 61,
    4805 => 61,
    4806 => 61,
    4807 => 61,
    4808 => 61,
    4809 => 61,
    4810 => 61,
    4811 => 61,
    4812 => 61,
    4813 => 61,
    4814 => 61,
    4815 => 61,
    4816 => 61,
    4817 => 61,
    4818 => 61,
    4819 => 61,
    4820 => 61,
    4821 => 61,
    4822 => 61,
    4823 => 61,
    4824 => 61,
    4825 => 61,
    4826 => 61,
    4827 => 61,
    4828 => 61,
    4829 => 61,
    4830 => 61,
    4831 => 61,
    4832 => 61,
    4833 => 61,
    4834 => 60,
    4835 => 60,
    4836 => 60,
    4837 => 60,
    4838 => 60,
    4839 => 60,
    4840 => 60,
    4841 => 60,
    4842 => 60,
    4843 => 60,
    4844 => 60,
    4845 => 60,
    4846 => 60,
    4847 => 60,
    4848 => 60,
    4849 => 60,
    4850 => 60,
    4851 => 60,
    4852 => 60,
    4853 => 60,
    4854 => 60,
    4855 => 60,
    4856 => 60,
    4857 => 60,
    4858 => 60,
    4859 => 60,
    4860 => 60,
    4861 => 60,
    4862 => 60,
    4863 => 60,
    4864 => 60,
    4865 => 60,
    4866 => 60,
    4867 => 60,
    4868 => 60,
    4869 => 60,
    4870 => 60,
    4871 => 60,
    4872 => 60,
    4873 => 60,
    4874 => 60,
    4875 => 60,
    4876 => 60,
    4877 => 60,
    4878 => 60,
    4879 => 60,
    4880 => 60,
    4881 => 60,
    4882 => 60,
    4883 => 60,
    4884 => 60,
    4885 => 60,
    4886 => 60,
    4887 => 60,
    4888 => 60,
    4889 => 60,
    4890 => 60,
    4891 => 60,
    4892 => 60,
    4893 => 60,
    4894 => 60,
    4895 => 60,
    4896 => 60,
    4897 => 60,
    4898 => 60,
    4899 => 60,
    4900 => 60,
    4901 => 60,
    4902 => 60,
    4903 => 60,
    4904 => 60,
    4905 => 60,
    4906 => 60,
    4907 => 60,
    4908 => 60,
    4909 => 60,
    4910 => 60,
    4911 => 60,
    4912 => 60,
    4913 => 60,
    4914 => 60,
    4915 => 60,
    4916 => 60,
    4917 => 60,
    4918 => 60,
    4919 => 60,
    4920 => 60,
    4921 => 60,
    4922 => 60,
    4923 => 60,
    4924 => 60,
    4925 => 60,
    4926 => 60,
    4927 => 60,
    4928 => 60,
    4929 => 60,
    4930 => 60,
    4931 => 60,
    4932 => 60,
    4933 => 60,
    4934 => 60,
    4935 => 60,
    4936 => 60,
    4937 => 60,
    4938 => 60,
    4939 => 60,
    4940 => 60,
    4941 => 60,
    4942 => 60,
    4943 => 60,
    4944 => 60,
    4945 => 60,
    4946 => 60,
    4947 => 60,
    4948 => 60,
    4949 => 60,
    4950 => 60,
    4951 => 60,
    4952 => 60,
    4953 => 60,
    4954 => 60,
    4955 => 60,
    4956 => 60,
    4957 => 60,
    4958 => 60,
    4959 => 60,
    4960 => 60,
    4961 => 60,
    4962 => 60,
    4963 => 60,
    4964 => 60,
    4965 => 60,
    4966 => 60,
    4967 => 60,
    4968 => 60,
    4969 => 60,
    4970 => 59,
    4971 => 59,
    4972 => 59,
    4973 => 59,
    4974 => 59,
    4975 => 59,
    4976 => 59,
    4977 => 59,
    4978 => 59,
    4979 => 59,
    4980 => 59,
    4981 => 59,
    4982 => 59,
    4983 => 59,
    4984 => 59,
    4985 => 59,
    4986 => 59,
    4987 => 59,
    4988 => 59,
    4989 => 59,
    4990 => 59,
    4991 => 59,
    4992 => 59,
    4993 => 59,
    4994 => 59,
    4995 => 59,
    4996 => 59,
    4997 => 59,
    4998 => 59,
    4999 => 59,
    5000 => 59,
    5001 => 59,
    5002 => 59,
    5003 => 59,
    5004 => 59,
    5005 => 59,
    5006 => 59,
    5007 => 59,
    5008 => 59,
    5009 => 59,
    5010 => 59,
    5011 => 59,
    5012 => 59,
    5013 => 59,
    5014 => 59,
    5015 => 59,
    5016 => 59,
    5017 => 59,
    5018 => 59,
    5019 => 59,
    5020 => 59,
    5021 => 59,
    5022 => 59,
    5023 => 59,
    5024 => 59,
    5025 => 59,
    5026 => 59,
    5027 => 59,
    5028 => 59,
    5029 => 59,
    5030 => 59,
    5031 => 59,
    5032 => 59,
    5033 => 59,
    5034 => 59,
    5035 => 59,
    5036 => 59,
    5037 => 59,
    5038 => 59,
    5039 => 59,
    5040 => 59,
    5041 => 59,
    5042 => 59,
    5043 => 59,
    5044 => 59,
    5045 => 59,
    5046 => 59,
    5047 => 59,
    5048 => 59,
    5049 => 59,
    5050 => 59,
    5051 => 59,
    5052 => 59,
    5053 => 59,
    5054 => 59,
    5055 => 59,
    5056 => 59,
    5057 => 59,
    5058 => 59,
    5059 => 59,
    5060 => 59,
    5061 => 59,
    5062 => 59,
    5063 => 59,
    5064 => 59,
    5065 => 59,
    5066 => 59,
    5067 => 59,
    5068 => 59,
    5069 => 59,
    5070 => 59,
    5071 => 59,
    5072 => 59,
    5073 => 59,
    5074 => 59,
    5075 => 59,
    5076 => 59,
    5077 => 59,
    5078 => 59,
    5079 => 59,
    5080 => 59,
    5081 => 59,
    5082 => 59,
    5083 => 59,
    5084 => 59,
    5085 => 59,
    5086 => 59,
    5087 => 59,
    5088 => 58,
    5089 => 58,
    5090 => 58,
    5091 => 58,
    5092 => 58,
    5093 => 58,
    5094 => 58,
    5095 => 58,
    5096 => 58,
    5097 => 58,
    5098 => 58,
    5099 => 58,
    5100 => 58,
    5101 => 58,
    5102 => 58,
    5103 => 58,
    5104 => 58,
    5105 => 58,
    5106 => 58,
    5107 => 58,
    5108 => 58,
    5109 => 58,
    5110 => 58,
    5111 => 58,
    5112 => 58,
    5113 => 58,
    5114 => 58,
    5115 => 58,
    5116 => 58,
    5117 => 58,
    5118 => 58,
    5119 => 58,
    5120 => 58,
    5121 => 58,
    5122 => 58,
    5123 => 58,
    5124 => 58,
    5125 => 58,
    5126 => 58,
    5127 => 58,
    5128 => 58,
    5129 => 58,
    5130 => 58,
    5131 => 58,
    5132 => 58,
    5133 => 58,
    5134 => 58,
    5135 => 58,
    5136 => 58,
    5137 => 58,
    5138 => 58,
    5139 => 58,
    5140 => 58,
    5141 => 58,
    5142 => 58,
    5143 => 58,
    5144 => 58,
    5145 => 58,
    5146 => 58,
    5147 => 58,
    5148 => 58,
    5149 => 58,
    5150 => 58,
    5151 => 58,
    5152 => 58,
    5153 => 58,
    5154 => 58,
    5155 => 58,
    5156 => 58,
    5157 => 58,
    5158 => 58,
    5159 => 58,
    5160 => 58,
    5161 => 58,
    5162 => 58,
    5163 => 58,
    5164 => 58,
    5165 => 58,
    5166 => 58,
    5167 => 58,
    5168 => 58,
    5169 => 58,
    5170 => 58,
    5171 => 58,
    5172 => 58,
    5173 => 58,
    5174 => 58,
    5175 => 58,
    5176 => 58,
    5177 => 58,
    5178 => 58,
    5179 => 58,
    5180 => 58,
    5181 => 58,
    5182 => 58,
    5183 => 58,
    5184 => 58,
    5185 => 58,
    5186 => 58,
    5187 => 58,
    5188 => 58,
    5189 => 58,
    5190 => 58,
    5191 => 58,
    5192 => 58,
    5193 => 58,
    5194 => 57,
    5195 => 57,
    5196 => 57,
    5197 => 57,
    5198 => 57,
    5199 => 57,
    5200 => 57,
    5201 => 57,
    5202 => 57,
    5203 => 57,
    5204 => 57,
    5205 => 57,
    5206 => 57,
    5207 => 57,
    5208 => 57,
    5209 => 57,
    5210 => 57,
    5211 => 57,
    5212 => 57,
    5213 => 57,
    5214 => 57,
    5215 => 57,
    5216 => 57,
    5217 => 57,
    5218 => 57,
    5219 => 57,
    5220 => 57,
    5221 => 57,
    5222 => 57,
    5223 => 57,
    5224 => 57,
    5225 => 57,
    5226 => 57,
    5227 => 57,
    5228 => 57,
    5229 => 57,
    5230 => 57,
    5231 => 57,
    5232 => 57,
    5233 => 57,
    5234 => 57,
    5235 => 57,
    5236 => 57,
    5237 => 57,
    5238 => 57,
    5239 => 57,
    5240 => 57,
    5241 => 57,
    5242 => 57,
    5243 => 57,
    5244 => 57,
    5245 => 57,
    5246 => 57,
    5247 => 57,
    5248 => 57,
    5249 => 57,
    5250 => 57,
    5251 => 57,
    5252 => 57,
    5253 => 57,
    5254 => 57,
    5255 => 57,
    5256 => 57,
    5257 => 57,
    5258 => 57,
    5259 => 57,
    5260 => 57,
    5261 => 57,
    5262 => 57,
    5263 => 57,
    5264 => 57,
    5265 => 57,
    5266 => 57,
    5267 => 57,
    5268 => 57,
    5269 => 57,
    5270 => 57,
    5271 => 57,
    5272 => 57,
    5273 => 57,
    5274 => 57,
    5275 => 57,
    5276 => 57,
    5277 => 57,
    5278 => 57,
    5279 => 57,
    5280 => 57,
    5281 => 57,
    5282 => 57,
    5283 => 57,
    5284 => 57,
    5285 => 57,
    5286 => 57,
    5287 => 57,
    5288 => 57,
    5289 => 57,
    5290 => 57,
    5291 => 56,
    5292 => 56,
    5293 => 56,
    5294 => 56,
    5295 => 56,
    5296 => 56,
    5297 => 56,
    5298 => 56,
    5299 => 56,
    5300 => 56,
    5301 => 56,
    5302 => 56,
    5303 => 56,
    5304 => 56,
    5305 => 56,
    5306 => 56,
    5307 => 56,
    5308 => 56,
    5309 => 56,
    5310 => 56,
    5311 => 56,
    5312 => 56,
    5313 => 56,
    5314 => 56,
    5315 => 56,
    5316 => 56,
    5317 => 56,
    5318 => 56,
    5319 => 56,
    5320 => 56,
    5321 => 56,
    5322 => 56,
    5323 => 56,
    5324 => 56,
    5325 => 56,
    5326 => 56,
    5327 => 56,
    5328 => 56,
    5329 => 56,
    5330 => 56,
    5331 => 56,
    5332 => 56,
    5333 => 56,
    5334 => 56,
    5335 => 56,
    5336 => 56,
    5337 => 56,
    5338 => 56,
    5339 => 56,
    5340 => 56,
    5341 => 56,
    5342 => 56,
    5343 => 56,
    5344 => 56,
    5345 => 56,
    5346 => 56,
    5347 => 56,
    5348 => 56,
    5349 => 56,
    5350 => 56,
    5351 => 56,
    5352 => 56,
    5353 => 56,
    5354 => 56,
    5355 => 56,
    5356 => 56,
    5357 => 56,
    5358 => 56,
    5359 => 56,
    5360 => 56,
    5361 => 56,
    5362 => 56,
    5363 => 56,
    5364 => 56,
    5365 => 56,
    5366 => 56,
    5367 => 56,
    5368 => 56,
    5369 => 56,
    5370 => 56,
    5371 => 56,
    5372 => 56,
    5373 => 56,
    5374 => 56,
    5375 => 56,
    5376 => 56,
    5377 => 56,
    5378 => 56,
    5379 => 56,
    5380 => 56,
    5381 => 56,
    5382 => 55,
    5383 => 55,
    5384 => 55,
    5385 => 55,
    5386 => 55,
    5387 => 55,
    5388 => 55,
    5389 => 55,
    5390 => 55,
    5391 => 55,
    5392 => 55,
    5393 => 55,
    5394 => 55,
    5395 => 55,
    5396 => 55,
    5397 => 55,
    5398 => 55,
    5399 => 55,
    5400 => 55,
    5401 => 55,
    5402 => 55,
    5403 => 55,
    5404 => 55,
    5405 => 55,
    5406 => 55,
    5407 => 55,
    5408 => 55,
    5409 => 55,
    5410 => 55,
    5411 => 55,
    5412 => 55,
    5413 => 55,
    5414 => 55,
    5415 => 55,
    5416 => 55,
    5417 => 55,
    5418 => 55,
    5419 => 55,
    5420 => 55,
    5421 => 55,
    5422 => 55,
    5423 => 55,
    5424 => 55,
    5425 => 55,
    5426 => 55,
    5427 => 55,
    5428 => 55,
    5429 => 55,
    5430 => 55,
    5431 => 55,
    5432 => 55,
    5433 => 55,
    5434 => 55,
    5435 => 55,
    5436 => 55,
    5437 => 55,
    5438 => 55,
    5439 => 55,
    5440 => 55,
    5441 => 55,
    5442 => 55,
    5443 => 55,
    5444 => 55,
    5445 => 55,
    5446 => 55,
    5447 => 55,
    5448 => 55,
    5449 => 55,
    5450 => 55,
    5451 => 55,
    5452 => 55,
    5453 => 55,
    5454 => 55,
    5455 => 55,
    5456 => 55,
    5457 => 55,
    5458 => 55,
    5459 => 55,
    5460 => 55,
    5461 => 55,
    5462 => 55,
    5463 => 55,
    5464 => 55,
    5465 => 55,
    5466 => 55,
    5467 => 54,
    5468 => 54,
    5469 => 54,
    5470 => 54,
    5471 => 54,
    5472 => 54,
    5473 => 54,
    5474 => 54,
    5475 => 54,
    5476 => 54,
    5477 => 54,
    5478 => 54,
    5479 => 54,
    5480 => 54,
    5481 => 54,
    5482 => 54,
    5483 => 54,
    5484 => 54,
    5485 => 54,
    5486 => 54,
    5487 => 54,
    5488 => 54,
    5489 => 54,
    5490 => 54,
    5491 => 54,
    5492 => 54,
    5493 => 54,
    5494 => 54,
    5495 => 54,
    5496 => 54,
    5497 => 54,
    5498 => 54,
    5499 => 54,
    5500 => 54,
    5501 => 54,
    5502 => 54,
    5503 => 54,
    5504 => 54,
    5505 => 54,
    5506 => 54,
    5507 => 54,
    5508 => 54,
    5509 => 54,
    5510 => 54,
    5511 => 54,
    5512 => 54,
    5513 => 54,
    5514 => 54,
    5515 => 54,
    5516 => 54,
    5517 => 54,
    5518 => 54,
    5519 => 54,
    5520 => 54,
    5521 => 54,
    5522 => 54,
    5523 => 54,
    5524 => 54,
    5525 => 54,
    5526 => 54,
    5527 => 54,
    5528 => 54,
    5529 => 54,
    5530 => 54,
    5531 => 54,
    5532 => 54,
    5533 => 54,
    5534 => 54,
    5535 => 54,
    5536 => 54,
    5537 => 54,
    5538 => 54,
    5539 => 54,
    5540 => 54,
    5541 => 54,
    5542 => 54,
    5543 => 54,
    5544 => 54,
    5545 => 54,
    5546 => 54,
    5547 => 53,
    5548 => 53,
    5549 => 53,
    5550 => 53,
    5551 => 53,
    5552 => 53,
    5553 => 53,
    5554 => 53,
    5555 => 53,
    5556 => 53,
    5557 => 53,
    5558 => 53,
    5559 => 53,
    5560 => 53,
    5561 => 53,
    5562 => 53,
    5563 => 53,
    5564 => 53,
    5565 => 53,
    5566 => 53,
    5567 => 53,
    5568 => 53,
    5569 => 53,
    5570 => 53,
    5571 => 53,
    5572 => 53,
    5573 => 53,
    5574 => 53,
    5575 => 53,
    5576 => 53,
    5577 => 53,
    5578 => 53,
    5579 => 53,
    5580 => 53,
    5581 => 53,
    5582 => 53,
    5583 => 53,
    5584 => 53,
    5585 => 53,
    5586 => 53,
    5587 => 53,
    5588 => 53,
    5589 => 53,
    5590 => 53,
    5591 => 53,
    5592 => 53,
    5593 => 53,
    5594 => 53,
    5595 => 53,
    5596 => 53,
    5597 => 53,
    5598 => 53,
    5599 => 53,
    5600 => 53,
    5601 => 53,
    5602 => 53,
    5603 => 53,
    5604 => 53,
    5605 => 53,
    5606 => 53,
    5607 => 53,
    5608 => 53,
    5609 => 53,
    5610 => 53,
    5611 => 53,
    5612 => 53,
    5613 => 53,
    5614 => 53,
    5615 => 53,
    5616 => 53,
    5617 => 53,
    5618 => 53,
    5619 => 53,
    5620 => 53,
    5621 => 53,
    5622 => 53,
    5623 => 53,
    5624 => 52,
    5625 => 52,
    5626 => 52,
    5627 => 52,
    5628 => 52,
    5629 => 52,
    5630 => 52,
    5631 => 52,
    5632 => 52,
    5633 => 52,
    5634 => 52,
    5635 => 52,
    5636 => 52,
    5637 => 52,
    5638 => 52,
    5639 => 52,
    5640 => 52,
    5641 => 52,
    5642 => 52,
    5643 => 52,
    5644 => 52,
    5645 => 52,
    5646 => 52,
    5647 => 52,
    5648 => 52,
    5649 => 52,
    5650 => 52,
    5651 => 52,
    5652 => 52,
    5653 => 52,
    5654 => 52,
    5655 => 52,
    5656 => 52,
    5657 => 52,
    5658 => 52,
    5659 => 52,
    5660 => 52,
    5661 => 52,
    5662 => 52,
    5663 => 52,
    5664 => 52,
    5665 => 52,
    5666 => 52,
    5667 => 52,
    5668 => 52,
    5669 => 52,
    5670 => 52,
    5671 => 52,
    5672 => 52,
    5673 => 52,
    5674 => 52,
    5675 => 52,
    5676 => 52,
    5677 => 52,
    5678 => 52,
    5679 => 52,
    5680 => 52,
    5681 => 52,
    5682 => 52,
    5683 => 52,
    5684 => 52,
    5685 => 52,
    5686 => 52,
    5687 => 52,
    5688 => 52,
    5689 => 52,
    5690 => 52,
    5691 => 52,
    5692 => 52,
    5693 => 52,
    5694 => 52,
    5695 => 52,
    5696 => 52,
    5697 => 51,
    5698 => 51,
    5699 => 51,
    5700 => 51,
    5701 => 51,
    5702 => 51,
    5703 => 51,
    5704 => 51,
    5705 => 51,
    5706 => 51,
    5707 => 51,
    5708 => 51,
    5709 => 51,
    5710 => 51,
    5711 => 51,
    5712 => 51,
    5713 => 51,
    5714 => 51,
    5715 => 51,
    5716 => 51,
    5717 => 51,
    5718 => 51,
    5719 => 51,
    5720 => 51,
    5721 => 51,
    5722 => 51,
    5723 => 51,
    5724 => 51,
    5725 => 51,
    5726 => 51,
    5727 => 51,
    5728 => 51,
    5729 => 51,
    5730 => 51,
    5731 => 51,
    5732 => 51,
    5733 => 51,
    5734 => 51,
    5735 => 51,
    5736 => 51,
    5737 => 51,
    5738 => 51,
    5739 => 51,
    5740 => 51,
    5741 => 51,
    5742 => 51,
    5743 => 51,
    5744 => 51,
    5745 => 51,
    5746 => 51,
    5747 => 51,
    5748 => 51,
    5749 => 51,
    5750 => 51,
    5751 => 51,
    5752 => 51,
    5753 => 51,
    5754 => 51,
    5755 => 51,
    5756 => 51,
    5757 => 51,
    5758 => 51,
    5759 => 51,
    5760 => 51,
    5761 => 51,
    5762 => 51,
    5763 => 51,
    5764 => 51,
    5765 => 51,
    5766 => 51,
    5767 => 51,
    5768 => 50,
    5769 => 50,
    5770 => 50,
    5771 => 50,
    5772 => 50,
    5773 => 50,
    5774 => 50,
    5775 => 50,
    5776 => 50,
    5777 => 50,
    5778 => 50,
    5779 => 50,
    5780 => 50,
    5781 => 50,
    5782 => 50,
    5783 => 50,
    5784 => 50,
    5785 => 50,
    5786 => 50,
    5787 => 50,
    5788 => 50,
    5789 => 50,
    5790 => 50,
    5791 => 50,
    5792 => 50,
    5793 => 50,
    5794 => 50,
    5795 => 50,
    5796 => 50,
    5797 => 50,
    5798 => 50,
    5799 => 50,
    5800 => 50,
    5801 => 50,
    5802 => 50,
    5803 => 50,
    5804 => 50,
    5805 => 50,
    5806 => 50,
    5807 => 50,
    5808 => 50,
    5809 => 50,
    5810 => 50,
    5811 => 50,
    5812 => 50,
    5813 => 50,
    5814 => 50,
    5815 => 50,
    5816 => 50,
    5817 => 50,
    5818 => 50,
    5819 => 50,
    5820 => 50,
    5821 => 50,
    5822 => 50,
    5823 => 50,
    5824 => 50,
    5825 => 50,
    5826 => 50,
    5827 => 50,
    5828 => 50,
    5829 => 50,
    5830 => 50,
    5831 => 50,
    5832 => 50,
    5833 => 50,
    5834 => 50,
    5835 => 50,
    5836 => 49,
    5837 => 49,
    5838 => 49,
    5839 => 49,
    5840 => 49,
    5841 => 49,
    5842 => 49,
    5843 => 49,
    5844 => 49,
    5845 => 49,
    5846 => 49,
    5847 => 49,
    5848 => 49,
    5849 => 49,
    5850 => 49,
    5851 => 49,
    5852 => 49,
    5853 => 49,
    5854 => 49,
    5855 => 49,
    5856 => 49,
    5857 => 49,
    5858 => 49,
    5859 => 49,
    5860 => 49,
    5861 => 49,
    5862 => 49,
    5863 => 49,
    5864 => 49,
    5865 => 49,
    5866 => 49,
    5867 => 49,
    5868 => 49,
    5869 => 49,
    5870 => 49,
    5871 => 49,
    5872 => 49,
    5873 => 49,
    5874 => 49,
    5875 => 49,
    5876 => 49,
    5877 => 49,
    5878 => 49,
    5879 => 49,
    5880 => 49,
    5881 => 49,
    5882 => 49,
    5883 => 49,
    5884 => 49,
    5885 => 49,
    5886 => 49,
    5887 => 49,
    5888 => 49,
    5889 => 49,
    5890 => 49,
    5891 => 49,
    5892 => 49,
    5893 => 49,
    5894 => 49,
    5895 => 49,
    5896 => 49,
    5897 => 49,
    5898 => 49,
    5899 => 49,
    5900 => 49,
    5901 => 48,
    5902 => 48,
    5903 => 48,
    5904 => 48,
    5905 => 48,
    5906 => 48,
    5907 => 48,
    5908 => 48,
    5909 => 48,
    5910 => 48,
    5911 => 48,
    5912 => 48,
    5913 => 48,
    5914 => 48,
    5915 => 48,
    5916 => 48,
    5917 => 48,
    5918 => 48,
    5919 => 48,
    5920 => 48,
    5921 => 48,
    5922 => 48,
    5923 => 48,
    5924 => 48,
    5925 => 48,
    5926 => 48,
    5927 => 48,
    5928 => 48,
    5929 => 48,
    5930 => 48,
    5931 => 48,
    5932 => 48,
    5933 => 48,
    5934 => 48,
    5935 => 48,
    5936 => 48,
    5937 => 48,
    5938 => 48,
    5939 => 48,
    5940 => 48,
    5941 => 48,
    5942 => 48,
    5943 => 48,
    5944 => 48,
    5945 => 48,
    5946 => 48,
    5947 => 48,
    5948 => 48,
    5949 => 48,
    5950 => 48,
    5951 => 48,
    5952 => 48,
    5953 => 48,
    5954 => 48,
    5955 => 48,
    5956 => 48,
    5957 => 48,
    5958 => 48,
    5959 => 48,
    5960 => 48,
    5961 => 48,
    5962 => 48,
    5963 => 48,
    5964 => 48,
    5965 => 47,
    5966 => 47,
    5967 => 47,
    5968 => 47,
    5969 => 47,
    5970 => 47,
    5971 => 47,
    5972 => 47,
    5973 => 47,
    5974 => 47,
    5975 => 47,
    5976 => 47,
    5977 => 47,
    5978 => 47,
    5979 => 47,
    5980 => 47,
    5981 => 47,
    5982 => 47,
    5983 => 47,
    5984 => 47,
    5985 => 47,
    5986 => 47,
    5987 => 47,
    5988 => 47,
    5989 => 47,
    5990 => 47,
    5991 => 47,
    5992 => 47,
    5993 => 47,
    5994 => 47,
    5995 => 47,
    5996 => 47,
    5997 => 47,
    5998 => 47,
    5999 => 47,
    6000 => 47,
    6001 => 47,
    6002 => 47,
    6003 => 47,
    6004 => 47,
    6005 => 47,
    6006 => 47,
    6007 => 47,
    6008 => 47,
    6009 => 47,
    6010 => 47,
    6011 => 47,
    6012 => 47,
    6013 => 47,
    6014 => 47,
    6015 => 47,
    6016 => 47,
    6017 => 47,
    6018 => 47,
    6019 => 47,
    6020 => 47,
    6021 => 47,
    6022 => 47,
    6023 => 47,
    6024 => 47,
    6025 => 47,
    6026 => 47,
    6027 => 47,
    6028 => 46,
    6029 => 46,
    6030 => 46,
    6031 => 46,
    6032 => 46,
    6033 => 46,
    6034 => 46,
    6035 => 46,
    6036 => 46,
    6037 => 46,
    6038 => 46,
    6039 => 46,
    6040 => 46,
    6041 => 46,
    6042 => 46,
    6043 => 46,
    6044 => 46,
    6045 => 46,
    6046 => 46,
    6047 => 46,
    6048 => 46,
    6049 => 46,
    6050 => 46,
    6051 => 46,
    6052 => 46,
    6053 => 46,
    6054 => 46,
    6055 => 46,
    6056 => 46,
    6057 => 46,
    6058 => 46,
    6059 => 46,
    6060 => 46,
    6061 => 46,
    6062 => 46,
    6063 => 46,
    6064 => 46,
    6065 => 46,
    6066 => 46,
    6067 => 46,
    6068 => 46,
    6069 => 46,
    6070 => 46,
    6071 => 46,
    6072 => 46,
    6073 => 46,
    6074 => 46,
    6075 => 46,
    6076 => 46,
    6077 => 46,
    6078 => 46,
    6079 => 46,
    6080 => 46,
    6081 => 46,
    6082 => 46,
    6083 => 46,
    6084 => 46,
    6085 => 46,
    6086 => 46,
    6087 => 46,
    6088 => 45,
    6089 => 45,
    6090 => 45,
    6091 => 45,
    6092 => 45,
    6093 => 45,
    6094 => 45,
    6095 => 45,
    6096 => 45,
    6097 => 45,
    6098 => 45,
    6099 => 45,
    6100 => 45,
    6101 => 45,
    6102 => 45,
    6103 => 45,
    6104 => 45,
    6105 => 45,
    6106 => 45,
    6107 => 45,
    6108 => 45,
    6109 => 45,
    6110 => 45,
    6111 => 45,
    6112 => 45,
    6113 => 45,
    6114 => 45,
    6115 => 45,
    6116 => 45,
    6117 => 45,
    6118 => 45,
    6119 => 45,
    6120 => 45,
    6121 => 45,
    6122 => 45,
    6123 => 45,
    6124 => 45,
    6125 => 45,
    6126 => 45,
    6127 => 45,
    6128 => 45,
    6129 => 45,
    6130 => 45,
    6131 => 45,
    6132 => 45,
    6133 => 45,
    6134 => 45,
    6135 => 45,
    6136 => 45,
    6137 => 45,
    6138 => 45,
    6139 => 45,
    6140 => 45,
    6141 => 45,
    6142 => 45,
    6143 => 45,
    6144 => 45,
    6145 => 45,
    6146 => 45,
    6147 => 44,
    6148 => 44,
    6149 => 44,
    6150 => 44,
    6151 => 44,
    6152 => 44,
    6153 => 44,
    6154 => 44,
    6155 => 44,
    6156 => 44,
    6157 => 44,
    6158 => 44,
    6159 => 44,
    6160 => 44,
    6161 => 44,
    6162 => 44,
    6163 => 44,
    6164 => 44,
    6165 => 44,
    6166 => 44,
    6167 => 44,
    6168 => 44,
    6169 => 44,
    6170 => 44,
    6171 => 44,
    6172 => 44,
    6173 => 44,
    6174 => 44,
    6175 => 44,
    6176 => 44,
    6177 => 44,
    6178 => 44,
    6179 => 44,
    6180 => 44,
    6181 => 44,
    6182 => 44,
    6183 => 44,
    6184 => 44,
    6185 => 44,
    6186 => 44,
    6187 => 44,
    6188 => 44,
    6189 => 44,
    6190 => 44,
    6191 => 44,
    6192 => 44,
    6193 => 44,
    6194 => 44,
    6195 => 44,
    6196 => 44,
    6197 => 44,
    6198 => 44,
    6199 => 44,
    6200 => 44,
    6201 => 44,
    6202 => 44,
    6203 => 44,
    6204 => 44,
    6205 => 43,
    6206 => 43,
    6207 => 43,
    6208 => 43,
    6209 => 43,
    6210 => 43,
    6211 => 43,
    6212 => 43,
    6213 => 43,
    6214 => 43,
    6215 => 43,
    6216 => 43,
    6217 => 43,
    6218 => 43,
    6219 => 43,
    6220 => 43,
    6221 => 43,
    6222 => 43,
    6223 => 43,
    6224 => 43,
    6225 => 43,
    6226 => 43,
    6227 => 43,
    6228 => 43,
    6229 => 43,
    6230 => 43,
    6231 => 43,
    6232 => 43,
    6233 => 43,
    6234 => 43,
    6235 => 43,
    6236 => 43,
    6237 => 43,
    6238 => 43,
    6239 => 43,
    6240 => 43,
    6241 => 43,
    6242 => 43,
    6243 => 43,
    6244 => 43,
    6245 => 43,
    6246 => 43,
    6247 => 43,
    6248 => 43,
    6249 => 43,
    6250 => 43,
    6251 => 43,
    6252 => 43,
    6253 => 43,
    6254 => 43,
    6255 => 43,
    6256 => 43,
    6257 => 43,
    6258 => 43,
    6259 => 43,
    6260 => 43,
    6261 => 43,
    6262 => 42,
    6263 => 42,
    6264 => 42,
    6265 => 42,
    6266 => 42,
    6267 => 42,
    6268 => 42,
    6269 => 42,
    6270 => 42,
    6271 => 42,
    6272 => 42,
    6273 => 42,
    6274 => 42,
    6275 => 42,
    6276 => 42,
    6277 => 42,
    6278 => 42,
    6279 => 42,
    6280 => 42,
    6281 => 42,
    6282 => 42,
    6283 => 42,
    6284 => 42,
    6285 => 42,
    6286 => 42,
    6287 => 42,
    6288 => 42,
    6289 => 42,
    6290 => 42,
    6291 => 42,
    6292 => 42,
    6293 => 42,
    6294 => 42,
    6295 => 42,
    6296 => 42,
    6297 => 42,
    6298 => 42,
    6299 => 42,
    6300 => 42,
    6301 => 42,
    6302 => 42,
    6303 => 42,
    6304 => 42,
    6305 => 42,
    6306 => 42,
    6307 => 42,
    6308 => 42,
    6309 => 42,
    6310 => 42,
    6311 => 42,
    6312 => 42,
    6313 => 42,
    6314 => 42,
    6315 => 42,
    6316 => 42,
    6317 => 41,
    6318 => 41,
    6319 => 41,
    6320 => 41,
    6321 => 41,
    6322 => 41,
    6323 => 41,
    6324 => 41,
    6325 => 41,
    6326 => 41,
    6327 => 41,
    6328 => 41,
    6329 => 41,
    6330 => 41,
    6331 => 41,
    6332 => 41,
    6333 => 41,
    6334 => 41,
    6335 => 41,
    6336 => 41,
    6337 => 41,
    6338 => 41,
    6339 => 41,
    6340 => 41,
    6341 => 41,
    6342 => 41,
    6343 => 41,
    6344 => 41,
    6345 => 41,
    6346 => 41,
    6347 => 41,
    6348 => 41,
    6349 => 41,
    6350 => 41,
    6351 => 41,
    6352 => 41,
    6353 => 41,
    6354 => 41,
    6355 => 41,
    6356 => 41,
    6357 => 41,
    6358 => 41,
    6359 => 41,
    6360 => 41,
    6361 => 41,
    6362 => 41,
    6363 => 41,
    6364 => 41,
    6365 => 41,
    6366 => 41,
    6367 => 41,
    6368 => 41,
    6369 => 41,
    6370 => 41,
    6371 => 41,
    6372 => 40,
    6373 => 40,
    6374 => 40,
    6375 => 40,
    6376 => 40,
    6377 => 40,
    6378 => 40,
    6379 => 40,
    6380 => 40,
    6381 => 40,
    6382 => 40,
    6383 => 40,
    6384 => 40,
    6385 => 40,
    6386 => 40,
    6387 => 40,
    6388 => 40,
    6389 => 40,
    6390 => 40,
    6391 => 40,
    6392 => 40,
    6393 => 40,
    6394 => 40,
    6395 => 40,
    6396 => 40,
    6397 => 40,
    6398 => 40,
    6399 => 40,
    6400 => 40,
    6401 => 40,
    6402 => 40,
    6403 => 40,
    6404 => 40,
    6405 => 40,
    6406 => 40,
    6407 => 40,
    6408 => 40,
    6409 => 40,
    6410 => 40,
    6411 => 40,
    6412 => 40,
    6413 => 40,
    6414 => 40,
    6415 => 40,
    6416 => 40,
    6417 => 40,
    6418 => 40,
    6419 => 40,
    6420 => 40,
    6421 => 40,
    6422 => 40,
    6423 => 40,
    6424 => 40,
    6425 => 39,
    6426 => 39,
    6427 => 39,
    6428 => 39,
    6429 => 39,
    6430 => 39,
    6431 => 39,
    6432 => 39,
    6433 => 39,
    6434 => 39,
    6435 => 39,
    6436 => 39,
    6437 => 39,
    6438 => 39,
    6439 => 39,
    6440 => 39,
    6441 => 39,
    6442 => 39,
    6443 => 39,
    6444 => 39,
    6445 => 39,
    6446 => 39,
    6447 => 39,
    6448 => 39,
    6449 => 39,
    6450 => 39,
    6451 => 39,
    6452 => 39,
    6453 => 39,
    6454 => 39,
    6455 => 39,
    6456 => 39,
    6457 => 39,
    6458 => 39,
    6459 => 39,
    6460 => 39,
    6461 => 39,
    6462 => 39,
    6463 => 39,
    6464 => 39,
    6465 => 39,
    6466 => 39,
    6467 => 39,
    6468 => 39,
    6469 => 39,
    6470 => 39,
    6471 => 39,
    6472 => 39,
    6473 => 39,
    6474 => 39,
    6475 => 39,
    6476 => 39,
    6477 => 39,
    6478 => 38,
    6479 => 38,
    6480 => 38,
    6481 => 38,
    6482 => 38,
    6483 => 38,
    6484 => 38,
    6485 => 38,
    6486 => 38,
    6487 => 38,
    6488 => 38,
    6489 => 38,
    6490 => 38,
    6491 => 38,
    6492 => 38,
    6493 => 38,
    6494 => 38,
    6495 => 38,
    6496 => 38,
    6497 => 38,
    6498 => 38,
    6499 => 38,
    6500 => 38,
    6501 => 38,
    6502 => 38,
    6503 => 38,
    6504 => 38,
    6505 => 38,
    6506 => 38,
    6507 => 38,
    6508 => 38,
    6509 => 38,
    6510 => 38,
    6511 => 38,
    6512 => 38,
    6513 => 38,
    6514 => 38,
    6515 => 38,
    6516 => 38,
    6517 => 38,
    6518 => 38,
    6519 => 38,
    6520 => 38,
    6521 => 38,
    6522 => 38,
    6523 => 38,
    6524 => 38,
    6525 => 38,
    6526 => 38,
    6527 => 38,
    6528 => 38,
    6529 => 38,
    6530 => 37,
    6531 => 37,
    6532 => 37,
    6533 => 37,
    6534 => 37,
    6535 => 37,
    6536 => 37,
    6537 => 37,
    6538 => 37,
    6539 => 37,
    6540 => 37,
    6541 => 37,
    6542 => 37,
    6543 => 37,
    6544 => 37,
    6545 => 37,
    6546 => 37,
    6547 => 37,
    6548 => 37,
    6549 => 37,
    6550 => 37,
    6551 => 37,
    6552 => 37,
    6553 => 37,
    6554 => 37,
    6555 => 37,
    6556 => 37,
    6557 => 37,
    6558 => 37,
    6559 => 37,
    6560 => 37,
    6561 => 37,
    6562 => 37,
    6563 => 37,
    6564 => 37,
    6565 => 37,
    6566 => 37,
    6567 => 37,
    6568 => 37,
    6569 => 37,
    6570 => 37,
    6571 => 37,
    6572 => 37,
    6573 => 37,
    6574 => 37,
    6575 => 37,
    6576 => 37,
    6577 => 37,
    6578 => 37,
    6579 => 37,
    6580 => 37,
    6581 => 36,
    6582 => 36,
    6583 => 36,
    6584 => 36,
    6585 => 36,
    6586 => 36,
    6587 => 36,
    6588 => 36,
    6589 => 36,
    6590 => 36,
    6591 => 36,
    6592 => 36,
    6593 => 36,
    6594 => 36,
    6595 => 36,
    6596 => 36,
    6597 => 36,
    6598 => 36,
    6599 => 36,
    6600 => 36,
    6601 => 36,
    6602 => 36,
    6603 => 36,
    6604 => 36,
    6605 => 36,
    6606 => 36,
    6607 => 36,
    6608 => 36,
    6609 => 36,
    6610 => 36,
    6611 => 36,
    6612 => 36,
    6613 => 36,
    6614 => 36,
    6615 => 36,
    6616 => 36,
    6617 => 36,
    6618 => 36,
    6619 => 36,
    6620 => 36,
    6621 => 36,
    6622 => 36,
    6623 => 36,
    6624 => 36,
    6625 => 36,
    6626 => 36,
    6627 => 36,
    6628 => 36,
    6629 => 36,
    6630 => 36,
    6631 => 36,
    6632 => 35,
    6633 => 35,
    6634 => 35,
    6635 => 35,
    6636 => 35,
    6637 => 35,
    6638 => 35,
    6639 => 35,
    6640 => 35,
    6641 => 35,
    6642 => 35,
    6643 => 35,
    6644 => 35,
    6645 => 35,
    6646 => 35,
    6647 => 35,
    6648 => 35,
    6649 => 35,
    6650 => 35,
    6651 => 35,
    6652 => 35,
    6653 => 35,
    6654 => 35,
    6655 => 35,
    6656 => 35,
    6657 => 35,
    6658 => 35,
    6659 => 35,
    6660 => 35,
    6661 => 35,
    6662 => 35,
    6663 => 35,
    6664 => 35,
    6665 => 35,
    6666 => 35,
    6667 => 35,
    6668 => 35,
    6669 => 35,
    6670 => 35,
    6671 => 35,
    6672 => 35,
    6673 => 35,
    6674 => 35,
    6675 => 35,
    6676 => 35,
    6677 => 35,
    6678 => 35,
    6679 => 35,
    6680 => 35,
    6681 => 34,
    6682 => 34,
    6683 => 34,
    6684 => 34,
    6685 => 34,
    6686 => 34,
    6687 => 34,
    6688 => 34,
    6689 => 34,
    6690 => 34,
    6691 => 34,
    6692 => 34,
    6693 => 34,
    6694 => 34,
    6695 => 34,
    6696 => 34,
    6697 => 34,
    6698 => 34,
    6699 => 34,
    6700 => 34,
    6701 => 34,
    6702 => 34,
    6703 => 34,
    6704 => 34,
    6705 => 34,
    6706 => 34,
    6707 => 34,
    6708 => 34,
    6709 => 34,
    6710 => 34,
    6711 => 34,
    6712 => 34,
    6713 => 34,
    6714 => 34,
    6715 => 34,
    6716 => 34,
    6717 => 34,
    6718 => 34,
    6719 => 34,
    6720 => 34,
    6721 => 34,
    6722 => 34,
    6723 => 34,
    6724 => 34,
    6725 => 34,
    6726 => 34,
    6727 => 34,
    6728 => 34,
    6729 => 34,
    6730 => 34,
    6731 => 33,
    6732 => 33,
    6733 => 33,
    6734 => 33,
    6735 => 33,
    6736 => 33,
    6737 => 33,
    6738 => 33,
    6739 => 33,
    6740 => 33,
    6741 => 33,
    6742 => 33,
    6743 => 33,
    6744 => 33,
    6745 => 33,
    6746 => 33,
    6747 => 33,
    6748 => 33,
    6749 => 33,
    6750 => 33,
    6751 => 33,
    6752 => 33,
    6753 => 33,
    6754 => 33,
    6755 => 33,
    6756 => 33,
    6757 => 33,
    6758 => 33,
    6759 => 33,
    6760 => 33,
    6761 => 33,
    6762 => 33,
    6763 => 33,
    6764 => 33,
    6765 => 33,
    6766 => 33,
    6767 => 33,
    6768 => 33,
    6769 => 33,
    6770 => 33,
    6771 => 33,
    6772 => 33,
    6773 => 33,
    6774 => 33,
    6775 => 33,
    6776 => 33,
    6777 => 33,
    6778 => 33,
    6779 => 32,
    6780 => 32,
    6781 => 32,
    6782 => 32,
    6783 => 32,
    6784 => 32,
    6785 => 32,
    6786 => 32,
    6787 => 32,
    6788 => 32,
    6789 => 32,
    6790 => 32,
    6791 => 32,
    6792 => 32,
    6793 => 32,
    6794 => 32,
    6795 => 32,
    6796 => 32,
    6797 => 32,
    6798 => 32,
    6799 => 32,
    6800 => 32,
    6801 => 32,
    6802 => 32,
    6803 => 32,
    6804 => 32,
    6805 => 32,
    6806 => 32,
    6807 => 32,
    6808 => 32,
    6809 => 32,
    6810 => 32,
    6811 => 32,
    6812 => 32,
    6813 => 32,
    6814 => 32,
    6815 => 32,
    6816 => 32,
    6817 => 32,
    6818 => 32,
    6819 => 32,
    6820 => 32,
    6821 => 32,
    6822 => 32,
    6823 => 32,
    6824 => 32,
    6825 => 32,
    6826 => 32,
    6827 => 31,
    6828 => 31,
    6829 => 31,
    6830 => 31,
    6831 => 31,
    6832 => 31,
    6833 => 31,
    6834 => 31,
    6835 => 31,
    6836 => 31,
    6837 => 31,
    6838 => 31,
    6839 => 31,
    6840 => 31,
    6841 => 31,
    6842 => 31,
    6843 => 31,
    6844 => 31,
    6845 => 31,
    6846 => 31,
    6847 => 31,
    6848 => 31,
    6849 => 31,
    6850 => 31,
    6851 => 31,
    6852 => 31,
    6853 => 31,
    6854 => 31,
    6855 => 31,
    6856 => 31,
    6857 => 31,
    6858 => 31,
    6859 => 31,
    6860 => 31,
    6861 => 31,
    6862 => 31,
    6863 => 31,
    6864 => 31,
    6865 => 31,
    6866 => 31,
    6867 => 31,
    6868 => 31,
    6869 => 31,
    6870 => 31,
    6871 => 31,
    6872 => 31,
    6873 => 31,
    6874 => 31,
    6875 => 30,
    6876 => 30,
    6877 => 30,
    6878 => 30,
    6879 => 30,
    6880 => 30,
    6881 => 30,
    6882 => 30,
    6883 => 30,
    6884 => 30,
    6885 => 30,
    6886 => 30,
    6887 => 30,
    6888 => 30,
    6889 => 30,
    6890 => 30,
    6891 => 30,
    6892 => 30,
    6893 => 30,
    6894 => 30,
    6895 => 30,
    6896 => 30,
    6897 => 30,
    6898 => 30,
    6899 => 30,
    6900 => 30,
    6901 => 30,
    6902 => 30,
    6903 => 30,
    6904 => 30,
    6905 => 30,
    6906 => 30,
    6907 => 30,
    6908 => 30,
    6909 => 30,
    6910 => 30,
    6911 => 30,
    6912 => 30,
    6913 => 30,
    6914 => 30,
    6915 => 30,
    6916 => 30,
    6917 => 30,
    6918 => 30,
    6919 => 30,
    6920 => 30,
    6921 => 30,
    6922 => 29,
    6923 => 29,
    6924 => 29,
    6925 => 29,
    6926 => 29,
    6927 => 29,
    6928 => 29,
    6929 => 29,
    6930 => 29,
    6931 => 29,
    6932 => 29,
    6933 => 29,
    6934 => 29,
    6935 => 29,
    6936 => 29,
    6937 => 29,
    6938 => 29,
    6939 => 29,
    6940 => 29,
    6941 => 29,
    6942 => 29,
    6943 => 29,
    6944 => 29,
    6945 => 29,
    6946 => 29,
    6947 => 29,
    6948 => 29,
    6949 => 29,
    6950 => 29,
    6951 => 29,
    6952 => 29,
    6953 => 29,
    6954 => 29,
    6955 => 29,
    6956 => 29,
    6957 => 29,
    6958 => 29,
    6959 => 29,
    6960 => 29,
    6961 => 29,
    6962 => 29,
    6963 => 29,
    6964 => 29,
    6965 => 29,
    6966 => 29,
    6967 => 29,
    6968 => 28,
    6969 => 28,
    6970 => 28,
    6971 => 28,
    6972 => 28,
    6973 => 28,
    6974 => 28,
    6975 => 28,
    6976 => 28,
    6977 => 28,
    6978 => 28,
    6979 => 28,
    6980 => 28,
    6981 => 28,
    6982 => 28,
    6983 => 28,
    6984 => 28,
    6985 => 28,
    6986 => 28,
    6987 => 28,
    6988 => 28,
    6989 => 28,
    6990 => 28,
    6991 => 28,
    6992 => 28,
    6993 => 28,
    6994 => 28,
    6995 => 28,
    6996 => 28,
    6997 => 28,
    6998 => 28,
    6999 => 28,
    7000 => 28,
    7001 => 28,
    7002 => 28,
    7003 => 28,
    7004 => 28,
    7005 => 28,
    7006 => 28,
    7007 => 28,
    7008 => 28,
    7009 => 28,
    7010 => 28,
    7011 => 28,
    7012 => 28,
    7013 => 28,
    7014 => 28,
    7015 => 27,
    7016 => 27,
    7017 => 27,
    7018 => 27,
    7019 => 27,
    7020 => 27,
    7021 => 27,
    7022 => 27,
    7023 => 27,
    7024 => 27,
    7025 => 27,
    7026 => 27,
    7027 => 27,
    7028 => 27,
    7029 => 27,
    7030 => 27,
    7031 => 27,
    7032 => 27,
    7033 => 27,
    7034 => 27,
    7035 => 27,
    7036 => 27,
    7037 => 27,
    7038 => 27,
    7039 => 27,
    7040 => 27,
    7041 => 27,
    7042 => 27,
    7043 => 27,
    7044 => 27,
    7045 => 27,
    7046 => 27,
    7047 => 27,
    7048 => 27,
    7049 => 27,
    7050 => 27,
    7051 => 27,
    7052 => 27,
    7053 => 27,
    7054 => 27,
    7055 => 27,
    7056 => 27,
    7057 => 27,
    7058 => 27,
    7059 => 27,
    7060 => 26,
    7061 => 26,
    7062 => 26,
    7063 => 26,
    7064 => 26,
    7065 => 26,
    7066 => 26,
    7067 => 26,
    7068 => 26,
    7069 => 26,
    7070 => 26,
    7071 => 26,
    7072 => 26,
    7073 => 26,
    7074 => 26,
    7075 => 26,
    7076 => 26,
    7077 => 26,
    7078 => 26,
    7079 => 26,
    7080 => 26,
    7081 => 26,
    7082 => 26,
    7083 => 26,
    7084 => 26,
    7085 => 26,
    7086 => 26,
    7087 => 26,
    7088 => 26,
    7089 => 26,
    7090 => 26,
    7091 => 26,
    7092 => 26,
    7093 => 26,
    7094 => 26,
    7095 => 26,
    7096 => 26,
    7097 => 26,
    7098 => 26,
    7099 => 26,
    7100 => 26,
    7101 => 26,
    7102 => 26,
    7103 => 26,
    7104 => 26,
    7105 => 26,
    7106 => 25,
    7107 => 25,
    7108 => 25,
    7109 => 25,
    7110 => 25,
    7111 => 25,
    7112 => 25,
    7113 => 25,
    7114 => 25,
    7115 => 25,
    7116 => 25,
    7117 => 25,
    7118 => 25,
    7119 => 25,
    7120 => 25,
    7121 => 25,
    7122 => 25,
    7123 => 25,
    7124 => 25,
    7125 => 25,
    7126 => 25,
    7127 => 25,
    7128 => 25,
    7129 => 25,
    7130 => 25,
    7131 => 25,
    7132 => 25,
    7133 => 25,
    7134 => 25,
    7135 => 25,
    7136 => 25,
    7137 => 25,
    7138 => 25,
    7139 => 25,
    7140 => 25,
    7141 => 25,
    7142 => 25,
    7143 => 25,
    7144 => 25,
    7145 => 25,
    7146 => 25,
    7147 => 25,
    7148 => 25,
    7149 => 25,
    7150 => 25,
    7151 => 24,
    7152 => 24,
    7153 => 24,
    7154 => 24,
    7155 => 24,
    7156 => 24,
    7157 => 24,
    7158 => 24,
    7159 => 24,
    7160 => 24,
    7161 => 24,
    7162 => 24,
    7163 => 24,
    7164 => 24,
    7165 => 24,
    7166 => 24,
    7167 => 24,
    7168 => 24,
    7169 => 24,
    7170 => 24,
    7171 => 24,
    7172 => 24,
    7173 => 24,
    7174 => 24,
    7175 => 24,
    7176 => 24,
    7177 => 24,
    7178 => 24,
    7179 => 24,
    7180 => 24,
    7181 => 24,
    7182 => 24,
    7183 => 24,
    7184 => 24,
    7185 => 24,
    7186 => 24,
    7187 => 24,
    7188 => 24,
    7189 => 24,
    7190 => 24,
    7191 => 24,
    7192 => 24,
    7193 => 24,
    7194 => 24,
    7195 => 24,
    7196 => 23,
    7197 => 23,
    7198 => 23,
    7199 => 23,
    7200 => 23,
    7201 => 23,
    7202 => 23,
    7203 => 23,
    7204 => 23,
    7205 => 23,
    7206 => 23,
    7207 => 23,
    7208 => 23,
    7209 => 23,
    7210 => 23,
    7211 => 23,
    7212 => 23,
    7213 => 23,
    7214 => 23,
    7215 => 23,
    7216 => 23,
    7217 => 23,
    7218 => 23,
    7219 => 23,
    7220 => 23,
    7221 => 23,
    7222 => 23,
    7223 => 23,
    7224 => 23,
    7225 => 23,
    7226 => 23,
    7227 => 23,
    7228 => 23,
    7229 => 23,
    7230 => 23,
    7231 => 23,
    7232 => 23,
    7233 => 23,
    7234 => 23,
    7235 => 23,
    7236 => 23,
    7237 => 23,
    7238 => 23,
    7239 => 23,
    7240 => 22,
    7241 => 22,
    7242 => 22,
    7243 => 22,
    7244 => 22,
    7245 => 22,
    7246 => 22,
    7247 => 22,
    7248 => 22,
    7249 => 22,
    7250 => 22,
    7251 => 22,
    7252 => 22,
    7253 => 22,
    7254 => 22,
    7255 => 22,
    7256 => 22,
    7257 => 22,
    7258 => 22,
    7259 => 22,
    7260 => 22,
    7261 => 22,
    7262 => 22,
    7263 => 22,
    7264 => 22,
    7265 => 22,
    7266 => 22,
    7267 => 22,
    7268 => 22,
    7269 => 22,
    7270 => 22,
    7271 => 22,
    7272 => 22,
    7273 => 22,
    7274 => 22,
    7275 => 22,
    7276 => 22,
    7277 => 22,
    7278 => 22,
    7279 => 22,
    7280 => 22,
    7281 => 22,
    7282 => 22,
    7283 => 22,
    7284 => 21,
    7285 => 21,
    7286 => 21,
    7287 => 21,
    7288 => 21,
    7289 => 21,
    7290 => 21,
    7291 => 21,
    7292 => 21,
    7293 => 21,
    7294 => 21,
    7295 => 21,
    7296 => 21,
    7297 => 21,
    7298 => 21,
    7299 => 21,
    7300 => 21,
    7301 => 21,
    7302 => 21,
    7303 => 21,
    7304 => 21,
    7305 => 21,
    7306 => 21,
    7307 => 21,
    7308 => 21,
    7309 => 21,
    7310 => 21,
    7311 => 21,
    7312 => 21,
    7313 => 21,
    7314 => 21,
    7315 => 21,
    7316 => 21,
    7317 => 21,
    7318 => 21,
    7319 => 21,
    7320 => 21,
    7321 => 21,
    7322 => 21,
    7323 => 21,
    7324 => 21,
    7325 => 21,
    7326 => 21,
    7327 => 21,
    7328 => 20,
    7329 => 20,
    7330 => 20,
    7331 => 20,
    7332 => 20,
    7333 => 20,
    7334 => 20,
    7335 => 20,
    7336 => 20,
    7337 => 20,
    7338 => 20,
    7339 => 20,
    7340 => 20,
    7341 => 20,
    7342 => 20,
    7343 => 20,
    7344 => 20,
    7345 => 20,
    7346 => 20,
    7347 => 20,
    7348 => 20,
    7349 => 20,
    7350 => 20,
    7351 => 20,
    7352 => 20,
    7353 => 20,
    7354 => 20,
    7355 => 20,
    7356 => 20,
    7357 => 20,
    7358 => 20,
    7359 => 20,
    7360 => 20,
    7361 => 20,
    7362 => 20,
    7363 => 20,
    7364 => 20,
    7365 => 20,
    7366 => 20,
    7367 => 20,
    7368 => 20,
    7369 => 20,
    7370 => 20,
    7371 => 20,
    7372 => 19,
    7373 => 19,
    7374 => 19,
    7375 => 19,
    7376 => 19,
    7377 => 19,
    7378 => 19,
    7379 => 19,
    7380 => 19,
    7381 => 19,
    7382 => 19,
    7383 => 19,
    7384 => 19,
    7385 => 19,
    7386 => 19,
    7387 => 19,
    7388 => 19,
    7389 => 19,
    7390 => 19,
    7391 => 19,
    7392 => 19,
    7393 => 19,
    7394 => 19,
    7395 => 19,
    7396 => 19,
    7397 => 19,
    7398 => 19,
    7399 => 19,
    7400 => 19,
    7401 => 19,
    7402 => 19,
    7403 => 19,
    7404 => 19,
    7405 => 19,
    7406 => 19,
    7407 => 19,
    7408 => 19,
    7409 => 19,
    7410 => 19,
    7411 => 19,
    7412 => 19,
    7413 => 19,
    7414 => 19,
    7415 => 18,
    7416 => 18,
    7417 => 18,
    7418 => 18,
    7419 => 18,
    7420 => 18,
    7421 => 18,
    7422 => 18,
    7423 => 18,
    7424 => 18,
    7425 => 18,
    7426 => 18,
    7427 => 18,
    7428 => 18,
    7429 => 18,
    7430 => 18,
    7431 => 18,
    7432 => 18,
    7433 => 18,
    7434 => 18,
    7435 => 18,
    7436 => 18,
    7437 => 18,
    7438 => 18,
    7439 => 18,
    7440 => 18,
    7441 => 18,
    7442 => 18,
    7443 => 18,
    7444 => 18,
    7445 => 18,
    7446 => 18,
    7447 => 18,
    7448 => 18,
    7449 => 18,
    7450 => 18,
    7451 => 18,
    7452 => 18,
    7453 => 18,
    7454 => 18,
    7455 => 18,
    7456 => 18,
    7457 => 18,
    7458 => 18,
    7459 => 17,
    7460 => 17,
    7461 => 17,
    7462 => 17,
    7463 => 17,
    7464 => 17,
    7465 => 17,
    7466 => 17,
    7467 => 17,
    7468 => 17,
    7469 => 17,
    7470 => 17,
    7471 => 17,
    7472 => 17,
    7473 => 17,
    7474 => 17,
    7475 => 17,
    7476 => 17,
    7477 => 17,
    7478 => 17,
    7479 => 17,
    7480 => 17,
    7481 => 17,
    7482 => 17,
    7483 => 17,
    7484 => 17,
    7485 => 17,
    7486 => 17,
    7487 => 17,
    7488 => 17,
    7489 => 17,
    7490 => 17,
    7491 => 17,
    7492 => 17,
    7493 => 17,
    7494 => 17,
    7495 => 17,
    7496 => 17,
    7497 => 17,
    7498 => 17,
    7499 => 17,
    7500 => 17,
    7501 => 16,
    7502 => 16,
    7503 => 16,
    7504 => 16,
    7505 => 16,
    7506 => 16,
    7507 => 16,
    7508 => 16,
    7509 => 16,
    7510 => 16,
    7511 => 16,
    7512 => 16,
    7513 => 16,
    7514 => 16,
    7515 => 16,
    7516 => 16,
    7517 => 16,
    7518 => 16,
    7519 => 16,
    7520 => 16,
    7521 => 16,
    7522 => 16,
    7523 => 16,
    7524 => 16,
    7525 => 16,
    7526 => 16,
    7527 => 16,
    7528 => 16,
    7529 => 16,
    7530 => 16,
    7531 => 16,
    7532 => 16,
    7533 => 16,
    7534 => 16,
    7535 => 16,
    7536 => 16,
    7537 => 16,
    7538 => 16,
    7539 => 16,
    7540 => 16,
    7541 => 16,
    7542 => 16,
    7543 => 16,
    7544 => 15,
    7545 => 15,
    7546 => 15,
    7547 => 15,
    7548 => 15,
    7549 => 15,
    7550 => 15,
    7551 => 15,
    7552 => 15,
    7553 => 15,
    7554 => 15,
    7555 => 15,
    7556 => 15,
    7557 => 15,
    7558 => 15,
    7559 => 15,
    7560 => 15,
    7561 => 15,
    7562 => 15,
    7563 => 15,
    7564 => 15,
    7565 => 15,
    7566 => 15,
    7567 => 15,
    7568 => 15,
    7569 => 15,
    7570 => 15,
    7571 => 15,
    7572 => 15,
    7573 => 15,
    7574 => 15,
    7575 => 15,
    7576 => 15,
    7577 => 15,
    7578 => 15,
    7579 => 15,
    7580 => 15,
    7581 => 15,
    7582 => 15,
    7583 => 15,
    7584 => 15,
    7585 => 15,
    7586 => 15,
    7587 => 14,
    7588 => 14,
    7589 => 14,
    7590 => 14,
    7591 => 14,
    7592 => 14,
    7593 => 14,
    7594 => 14,
    7595 => 14,
    7596 => 14,
    7597 => 14,
    7598 => 14,
    7599 => 14,
    7600 => 14,
    7601 => 14,
    7602 => 14,
    7603 => 14,
    7604 => 14,
    7605 => 14,
    7606 => 14,
    7607 => 14,
    7608 => 14,
    7609 => 14,
    7610 => 14,
    7611 => 14,
    7612 => 14,
    7613 => 14,
    7614 => 14,
    7615 => 14,
    7616 => 14,
    7617 => 14,
    7618 => 14,
    7619 => 14,
    7620 => 14,
    7621 => 14,
    7622 => 14,
    7623 => 14,
    7624 => 14,
    7625 => 14,
    7626 => 14,
    7627 => 14,
    7628 => 14,
    7629 => 13,
    7630 => 13,
    7631 => 13,
    7632 => 13,
    7633 => 13,
    7634 => 13,
    7635 => 13,
    7636 => 13,
    7637 => 13,
    7638 => 13,
    7639 => 13,
    7640 => 13,
    7641 => 13,
    7642 => 13,
    7643 => 13,
    7644 => 13,
    7645 => 13,
    7646 => 13,
    7647 => 13,
    7648 => 13,
    7649 => 13,
    7650 => 13,
    7651 => 13,
    7652 => 13,
    7653 => 13,
    7654 => 13,
    7655 => 13,
    7656 => 13,
    7657 => 13,
    7658 => 13,
    7659 => 13,
    7660 => 13,
    7661 => 13,
    7662 => 13,
    7663 => 13,
    7664 => 13,
    7665 => 13,
    7666 => 13,
    7667 => 13,
    7668 => 13,
    7669 => 13,
    7670 => 13,
    7671 => 13,
    7672 => 12,
    7673 => 12,
    7674 => 12,
    7675 => 12,
    7676 => 12,
    7677 => 12,
    7678 => 12,
    7679 => 12,
    7680 => 12,
    7681 => 12,
    7682 => 12,
    7683 => 12,
    7684 => 12,
    7685 => 12,
    7686 => 12,
    7687 => 12,
    7688 => 12,
    7689 => 12,
    7690 => 12,
    7691 => 12,
    7692 => 12,
    7693 => 12,
    7694 => 12,
    7695 => 12,
    7696 => 12,
    7697 => 12,
    7698 => 12,
    7699 => 12,
    7700 => 12,
    7701 => 12,
    7702 => 12,
    7703 => 12,
    7704 => 12,
    7705 => 12,
    7706 => 12,
    7707 => 12,
    7708 => 12,
    7709 => 12,
    7710 => 12,
    7711 => 12,
    7712 => 12,
    7713 => 12,
    7714 => 11,
    7715 => 11,
    7716 => 11,
    7717 => 11,
    7718 => 11,
    7719 => 11,
    7720 => 11,
    7721 => 11,
    7722 => 11,
    7723 => 11,
    7724 => 11,
    7725 => 11,
    7726 => 11,
    7727 => 11,
    7728 => 11,
    7729 => 11,
    7730 => 11,
    7731 => 11,
    7732 => 11,
    7733 => 11,
    7734 => 11,
    7735 => 11,
    7736 => 11,
    7737 => 11,
    7738 => 11,
    7739 => 11,
    7740 => 11,
    7741 => 11,
    7742 => 11,
    7743 => 11,
    7744 => 11,
    7745 => 11,
    7746 => 11,
    7747 => 11,
    7748 => 11,
    7749 => 11,
    7750 => 11,
    7751 => 11,
    7752 => 11,
    7753 => 11,
    7754 => 11,
    7755 => 11,
    7756 => 10,
    7757 => 10,
    7758 => 10,
    7759 => 10,
    7760 => 10,
    7761 => 10,
    7762 => 10,
    7763 => 10,
    7764 => 10,
    7765 => 10,
    7766 => 10,
    7767 => 10,
    7768 => 10,
    7769 => 10,
    7770 => 10,
    7771 => 10,
    7772 => 10,
    7773 => 10,
    7774 => 10,
    7775 => 10,
    7776 => 10,
    7777 => 10,
    7778 => 10,
    7779 => 10,
    7780 => 10,
    7781 => 10,
    7782 => 10,
    7783 => 10,
    7784 => 10,
    7785 => 10,
    7786 => 10,
    7787 => 10,
    7788 => 10,
    7789 => 10,
    7790 => 10,
    7791 => 10,
    7792 => 10,
    7793 => 10,
    7794 => 10,
    7795 => 10,
    7796 => 10,
    7797 => 10,
    7798 => 9,
    7799 => 9,
    7800 => 9,
    7801 => 9,
    7802 => 9,
    7803 => 9,
    7804 => 9,
    7805 => 9,
    7806 => 9,
    7807 => 9,
    7808 => 9,
    7809 => 9,
    7810 => 9,
    7811 => 9,
    7812 => 9,
    7813 => 9,
    7814 => 9,
    7815 => 9,
    7816 => 9,
    7817 => 9,
    7818 => 9,
    7819 => 9,
    7820 => 9,
    7821 => 9,
    7822 => 9,
    7823 => 9,
    7824 => 9,
    7825 => 9,
    7826 => 9,
    7827 => 9,
    7828 => 9,
    7829 => 9,
    7830 => 9,
    7831 => 9,
    7832 => 9,
    7833 => 9,
    7834 => 9,
    7835 => 9,
    7836 => 9,
    7837 => 9,
    7838 => 9,
    7839 => 9,
    7840 => 8,
    7841 => 8,
    7842 => 8,
    7843 => 8,
    7844 => 8,
    7845 => 8,
    7846 => 8,
    7847 => 8,
    7848 => 8,
    7849 => 8,
    7850 => 8,
    7851 => 8,
    7852 => 8,
    7853 => 8,
    7854 => 8,
    7855 => 8,
    7856 => 8,
    7857 => 8,
    7858 => 8,
    7859 => 8,
    7860 => 8,
    7861 => 8,
    7862 => 8,
    7863 => 8,
    7864 => 8,
    7865 => 8,
    7866 => 8,
    7867 => 8,
    7868 => 8,
    7869 => 8,
    7870 => 8,
    7871 => 8,
    7872 => 8,
    7873 => 8,
    7874 => 8,
    7875 => 8,
    7876 => 8,
    7877 => 8,
    7878 => 8,
    7879 => 8,
    7880 => 8,
    7881 => 7,
    7882 => 7,
    7883 => 7,
    7884 => 7,
    7885 => 7,
    7886 => 7,
    7887 => 7,
    7888 => 7,
    7889 => 7,
    7890 => 7,
    7891 => 7,
    7892 => 7,
    7893 => 7,
    7894 => 7,
    7895 => 7,
    7896 => 7,
    7897 => 7,
    7898 => 7,
    7899 => 7,
    7900 => 7,
    7901 => 7,
    7902 => 7,
    7903 => 7,
    7904 => 7,
    7905 => 7,
    7906 => 7,
    7907 => 7,
    7908 => 7,
    7909 => 7,
    7910 => 7,
    7911 => 7,
    7912 => 7,
    7913 => 7,
    7914 => 7,
    7915 => 7,
    7916 => 7,
    7917 => 7,
    7918 => 7,
    7919 => 7,
    7920 => 7,
    7921 => 7,
    7922 => 7,
    7923 => 6,
    7924 => 6,
    7925 => 6,
    7926 => 6,
    7927 => 6,
    7928 => 6,
    7929 => 6,
    7930 => 6,
    7931 => 6,
    7932 => 6,
    7933 => 6,
    7934 => 6,
    7935 => 6,
    7936 => 6,
    7937 => 6,
    7938 => 6,
    7939 => 6,
    7940 => 6,
    7941 => 6,
    7942 => 6,
    7943 => 6,
    7944 => 6,
    7945 => 6,
    7946 => 6,
    7947 => 6,
    7948 => 6,
    7949 => 6,
    7950 => 6,
    7951 => 6,
    7952 => 6,
    7953 => 6,
    7954 => 6,
    7955 => 6,
    7956 => 6,
    7957 => 6,
    7958 => 6,
    7959 => 6,
    7960 => 6,
    7961 => 6,
    7962 => 6,
    7963 => 6,
    7964 => 6,
    7965 => 5,
    7966 => 5,
    7967 => 5,
    7968 => 5,
    7969 => 5,
    7970 => 5,
    7971 => 5,
    7972 => 5,
    7973 => 5,
    7974 => 5,
    7975 => 5,
    7976 => 5,
    7977 => 5,
    7978 => 5,
    7979 => 5,
    7980 => 5,
    7981 => 5,
    7982 => 5,
    7983 => 5,
    7984 => 5,
    7985 => 5,
    7986 => 5,
    7987 => 5,
    7988 => 5,
    7989 => 5,
    7990 => 5,
    7991 => 5,
    7992 => 5,
    7993 => 5,
    7994 => 5,
    7995 => 5,
    7996 => 5,
    7997 => 5,
    7998 => 5,
    7999 => 5,
    8000 => 5,
    8001 => 5,
    8002 => 5,
    8003 => 5,
    8004 => 5,
    8005 => 5,
    8006 => 4,
    8007 => 4,
    8008 => 4,
    8009 => 4,
    8010 => 4,
    8011 => 4,
    8012 => 4,
    8013 => 4,
    8014 => 4,
    8015 => 4,
    8016 => 4,
    8017 => 4,
    8018 => 4,
    8019 => 4,
    8020 => 4,
    8021 => 4,
    8022 => 4,
    8023 => 4,
    8024 => 4,
    8025 => 4,
    8026 => 4,
    8027 => 4,
    8028 => 4,
    8029 => 4,
    8030 => 4,
    8031 => 4,
    8032 => 4,
    8033 => 4,
    8034 => 4,
    8035 => 4,
    8036 => 4,
    8037 => 4,
    8038 => 4,
    8039 => 4,
    8040 => 4,
    8041 => 4,
    8042 => 4,
    8043 => 4,
    8044 => 4,
    8045 => 4,
    8046 => 4,
    8047 => 4,
    8048 => 3,
    8049 => 3,
    8050 => 3,
    8051 => 3,
    8052 => 3,
    8053 => 3,
    8054 => 3,
    8055 => 3,
    8056 => 3,
    8057 => 3,
    8058 => 3,
    8059 => 3,
    8060 => 3,
    8061 => 3,
    8062 => 3,
    8063 => 3,
    8064 => 3,
    8065 => 3,
    8066 => 3,
    8067 => 3,
    8068 => 3,
    8069 => 3,
    8070 => 3,
    8071 => 3,
    8072 => 3,
    8073 => 3,
    8074 => 3,
    8075 => 3,
    8076 => 3,
    8077 => 3,
    8078 => 3,
    8079 => 3,
    8080 => 3,
    8081 => 3,
    8082 => 3,
    8083 => 3,
    8084 => 3,
    8085 => 3,
    8086 => 3,
    8087 => 3,
    8088 => 3,
    8089 => 2,
    8090 => 2,
    8091 => 2,
    8092 => 2,
    8093 => 2,
    8094 => 2,
    8095 => 2,
    8096 => 2,
    8097 => 2,
    8098 => 2,
    8099 => 2,
    8100 => 2,
    8101 => 2,
    8102 => 2,
    8103 => 2,
    8104 => 2,
    8105 => 2,
    8106 => 2,
    8107 => 2,
    8108 => 2,
    8109 => 2,
    8110 => 2,
    8111 => 2,
    8112 => 2,
    8113 => 2,
    8114 => 2,
    8115 => 2,
    8116 => 2,
    8117 => 2,
    8118 => 2,
    8119 => 2,
    8120 => 2,
    8121 => 2,
    8122 => 2,
    8123 => 2,
    8124 => 2,
    8125 => 2,
    8126 => 2,
    8127 => 2,
    8128 => 2,
    8129 => 2,
    8130 => 1,
    8131 => 1,
    8132 => 1,
    8133 => 1,
    8134 => 1,
    8135 => 1,
    8136 => 1,
    8137 => 1,
    8138 => 1,
    8139 => 1,
    8140 => 1,
    8141 => 1,
    8142 => 1,
    8143 => 1,
    8144 => 1,
    8145 => 1,
    8146 => 1,
    8147 => 1,
    8148 => 1,
    8149 => 1,
    8150 => 1,
    8151 => 1,
    8152 => 1,
    8153 => 1,
    8154 => 1,
    8155 => 1,
    8156 => 1,
    8157 => 1,
    8158 => 1,
    8159 => 1,
    8160 => 1,
    8161 => 1,
    8162 => 1,
    8163 => 1,
    8164 => 1,
    8165 => 1,
    8166 => 1,
    8167 => 1,
    8168 => 1,
    8169 => 1,
    8170 => 1,
    8171 => 1,
    8172 => 0,
    8173 => 0,
    8174 => 0,
    8175 => 0,
    8176 => 0,
    8177 => 0,
    8178 => 0,
    8179 => 0,
    8180 => 0,
    8181 => 0,
    8182 => 0,
    8183 => 0,
    8184 => 0,
    8185 => 0,
    8186 => 0,
    8187 => 0,
    8188 => 0,
    8189 => 0,
    8190 => 0,
    8191 => 0,
    8192 => 0,
    8193 => 0,
    8194 => 0,
    8195 => 0,
    8196 => 0,
    8197 => 0,
    8198 => 0,
    8199 => 0,
    8200 => 0,
    8201 => 0,
    8202 => 0,
    8203 => 0,
    8204 => 0,
    8205 => 0,
    8206 => 0,
    8207 => 0,
    8208 => 0,
    8209 => 0,
    8210 => 0,
    8211 => 0,
    8212 => 0,
    8213 => -1,
    8214 => -1,
    8215 => -1,
    8216 => -1,
    8217 => -1,
    8218 => -1,
    8219 => -1,
    8220 => -1,
    8221 => -1,
    8222 => -1,
    8223 => -1,
    8224 => -1,
    8225 => -1,
    8226 => -1,
    8227 => -1,
    8228 => -1,
    8229 => -1,
    8230 => -1,
    8231 => -1,
    8232 => -1,
    8233 => -1,
    8234 => -1,
    8235 => -1,
    8236 => -1,
    8237 => -1,
    8238 => -1,
    8239 => -1,
    8240 => -1,
    8241 => -1,
    8242 => -1,
    8243 => -1,
    8244 => -1,
    8245 => -1,
    8246 => -1,
    8247 => -1,
    8248 => -1,
    8249 => -1,
    8250 => -1,
    8251 => -1,
    8252 => -1,
    8253 => -1,
    8254 => -1,
    8255 => -2,
    8256 => -2,
    8257 => -2,
    8258 => -2,
    8259 => -2,
    8260 => -2,
    8261 => -2,
    8262 => -2,
    8263 => -2,
    8264 => -2,
    8265 => -2,
    8266 => -2,
    8267 => -2,
    8268 => -2,
    8269 => -2,
    8270 => -2,
    8271 => -2,
    8272 => -2,
    8273 => -2,
    8274 => -2,
    8275 => -2,
    8276 => -2,
    8277 => -2,
    8278 => -2,
    8279 => -2,
    8280 => -2,
    8281 => -2,
    8282 => -2,
    8283 => -2,
    8284 => -2,
    8285 => -2,
    8286 => -2,
    8287 => -2,
    8288 => -2,
    8289 => -2,
    8290 => -2,
    8291 => -2,
    8292 => -2,
    8293 => -2,
    8294 => -2,
    8295 => -2,
    8296 => -3,
    8297 => -3,
    8298 => -3,
    8299 => -3,
    8300 => -3,
    8301 => -3,
    8302 => -3,
    8303 => -3,
    8304 => -3,
    8305 => -3,
    8306 => -3,
    8307 => -3,
    8308 => -3,
    8309 => -3,
    8310 => -3,
    8311 => -3,
    8312 => -3,
    8313 => -3,
    8314 => -3,
    8315 => -3,
    8316 => -3,
    8317 => -3,
    8318 => -3,
    8319 => -3,
    8320 => -3,
    8321 => -3,
    8322 => -3,
    8323 => -3,
    8324 => -3,
    8325 => -3,
    8326 => -3,
    8327 => -3,
    8328 => -3,
    8329 => -3,
    8330 => -3,
    8331 => -3,
    8332 => -3,
    8333 => -3,
    8334 => -3,
    8335 => -3,
    8336 => -3,
    8337 => -4,
    8338 => -4,
    8339 => -4,
    8340 => -4,
    8341 => -4,
    8342 => -4,
    8343 => -4,
    8344 => -4,
    8345 => -4,
    8346 => -4,
    8347 => -4,
    8348 => -4,
    8349 => -4,
    8350 => -4,
    8351 => -4,
    8352 => -4,
    8353 => -4,
    8354 => -4,
    8355 => -4,
    8356 => -4,
    8357 => -4,
    8358 => -4,
    8359 => -4,
    8360 => -4,
    8361 => -4,
    8362 => -4,
    8363 => -4,
    8364 => -4,
    8365 => -4,
    8366 => -4,
    8367 => -4,
    8368 => -4,
    8369 => -4,
    8370 => -4,
    8371 => -4,
    8372 => -4,
    8373 => -4,
    8374 => -4,
    8375 => -4,
    8376 => -4,
    8377 => -4,
    8378 => -4,
    8379 => -5,
    8380 => -5,
    8381 => -5,
    8382 => -5,
    8383 => -5,
    8384 => -5,
    8385 => -5,
    8386 => -5,
    8387 => -5,
    8388 => -5,
    8389 => -5,
    8390 => -5,
    8391 => -5,
    8392 => -5,
    8393 => -5,
    8394 => -5,
    8395 => -5,
    8396 => -5,
    8397 => -5,
    8398 => -5,
    8399 => -5,
    8400 => -5,
    8401 => -5,
    8402 => -5,
    8403 => -5,
    8404 => -5,
    8405 => -5,
    8406 => -5,
    8407 => -5,
    8408 => -5,
    8409 => -5,
    8410 => -5,
    8411 => -5,
    8412 => -5,
    8413 => -5,
    8414 => -5,
    8415 => -5,
    8416 => -5,
    8417 => -5,
    8418 => -5,
    8419 => -5,
    8420 => -6,
    8421 => -6,
    8422 => -6,
    8423 => -6,
    8424 => -6,
    8425 => -6,
    8426 => -6,
    8427 => -6,
    8428 => -6,
    8429 => -6,
    8430 => -6,
    8431 => -6,
    8432 => -6,
    8433 => -6,
    8434 => -6,
    8435 => -6,
    8436 => -6,
    8437 => -6,
    8438 => -6,
    8439 => -6,
    8440 => -6,
    8441 => -6,
    8442 => -6,
    8443 => -6,
    8444 => -6,
    8445 => -6,
    8446 => -6,
    8447 => -6,
    8448 => -6,
    8449 => -6,
    8450 => -6,
    8451 => -6,
    8452 => -6,
    8453 => -6,
    8454 => -6,
    8455 => -6,
    8456 => -6,
    8457 => -6,
    8458 => -6,
    8459 => -6,
    8460 => -6,
    8461 => -6,
    8462 => -7,
    8463 => -7,
    8464 => -7,
    8465 => -7,
    8466 => -7,
    8467 => -7,
    8468 => -7,
    8469 => -7,
    8470 => -7,
    8471 => -7,
    8472 => -7,
    8473 => -7,
    8474 => -7,
    8475 => -7,
    8476 => -7,
    8477 => -7,
    8478 => -7,
    8479 => -7,
    8480 => -7,
    8481 => -7,
    8482 => -7,
    8483 => -7,
    8484 => -7,
    8485 => -7,
    8486 => -7,
    8487 => -7,
    8488 => -7,
    8489 => -7,
    8490 => -7,
    8491 => -7,
    8492 => -7,
    8493 => -7,
    8494 => -7,
    8495 => -7,
    8496 => -7,
    8497 => -7,
    8498 => -7,
    8499 => -7,
    8500 => -7,
    8501 => -7,
    8502 => -7,
    8503 => -7,
    8504 => -8,
    8505 => -8,
    8506 => -8,
    8507 => -8,
    8508 => -8,
    8509 => -8,
    8510 => -8,
    8511 => -8,
    8512 => -8,
    8513 => -8,
    8514 => -8,
    8515 => -8,
    8516 => -8,
    8517 => -8,
    8518 => -8,
    8519 => -8,
    8520 => -8,
    8521 => -8,
    8522 => -8,
    8523 => -8,
    8524 => -8,
    8525 => -8,
    8526 => -8,
    8527 => -8,
    8528 => -8,
    8529 => -8,
    8530 => -8,
    8531 => -8,
    8532 => -8,
    8533 => -8,
    8534 => -8,
    8535 => -8,
    8536 => -8,
    8537 => -8,
    8538 => -8,
    8539 => -8,
    8540 => -8,
    8541 => -8,
    8542 => -8,
    8543 => -8,
    8544 => -8,
    8545 => -9,
    8546 => -9,
    8547 => -9,
    8548 => -9,
    8549 => -9,
    8550 => -9,
    8551 => -9,
    8552 => -9,
    8553 => -9,
    8554 => -9,
    8555 => -9,
    8556 => -9,
    8557 => -9,
    8558 => -9,
    8559 => -9,
    8560 => -9,
    8561 => -9,
    8562 => -9,
    8563 => -9,
    8564 => -9,
    8565 => -9,
    8566 => -9,
    8567 => -9,
    8568 => -9,
    8569 => -9,
    8570 => -9,
    8571 => -9,
    8572 => -9,
    8573 => -9,
    8574 => -9,
    8575 => -9,
    8576 => -9,
    8577 => -9,
    8578 => -9,
    8579 => -9,
    8580 => -9,
    8581 => -9,
    8582 => -9,
    8583 => -9,
    8584 => -9,
    8585 => -9,
    8586 => -9,
    8587 => -10,
    8588 => -10,
    8589 => -10,
    8590 => -10,
    8591 => -10,
    8592 => -10,
    8593 => -10,
    8594 => -10,
    8595 => -10,
    8596 => -10,
    8597 => -10,
    8598 => -10,
    8599 => -10,
    8600 => -10,
    8601 => -10,
    8602 => -10,
    8603 => -10,
    8604 => -10,
    8605 => -10,
    8606 => -10,
    8607 => -10,
    8608 => -10,
    8609 => -10,
    8610 => -10,
    8611 => -10,
    8612 => -10,
    8613 => -10,
    8614 => -10,
    8615 => -10,
    8616 => -10,
    8617 => -10,
    8618 => -10,
    8619 => -10,
    8620 => -10,
    8621 => -10,
    8622 => -10,
    8623 => -10,
    8624 => -10,
    8625 => -10,
    8626 => -10,
    8627 => -10,
    8628 => -10,
    8629 => -11,
    8630 => -11,
    8631 => -11,
    8632 => -11,
    8633 => -11,
    8634 => -11,
    8635 => -11,
    8636 => -11,
    8637 => -11,
    8638 => -11,
    8639 => -11,
    8640 => -11,
    8641 => -11,
    8642 => -11,
    8643 => -11,
    8644 => -11,
    8645 => -11,
    8646 => -11,
    8647 => -11,
    8648 => -11,
    8649 => -11,
    8650 => -11,
    8651 => -11,
    8652 => -11,
    8653 => -11,
    8654 => -11,
    8655 => -11,
    8656 => -11,
    8657 => -11,
    8658 => -11,
    8659 => -11,
    8660 => -11,
    8661 => -11,
    8662 => -11,
    8663 => -11,
    8664 => -11,
    8665 => -11,
    8666 => -11,
    8667 => -11,
    8668 => -11,
    8669 => -11,
    8670 => -11,
    8671 => -12,
    8672 => -12,
    8673 => -12,
    8674 => -12,
    8675 => -12,
    8676 => -12,
    8677 => -12,
    8678 => -12,
    8679 => -12,
    8680 => -12,
    8681 => -12,
    8682 => -12,
    8683 => -12,
    8684 => -12,
    8685 => -12,
    8686 => -12,
    8687 => -12,
    8688 => -12,
    8689 => -12,
    8690 => -12,
    8691 => -12,
    8692 => -12,
    8693 => -12,
    8694 => -12,
    8695 => -12,
    8696 => -12,
    8697 => -12,
    8698 => -12,
    8699 => -12,
    8700 => -12,
    8701 => -12,
    8702 => -12,
    8703 => -12,
    8704 => -12,
    8705 => -12,
    8706 => -12,
    8707 => -12,
    8708 => -12,
    8709 => -12,
    8710 => -12,
    8711 => -12,
    8712 => -12,
    8713 => -13,
    8714 => -13,
    8715 => -13,
    8716 => -13,
    8717 => -13,
    8718 => -13,
    8719 => -13,
    8720 => -13,
    8721 => -13,
    8722 => -13,
    8723 => -13,
    8724 => -13,
    8725 => -13,
    8726 => -13,
    8727 => -13,
    8728 => -13,
    8729 => -13,
    8730 => -13,
    8731 => -13,
    8732 => -13,
    8733 => -13,
    8734 => -13,
    8735 => -13,
    8736 => -13,
    8737 => -13,
    8738 => -13,
    8739 => -13,
    8740 => -13,
    8741 => -13,
    8742 => -13,
    8743 => -13,
    8744 => -13,
    8745 => -13,
    8746 => -13,
    8747 => -13,
    8748 => -13,
    8749 => -13,
    8750 => -13,
    8751 => -13,
    8752 => -13,
    8753 => -13,
    8754 => -13,
    8755 => -13,
    8756 => -14,
    8757 => -14,
    8758 => -14,
    8759 => -14,
    8760 => -14,
    8761 => -14,
    8762 => -14,
    8763 => -14,
    8764 => -14,
    8765 => -14,
    8766 => -14,
    8767 => -14,
    8768 => -14,
    8769 => -14,
    8770 => -14,
    8771 => -14,
    8772 => -14,
    8773 => -14,
    8774 => -14,
    8775 => -14,
    8776 => -14,
    8777 => -14,
    8778 => -14,
    8779 => -14,
    8780 => -14,
    8781 => -14,
    8782 => -14,
    8783 => -14,
    8784 => -14,
    8785 => -14,
    8786 => -14,
    8787 => -14,
    8788 => -14,
    8789 => -14,
    8790 => -14,
    8791 => -14,
    8792 => -14,
    8793 => -14,
    8794 => -14,
    8795 => -14,
    8796 => -14,
    8797 => -14,
    8798 => -15,
    8799 => -15,
    8800 => -15,
    8801 => -15,
    8802 => -15,
    8803 => -15,
    8804 => -15,
    8805 => -15,
    8806 => -15,
    8807 => -15,
    8808 => -15,
    8809 => -15,
    8810 => -15,
    8811 => -15,
    8812 => -15,
    8813 => -15,
    8814 => -15,
    8815 => -15,
    8816 => -15,
    8817 => -15,
    8818 => -15,
    8819 => -15,
    8820 => -15,
    8821 => -15,
    8822 => -15,
    8823 => -15,
    8824 => -15,
    8825 => -15,
    8826 => -15,
    8827 => -15,
    8828 => -15,
    8829 => -15,
    8830 => -15,
    8831 => -15,
    8832 => -15,
    8833 => -15,
    8834 => -15,
    8835 => -15,
    8836 => -15,
    8837 => -15,
    8838 => -15,
    8839 => -15,
    8840 => -15,
    8841 => -16,
    8842 => -16,
    8843 => -16,
    8844 => -16,
    8845 => -16,
    8846 => -16,
    8847 => -16,
    8848 => -16,
    8849 => -16,
    8850 => -16,
    8851 => -16,
    8852 => -16,
    8853 => -16,
    8854 => -16,
    8855 => -16,
    8856 => -16,
    8857 => -16,
    8858 => -16,
    8859 => -16,
    8860 => -16,
    8861 => -16,
    8862 => -16,
    8863 => -16,
    8864 => -16,
    8865 => -16,
    8866 => -16,
    8867 => -16,
    8868 => -16,
    8869 => -16,
    8870 => -16,
    8871 => -16,
    8872 => -16,
    8873 => -16,
    8874 => -16,
    8875 => -16,
    8876 => -16,
    8877 => -16,
    8878 => -16,
    8879 => -16,
    8880 => -16,
    8881 => -16,
    8882 => -16,
    8883 => -16,
    8884 => -17,
    8885 => -17,
    8886 => -17,
    8887 => -17,
    8888 => -17,
    8889 => -17,
    8890 => -17,
    8891 => -17,
    8892 => -17,
    8893 => -17,
    8894 => -17,
    8895 => -17,
    8896 => -17,
    8897 => -17,
    8898 => -17,
    8899 => -17,
    8900 => -17,
    8901 => -17,
    8902 => -17,
    8903 => -17,
    8904 => -17,
    8905 => -17,
    8906 => -17,
    8907 => -17,
    8908 => -17,
    8909 => -17,
    8910 => -17,
    8911 => -17,
    8912 => -17,
    8913 => -17,
    8914 => -17,
    8915 => -17,
    8916 => -17,
    8917 => -17,
    8918 => -17,
    8919 => -17,
    8920 => -17,
    8921 => -17,
    8922 => -17,
    8923 => -17,
    8924 => -17,
    8925 => -17,
    8926 => -18,
    8927 => -18,
    8928 => -18,
    8929 => -18,
    8930 => -18,
    8931 => -18,
    8932 => -18,
    8933 => -18,
    8934 => -18,
    8935 => -18,
    8936 => -18,
    8937 => -18,
    8938 => -18,
    8939 => -18,
    8940 => -18,
    8941 => -18,
    8942 => -18,
    8943 => -18,
    8944 => -18,
    8945 => -18,
    8946 => -18,
    8947 => -18,
    8948 => -18,
    8949 => -18,
    8950 => -18,
    8951 => -18,
    8952 => -18,
    8953 => -18,
    8954 => -18,
    8955 => -18,
    8956 => -18,
    8957 => -18,
    8958 => -18,
    8959 => -18,
    8960 => -18,
    8961 => -18,
    8962 => -18,
    8963 => -18,
    8964 => -18,
    8965 => -18,
    8966 => -18,
    8967 => -18,
    8968 => -18,
    8969 => -18,
    8970 => -19,
    8971 => -19,
    8972 => -19,
    8973 => -19,
    8974 => -19,
    8975 => -19,
    8976 => -19,
    8977 => -19,
    8978 => -19,
    8979 => -19,
    8980 => -19,
    8981 => -19,
    8982 => -19,
    8983 => -19,
    8984 => -19,
    8985 => -19,
    8986 => -19,
    8987 => -19,
    8988 => -19,
    8989 => -19,
    8990 => -19,
    8991 => -19,
    8992 => -19,
    8993 => -19,
    8994 => -19,
    8995 => -19,
    8996 => -19,
    8997 => -19,
    8998 => -19,
    8999 => -19,
    9000 => -19,
    9001 => -19,
    9002 => -19,
    9003 => -19,
    9004 => -19,
    9005 => -19,
    9006 => -19,
    9007 => -19,
    9008 => -19,
    9009 => -19,
    9010 => -19,
    9011 => -19,
    9012 => -19,
    9013 => -20,
    9014 => -20,
    9015 => -20,
    9016 => -20,
    9017 => -20,
    9018 => -20,
    9019 => -20,
    9020 => -20,
    9021 => -20,
    9022 => -20,
    9023 => -20,
    9024 => -20,
    9025 => -20,
    9026 => -20,
    9027 => -20,
    9028 => -20,
    9029 => -20,
    9030 => -20,
    9031 => -20,
    9032 => -20,
    9033 => -20,
    9034 => -20,
    9035 => -20,
    9036 => -20,
    9037 => -20,
    9038 => -20,
    9039 => -20,
    9040 => -20,
    9041 => -20,
    9042 => -20,
    9043 => -20,
    9044 => -20,
    9045 => -20,
    9046 => -20,
    9047 => -20,
    9048 => -20,
    9049 => -20,
    9050 => -20,
    9051 => -20,
    9052 => -20,
    9053 => -20,
    9054 => -20,
    9055 => -20,
    9056 => -20,
    9057 => -21,
    9058 => -21,
    9059 => -21,
    9060 => -21,
    9061 => -21,
    9062 => -21,
    9063 => -21,
    9064 => -21,
    9065 => -21,
    9066 => -21,
    9067 => -21,
    9068 => -21,
    9069 => -21,
    9070 => -21,
    9071 => -21,
    9072 => -21,
    9073 => -21,
    9074 => -21,
    9075 => -21,
    9076 => -21,
    9077 => -21,
    9078 => -21,
    9079 => -21,
    9080 => -21,
    9081 => -21,
    9082 => -21,
    9083 => -21,
    9084 => -21,
    9085 => -21,
    9086 => -21,
    9087 => -21,
    9088 => -21,
    9089 => -21,
    9090 => -21,
    9091 => -21,
    9092 => -21,
    9093 => -21,
    9094 => -21,
    9095 => -21,
    9096 => -21,
    9097 => -21,
    9098 => -21,
    9099 => -21,
    9100 => -21,
    9101 => -22,
    9102 => -22,
    9103 => -22,
    9104 => -22,
    9105 => -22,
    9106 => -22,
    9107 => -22,
    9108 => -22,
    9109 => -22,
    9110 => -22,
    9111 => -22,
    9112 => -22,
    9113 => -22,
    9114 => -22,
    9115 => -22,
    9116 => -22,
    9117 => -22,
    9118 => -22,
    9119 => -22,
    9120 => -22,
    9121 => -22,
    9122 => -22,
    9123 => -22,
    9124 => -22,
    9125 => -22,
    9126 => -22,
    9127 => -22,
    9128 => -22,
    9129 => -22,
    9130 => -22,
    9131 => -22,
    9132 => -22,
    9133 => -22,
    9134 => -22,
    9135 => -22,
    9136 => -22,
    9137 => -22,
    9138 => -22,
    9139 => -22,
    9140 => -22,
    9141 => -22,
    9142 => -22,
    9143 => -22,
    9144 => -22,
    9145 => -23,
    9146 => -23,
    9147 => -23,
    9148 => -23,
    9149 => -23,
    9150 => -23,
    9151 => -23,
    9152 => -23,
    9153 => -23,
    9154 => -23,
    9155 => -23,
    9156 => -23,
    9157 => -23,
    9158 => -23,
    9159 => -23,
    9160 => -23,
    9161 => -23,
    9162 => -23,
    9163 => -23,
    9164 => -23,
    9165 => -23,
    9166 => -23,
    9167 => -23,
    9168 => -23,
    9169 => -23,
    9170 => -23,
    9171 => -23,
    9172 => -23,
    9173 => -23,
    9174 => -23,
    9175 => -23,
    9176 => -23,
    9177 => -23,
    9178 => -23,
    9179 => -23,
    9180 => -23,
    9181 => -23,
    9182 => -23,
    9183 => -23,
    9184 => -23,
    9185 => -23,
    9186 => -23,
    9187 => -23,
    9188 => -23,
    9189 => -24,
    9190 => -24,
    9191 => -24,
    9192 => -24,
    9193 => -24,
    9194 => -24,
    9195 => -24,
    9196 => -24,
    9197 => -24,
    9198 => -24,
    9199 => -24,
    9200 => -24,
    9201 => -24,
    9202 => -24,
    9203 => -24,
    9204 => -24,
    9205 => -24,
    9206 => -24,
    9207 => -24,
    9208 => -24,
    9209 => -24,
    9210 => -24,
    9211 => -24,
    9212 => -24,
    9213 => -24,
    9214 => -24,
    9215 => -24,
    9216 => -24,
    9217 => -24,
    9218 => -24,
    9219 => -24,
    9220 => -24,
    9221 => -24,
    9222 => -24,
    9223 => -24,
    9224 => -24,
    9225 => -24,
    9226 => -24,
    9227 => -24,
    9228 => -24,
    9229 => -24,
    9230 => -24,
    9231 => -24,
    9232 => -24,
    9233 => -24,
    9234 => -25,
    9235 => -25,
    9236 => -25,
    9237 => -25,
    9238 => -25,
    9239 => -25,
    9240 => -25,
    9241 => -25,
    9242 => -25,
    9243 => -25,
    9244 => -25,
    9245 => -25,
    9246 => -25,
    9247 => -25,
    9248 => -25,
    9249 => -25,
    9250 => -25,
    9251 => -25,
    9252 => -25,
    9253 => -25,
    9254 => -25,
    9255 => -25,
    9256 => -25,
    9257 => -25,
    9258 => -25,
    9259 => -25,
    9260 => -25,
    9261 => -25,
    9262 => -25,
    9263 => -25,
    9264 => -25,
    9265 => -25,
    9266 => -25,
    9267 => -25,
    9268 => -25,
    9269 => -25,
    9270 => -25,
    9271 => -25,
    9272 => -25,
    9273 => -25,
    9274 => -25,
    9275 => -25,
    9276 => -25,
    9277 => -25,
    9278 => -25,
    9279 => -26,
    9280 => -26,
    9281 => -26,
    9282 => -26,
    9283 => -26,
    9284 => -26,
    9285 => -26,
    9286 => -26,
    9287 => -26,
    9288 => -26,
    9289 => -26,
    9290 => -26,
    9291 => -26,
    9292 => -26,
    9293 => -26,
    9294 => -26,
    9295 => -26,
    9296 => -26,
    9297 => -26,
    9298 => -26,
    9299 => -26,
    9300 => -26,
    9301 => -26,
    9302 => -26,
    9303 => -26,
    9304 => -26,
    9305 => -26,
    9306 => -26,
    9307 => -26,
    9308 => -26,
    9309 => -26,
    9310 => -26,
    9311 => -26,
    9312 => -26,
    9313 => -26,
    9314 => -26,
    9315 => -26,
    9316 => -26,
    9317 => -26,
    9318 => -26,
    9319 => -26,
    9320 => -26,
    9321 => -26,
    9322 => -26,
    9323 => -26,
    9324 => -26,
    9325 => -27,
    9326 => -27,
    9327 => -27,
    9328 => -27,
    9329 => -27,
    9330 => -27,
    9331 => -27,
    9332 => -27,
    9333 => -27,
    9334 => -27,
    9335 => -27,
    9336 => -27,
    9337 => -27,
    9338 => -27,
    9339 => -27,
    9340 => -27,
    9341 => -27,
    9342 => -27,
    9343 => -27,
    9344 => -27,
    9345 => -27,
    9346 => -27,
    9347 => -27,
    9348 => -27,
    9349 => -27,
    9350 => -27,
    9351 => -27,
    9352 => -27,
    9353 => -27,
    9354 => -27,
    9355 => -27,
    9356 => -27,
    9357 => -27,
    9358 => -27,
    9359 => -27,
    9360 => -27,
    9361 => -27,
    9362 => -27,
    9363 => -27,
    9364 => -27,
    9365 => -27,
    9366 => -27,
    9367 => -27,
    9368 => -27,
    9369 => -27,
    9370 => -28,
    9371 => -28,
    9372 => -28,
    9373 => -28,
    9374 => -28,
    9375 => -28,
    9376 => -28,
    9377 => -28,
    9378 => -28,
    9379 => -28,
    9380 => -28,
    9381 => -28,
    9382 => -28,
    9383 => -28,
    9384 => -28,
    9385 => -28,
    9386 => -28,
    9387 => -28,
    9388 => -28,
    9389 => -28,
    9390 => -28,
    9391 => -28,
    9392 => -28,
    9393 => -28,
    9394 => -28,
    9395 => -28,
    9396 => -28,
    9397 => -28,
    9398 => -28,
    9399 => -28,
    9400 => -28,
    9401 => -28,
    9402 => -28,
    9403 => -28,
    9404 => -28,
    9405 => -28,
    9406 => -28,
    9407 => -28,
    9408 => -28,
    9409 => -28,
    9410 => -28,
    9411 => -28,
    9412 => -28,
    9413 => -28,
    9414 => -28,
    9415 => -28,
    9416 => -28,
    9417 => -29,
    9418 => -29,
    9419 => -29,
    9420 => -29,
    9421 => -29,
    9422 => -29,
    9423 => -29,
    9424 => -29,
    9425 => -29,
    9426 => -29,
    9427 => -29,
    9428 => -29,
    9429 => -29,
    9430 => -29,
    9431 => -29,
    9432 => -29,
    9433 => -29,
    9434 => -29,
    9435 => -29,
    9436 => -29,
    9437 => -29,
    9438 => -29,
    9439 => -29,
    9440 => -29,
    9441 => -29,
    9442 => -29,
    9443 => -29,
    9444 => -29,
    9445 => -29,
    9446 => -29,
    9447 => -29,
    9448 => -29,
    9449 => -29,
    9450 => -29,
    9451 => -29,
    9452 => -29,
    9453 => -29,
    9454 => -29,
    9455 => -29,
    9456 => -29,
    9457 => -29,
    9458 => -29,
    9459 => -29,
    9460 => -29,
    9461 => -29,
    9462 => -29,
    9463 => -30,
    9464 => -30,
    9465 => -30,
    9466 => -30,
    9467 => -30,
    9468 => -30,
    9469 => -30,
    9470 => -30,
    9471 => -30,
    9472 => -30,
    9473 => -30,
    9474 => -30,
    9475 => -30,
    9476 => -30,
    9477 => -30,
    9478 => -30,
    9479 => -30,
    9480 => -30,
    9481 => -30,
    9482 => -30,
    9483 => -30,
    9484 => -30,
    9485 => -30,
    9486 => -30,
    9487 => -30,
    9488 => -30,
    9489 => -30,
    9490 => -30,
    9491 => -30,
    9492 => -30,
    9493 => -30,
    9494 => -30,
    9495 => -30,
    9496 => -30,
    9497 => -30,
    9498 => -30,
    9499 => -30,
    9500 => -30,
    9501 => -30,
    9502 => -30,
    9503 => -30,
    9504 => -30,
    9505 => -30,
    9506 => -30,
    9507 => -30,
    9508 => -30,
    9509 => -30,
    9510 => -31,
    9511 => -31,
    9512 => -31,
    9513 => -31,
    9514 => -31,
    9515 => -31,
    9516 => -31,
    9517 => -31,
    9518 => -31,
    9519 => -31,
    9520 => -31,
    9521 => -31,
    9522 => -31,
    9523 => -31,
    9524 => -31,
    9525 => -31,
    9526 => -31,
    9527 => -31,
    9528 => -31,
    9529 => -31,
    9530 => -31,
    9531 => -31,
    9532 => -31,
    9533 => -31,
    9534 => -31,
    9535 => -31,
    9536 => -31,
    9537 => -31,
    9538 => -31,
    9539 => -31,
    9540 => -31,
    9541 => -31,
    9542 => -31,
    9543 => -31,
    9544 => -31,
    9545 => -31,
    9546 => -31,
    9547 => -31,
    9548 => -31,
    9549 => -31,
    9550 => -31,
    9551 => -31,
    9552 => -31,
    9553 => -31,
    9554 => -31,
    9555 => -31,
    9556 => -31,
    9557 => -31,
    9558 => -32,
    9559 => -32,
    9560 => -32,
    9561 => -32,
    9562 => -32,
    9563 => -32,
    9564 => -32,
    9565 => -32,
    9566 => -32,
    9567 => -32,
    9568 => -32,
    9569 => -32,
    9570 => -32,
    9571 => -32,
    9572 => -32,
    9573 => -32,
    9574 => -32,
    9575 => -32,
    9576 => -32,
    9577 => -32,
    9578 => -32,
    9579 => -32,
    9580 => -32,
    9581 => -32,
    9582 => -32,
    9583 => -32,
    9584 => -32,
    9585 => -32,
    9586 => -32,
    9587 => -32,
    9588 => -32,
    9589 => -32,
    9590 => -32,
    9591 => -32,
    9592 => -32,
    9593 => -32,
    9594 => -32,
    9595 => -32,
    9596 => -32,
    9597 => -32,
    9598 => -32,
    9599 => -32,
    9600 => -32,
    9601 => -32,
    9602 => -32,
    9603 => -32,
    9604 => -32,
    9605 => -32,
    9606 => -33,
    9607 => -33,
    9608 => -33,
    9609 => -33,
    9610 => -33,
    9611 => -33,
    9612 => -33,
    9613 => -33,
    9614 => -33,
    9615 => -33,
    9616 => -33,
    9617 => -33,
    9618 => -33,
    9619 => -33,
    9620 => -33,
    9621 => -33,
    9622 => -33,
    9623 => -33,
    9624 => -33,
    9625 => -33,
    9626 => -33,
    9627 => -33,
    9628 => -33,
    9629 => -33,
    9630 => -33,
    9631 => -33,
    9632 => -33,
    9633 => -33,
    9634 => -33,
    9635 => -33,
    9636 => -33,
    9637 => -33,
    9638 => -33,
    9639 => -33,
    9640 => -33,
    9641 => -33,
    9642 => -33,
    9643 => -33,
    9644 => -33,
    9645 => -33,
    9646 => -33,
    9647 => -33,
    9648 => -33,
    9649 => -33,
    9650 => -33,
    9651 => -33,
    9652 => -33,
    9653 => -33,
    9654 => -34,
    9655 => -34,
    9656 => -34,
    9657 => -34,
    9658 => -34,
    9659 => -34,
    9660 => -34,
    9661 => -34,
    9662 => -34,
    9663 => -34,
    9664 => -34,
    9665 => -34,
    9666 => -34,
    9667 => -34,
    9668 => -34,
    9669 => -34,
    9670 => -34,
    9671 => -34,
    9672 => -34,
    9673 => -34,
    9674 => -34,
    9675 => -34,
    9676 => -34,
    9677 => -34,
    9678 => -34,
    9679 => -34,
    9680 => -34,
    9681 => -34,
    9682 => -34,
    9683 => -34,
    9684 => -34,
    9685 => -34,
    9686 => -34,
    9687 => -34,
    9688 => -34,
    9689 => -34,
    9690 => -34,
    9691 => -34,
    9692 => -34,
    9693 => -34,
    9694 => -34,
    9695 => -34,
    9696 => -34,
    9697 => -34,
    9698 => -34,
    9699 => -34,
    9700 => -34,
    9701 => -34,
    9702 => -34,
    9703 => -34,
    9704 => -35,
    9705 => -35,
    9706 => -35,
    9707 => -35,
    9708 => -35,
    9709 => -35,
    9710 => -35,
    9711 => -35,
    9712 => -35,
    9713 => -35,
    9714 => -35,
    9715 => -35,
    9716 => -35,
    9717 => -35,
    9718 => -35,
    9719 => -35,
    9720 => -35,
    9721 => -35,
    9722 => -35,
    9723 => -35,
    9724 => -35,
    9725 => -35,
    9726 => -35,
    9727 => -35,
    9728 => -35,
    9729 => -35,
    9730 => -35,
    9731 => -35,
    9732 => -35,
    9733 => -35,
    9734 => -35,
    9735 => -35,
    9736 => -35,
    9737 => -35,
    9738 => -35,
    9739 => -35,
    9740 => -35,
    9741 => -35,
    9742 => -35,
    9743 => -35,
    9744 => -35,
    9745 => -35,
    9746 => -35,
    9747 => -35,
    9748 => -35,
    9749 => -35,
    9750 => -35,
    9751 => -35,
    9752 => -35,
    9753 => -36,
    9754 => -36,
    9755 => -36,
    9756 => -36,
    9757 => -36,
    9758 => -36,
    9759 => -36,
    9760 => -36,
    9761 => -36,
    9762 => -36,
    9763 => -36,
    9764 => -36,
    9765 => -36,
    9766 => -36,
    9767 => -36,
    9768 => -36,
    9769 => -36,
    9770 => -36,
    9771 => -36,
    9772 => -36,
    9773 => -36,
    9774 => -36,
    9775 => -36,
    9776 => -36,
    9777 => -36,
    9778 => -36,
    9779 => -36,
    9780 => -36,
    9781 => -36,
    9782 => -36,
    9783 => -36,
    9784 => -36,
    9785 => -36,
    9786 => -36,
    9787 => -36,
    9788 => -36,
    9789 => -36,
    9790 => -36,
    9791 => -36,
    9792 => -36,
    9793 => -36,
    9794 => -36,
    9795 => -36,
    9796 => -36,
    9797 => -36,
    9798 => -36,
    9799 => -36,
    9800 => -36,
    9801 => -36,
    9802 => -36,
    9803 => -36,
    9804 => -37,
    9805 => -37,
    9806 => -37,
    9807 => -37,
    9808 => -37,
    9809 => -37,
    9810 => -37,
    9811 => -37,
    9812 => -37,
    9813 => -37,
    9814 => -37,
    9815 => -37,
    9816 => -37,
    9817 => -37,
    9818 => -37,
    9819 => -37,
    9820 => -37,
    9821 => -37,
    9822 => -37,
    9823 => -37,
    9824 => -37,
    9825 => -37,
    9826 => -37,
    9827 => -37,
    9828 => -37,
    9829 => -37,
    9830 => -37,
    9831 => -37,
    9832 => -37,
    9833 => -37,
    9834 => -37,
    9835 => -37,
    9836 => -37,
    9837 => -37,
    9838 => -37,
    9839 => -37,
    9840 => -37,
    9841 => -37,
    9842 => -37,
    9843 => -37,
    9844 => -37,
    9845 => -37,
    9846 => -37,
    9847 => -37,
    9848 => -37,
    9849 => -37,
    9850 => -37,
    9851 => -37,
    9852 => -37,
    9853 => -37,
    9854 => -37,
    9855 => -38,
    9856 => -38,
    9857 => -38,
    9858 => -38,
    9859 => -38,
    9860 => -38,
    9861 => -38,
    9862 => -38,
    9863 => -38,
    9864 => -38,
    9865 => -38,
    9866 => -38,
    9867 => -38,
    9868 => -38,
    9869 => -38,
    9870 => -38,
    9871 => -38,
    9872 => -38,
    9873 => -38,
    9874 => -38,
    9875 => -38,
    9876 => -38,
    9877 => -38,
    9878 => -38,
    9879 => -38,
    9880 => -38,
    9881 => -38,
    9882 => -38,
    9883 => -38,
    9884 => -38,
    9885 => -38,
    9886 => -38,
    9887 => -38,
    9888 => -38,
    9889 => -38,
    9890 => -38,
    9891 => -38,
    9892 => -38,
    9893 => -38,
    9894 => -38,
    9895 => -38,
    9896 => -38,
    9897 => -38,
    9898 => -38,
    9899 => -38,
    9900 => -38,
    9901 => -38,
    9902 => -38,
    9903 => -38,
    9904 => -38,
    9905 => -38,
    9906 => -38,
    9907 => -39,
    9908 => -39,
    9909 => -39,
    9910 => -39,
    9911 => -39,
    9912 => -39,
    9913 => -39,
    9914 => -39,
    9915 => -39,
    9916 => -39,
    9917 => -39,
    9918 => -39,
    9919 => -39,
    9920 => -39,
    9921 => -39,
    9922 => -39,
    9923 => -39,
    9924 => -39,
    9925 => -39,
    9926 => -39,
    9927 => -39,
    9928 => -39,
    9929 => -39,
    9930 => -39,
    9931 => -39,
    9932 => -39,
    9933 => -39,
    9934 => -39,
    9935 => -39,
    9936 => -39,
    9937 => -39,
    9938 => -39,
    9939 => -39,
    9940 => -39,
    9941 => -39,
    9942 => -39,
    9943 => -39,
    9944 => -39,
    9945 => -39,
    9946 => -39,
    9947 => -39,
    9948 => -39,
    9949 => -39,
    9950 => -39,
    9951 => -39,
    9952 => -39,
    9953 => -39,
    9954 => -39,
    9955 => -39,
    9956 => -39,
    9957 => -39,
    9958 => -39,
    9959 => -39,
    9960 => -40,
    9961 => -40,
    9962 => -40,
    9963 => -40,
    9964 => -40,
    9965 => -40,
    9966 => -40,
    9967 => -40,
    9968 => -40,
    9969 => -40,
    9970 => -40,
    9971 => -40,
    9972 => -40,
    9973 => -40,
    9974 => -40,
    9975 => -40,
    9976 => -40,
    9977 => -40,
    9978 => -40,
    9979 => -40,
    9980 => -40,
    9981 => -40,
    9982 => -40,
    9983 => -40,
    9984 => -40,
    9985 => -40,
    9986 => -40,
    9987 => -40,
    9988 => -40,
    9989 => -40,
    9990 => -40,
    9991 => -40,
    9992 => -40,
    9993 => -40,
    9994 => -40,
    9995 => -40,
    9996 => -40,
    9997 => -40,
    9998 => -40,
    9999 => -40,
    10000 => -40,
    10001 => -40,
    10002 => -40,
    10003 => -40,
    10004 => -40,
    10005 => -40,
    10006 => -40,
    10007 => -40,
    10008 => -40,
    10009 => -40,
    10010 => -40,
    10011 => -40,
    10012 => -40,
    10013 => -41,
    10014 => -41,
    10015 => -41,
    10016 => -41,
    10017 => -41,
    10018 => -41,
    10019 => -41,
    10020 => -41,
    10021 => -41,
    10022 => -41,
    10023 => -41,
    10024 => -41,
    10025 => -41,
    10026 => -41,
    10027 => -41,
    10028 => -41,
    10029 => -41,
    10030 => -41,
    10031 => -41,
    10032 => -41,
    10033 => -41,
    10034 => -41,
    10035 => -41,
    10036 => -41,
    10037 => -41,
    10038 => -41,
    10039 => -41,
    10040 => -41,
    10041 => -41,
    10042 => -41,
    10043 => -41,
    10044 => -41,
    10045 => -41,
    10046 => -41,
    10047 => -41,
    10048 => -41,
    10049 => -41,
    10050 => -41,
    10051 => -41,
    10052 => -41,
    10053 => -41,
    10054 => -41,
    10055 => -41,
    10056 => -41,
    10057 => -41,
    10058 => -41,
    10059 => -41,
    10060 => -41,
    10061 => -41,
    10062 => -41,
    10063 => -41,
    10064 => -41,
    10065 => -41,
    10066 => -41,
    10067 => -41,
    10068 => -42,
    10069 => -42,
    10070 => -42,
    10071 => -42,
    10072 => -42,
    10073 => -42,
    10074 => -42,
    10075 => -42,
    10076 => -42,
    10077 => -42,
    10078 => -42,
    10079 => -42,
    10080 => -42,
    10081 => -42,
    10082 => -42,
    10083 => -42,
    10084 => -42,
    10085 => -42,
    10086 => -42,
    10087 => -42,
    10088 => -42,
    10089 => -42,
    10090 => -42,
    10091 => -42,
    10092 => -42,
    10093 => -42,
    10094 => -42,
    10095 => -42,
    10096 => -42,
    10097 => -42,
    10098 => -42,
    10099 => -42,
    10100 => -42,
    10101 => -42,
    10102 => -42,
    10103 => -42,
    10104 => -42,
    10105 => -42,
    10106 => -42,
    10107 => -42,
    10108 => -42,
    10109 => -42,
    10110 => -42,
    10111 => -42,
    10112 => -42,
    10113 => -42,
    10114 => -42,
    10115 => -42,
    10116 => -42,
    10117 => -42,
    10118 => -42,
    10119 => -42,
    10120 => -42,
    10121 => -42,
    10122 => -42,
    10123 => -43,
    10124 => -43,
    10125 => -43,
    10126 => -43,
    10127 => -43,
    10128 => -43,
    10129 => -43,
    10130 => -43,
    10131 => -43,
    10132 => -43,
    10133 => -43,
    10134 => -43,
    10135 => -43,
    10136 => -43,
    10137 => -43,
    10138 => -43,
    10139 => -43,
    10140 => -43,
    10141 => -43,
    10142 => -43,
    10143 => -43,
    10144 => -43,
    10145 => -43,
    10146 => -43,
    10147 => -43,
    10148 => -43,
    10149 => -43,
    10150 => -43,
    10151 => -43,
    10152 => -43,
    10153 => -43,
    10154 => -43,
    10155 => -43,
    10156 => -43,
    10157 => -43,
    10158 => -43,
    10159 => -43,
    10160 => -43,
    10161 => -43,
    10162 => -43,
    10163 => -43,
    10164 => -43,
    10165 => -43,
    10166 => -43,
    10167 => -43,
    10168 => -43,
    10169 => -43,
    10170 => -43,
    10171 => -43,
    10172 => -43,
    10173 => -43,
    10174 => -43,
    10175 => -43,
    10176 => -43,
    10177 => -43,
    10178 => -43,
    10179 => -43,
    10180 => -44,
    10181 => -44,
    10182 => -44,
    10183 => -44,
    10184 => -44,
    10185 => -44,
    10186 => -44,
    10187 => -44,
    10188 => -44,
    10189 => -44,
    10190 => -44,
    10191 => -44,
    10192 => -44,
    10193 => -44,
    10194 => -44,
    10195 => -44,
    10196 => -44,
    10197 => -44,
    10198 => -44,
    10199 => -44,
    10200 => -44,
    10201 => -44,
    10202 => -44,
    10203 => -44,
    10204 => -44,
    10205 => -44,
    10206 => -44,
    10207 => -44,
    10208 => -44,
    10209 => -44,
    10210 => -44,
    10211 => -44,
    10212 => -44,
    10213 => -44,
    10214 => -44,
    10215 => -44,
    10216 => -44,
    10217 => -44,
    10218 => -44,
    10219 => -44,
    10220 => -44,
    10221 => -44,
    10222 => -44,
    10223 => -44,
    10224 => -44,
    10225 => -44,
    10226 => -44,
    10227 => -44,
    10228 => -44,
    10229 => -44,
    10230 => -44,
    10231 => -44,
    10232 => -44,
    10233 => -44,
    10234 => -44,
    10235 => -44,
    10236 => -44,
    10237 => -44,
    10238 => -45,
    10239 => -45,
    10240 => -45,
    10241 => -45,
    10242 => -45,
    10243 => -45,
    10244 => -45,
    10245 => -45,
    10246 => -45,
    10247 => -45,
    10248 => -45,
    10249 => -45,
    10250 => -45,
    10251 => -45,
    10252 => -45,
    10253 => -45,
    10254 => -45,
    10255 => -45,
    10256 => -45,
    10257 => -45,
    10258 => -45,
    10259 => -45,
    10260 => -45,
    10261 => -45,
    10262 => -45,
    10263 => -45,
    10264 => -45,
    10265 => -45,
    10266 => -45,
    10267 => -45,
    10268 => -45,
    10269 => -45,
    10270 => -45,
    10271 => -45,
    10272 => -45,
    10273 => -45,
    10274 => -45,
    10275 => -45,
    10276 => -45,
    10277 => -45,
    10278 => -45,
    10279 => -45,
    10280 => -45,
    10281 => -45,
    10282 => -45,
    10283 => -45,
    10284 => -45,
    10285 => -45,
    10286 => -45,
    10287 => -45,
    10288 => -45,
    10289 => -45,
    10290 => -45,
    10291 => -45,
    10292 => -45,
    10293 => -45,
    10294 => -45,
    10295 => -45,
    10296 => -45,
    10297 => -46,
    10298 => -46,
    10299 => -46,
    10300 => -46,
    10301 => -46,
    10302 => -46,
    10303 => -46,
    10304 => -46,
    10305 => -46,
    10306 => -46,
    10307 => -46,
    10308 => -46,
    10309 => -46,
    10310 => -46,
    10311 => -46,
    10312 => -46,
    10313 => -46,
    10314 => -46,
    10315 => -46,
    10316 => -46,
    10317 => -46,
    10318 => -46,
    10319 => -46,
    10320 => -46,
    10321 => -46,
    10322 => -46,
    10323 => -46,
    10324 => -46,
    10325 => -46,
    10326 => -46,
    10327 => -46,
    10328 => -46,
    10329 => -46,
    10330 => -46,
    10331 => -46,
    10332 => -46,
    10333 => -46,
    10334 => -46,
    10335 => -46,
    10336 => -46,
    10337 => -46,
    10338 => -46,
    10339 => -46,
    10340 => -46,
    10341 => -46,
    10342 => -46,
    10343 => -46,
    10344 => -46,
    10345 => -46,
    10346 => -46,
    10347 => -46,
    10348 => -46,
    10349 => -46,
    10350 => -46,
    10351 => -46,
    10352 => -46,
    10353 => -46,
    10354 => -46,
    10355 => -46,
    10356 => -46,
    10357 => -47,
    10358 => -47,
    10359 => -47,
    10360 => -47,
    10361 => -47,
    10362 => -47,
    10363 => -47,
    10364 => -47,
    10365 => -47,
    10366 => -47,
    10367 => -47,
    10368 => -47,
    10369 => -47,
    10370 => -47,
    10371 => -47,
    10372 => -47,
    10373 => -47,
    10374 => -47,
    10375 => -47,
    10376 => -47,
    10377 => -47,
    10378 => -47,
    10379 => -47,
    10380 => -47,
    10381 => -47,
    10382 => -47,
    10383 => -47,
    10384 => -47,
    10385 => -47,
    10386 => -47,
    10387 => -47,
    10388 => -47,
    10389 => -47,
    10390 => -47,
    10391 => -47,
    10392 => -47,
    10393 => -47,
    10394 => -47,
    10395 => -47,
    10396 => -47,
    10397 => -47,
    10398 => -47,
    10399 => -47,
    10400 => -47,
    10401 => -47,
    10402 => -47,
    10403 => -47,
    10404 => -47,
    10405 => -47,
    10406 => -47,
    10407 => -47,
    10408 => -47,
    10409 => -47,
    10410 => -47,
    10411 => -47,
    10412 => -47,
    10413 => -47,
    10414 => -47,
    10415 => -47,
    10416 => -47,
    10417 => -47,
    10418 => -47,
    10419 => -47,
    10420 => -48,
    10421 => -48,
    10422 => -48,
    10423 => -48,
    10424 => -48,
    10425 => -48,
    10426 => -48,
    10427 => -48,
    10428 => -48,
    10429 => -48,
    10430 => -48,
    10431 => -48,
    10432 => -48,
    10433 => -48,
    10434 => -48,
    10435 => -48,
    10436 => -48,
    10437 => -48,
    10438 => -48,
    10439 => -48,
    10440 => -48,
    10441 => -48,
    10442 => -48,
    10443 => -48,
    10444 => -48,
    10445 => -48,
    10446 => -48,
    10447 => -48,
    10448 => -48,
    10449 => -48,
    10450 => -48,
    10451 => -48,
    10452 => -48,
    10453 => -48,
    10454 => -48,
    10455 => -48,
    10456 => -48,
    10457 => -48,
    10458 => -48,
    10459 => -48,
    10460 => -48,
    10461 => -48,
    10462 => -48,
    10463 => -48,
    10464 => -48,
    10465 => -48,
    10466 => -48,
    10467 => -48,
    10468 => -48,
    10469 => -48,
    10470 => -48,
    10471 => -48,
    10472 => -48,
    10473 => -48,
    10474 => -48,
    10475 => -48,
    10476 => -48,
    10477 => -48,
    10478 => -48,
    10479 => -48,
    10480 => -48,
    10481 => -48,
    10482 => -48,
    10483 => -48,
    10484 => -49,
    10485 => -49,
    10486 => -49,
    10487 => -49,
    10488 => -49,
    10489 => -49,
    10490 => -49,
    10491 => -49,
    10492 => -49,
    10493 => -49,
    10494 => -49,
    10495 => -49,
    10496 => -49,
    10497 => -49,
    10498 => -49,
    10499 => -49,
    10500 => -49,
    10501 => -49,
    10502 => -49,
    10503 => -49,
    10504 => -49,
    10505 => -49,
    10506 => -49,
    10507 => -49,
    10508 => -49,
    10509 => -49,
    10510 => -49,
    10511 => -49,
    10512 => -49,
    10513 => -49,
    10514 => -49,
    10515 => -49,
    10516 => -49,
    10517 => -49,
    10518 => -49,
    10519 => -49,
    10520 => -49,
    10521 => -49,
    10522 => -49,
    10523 => -49,
    10524 => -49,
    10525 => -49,
    10526 => -49,
    10527 => -49,
    10528 => -49,
    10529 => -49,
    10530 => -49,
    10531 => -49,
    10532 => -49,
    10533 => -49,
    10534 => -49,
    10535 => -49,
    10536 => -49,
    10537 => -49,
    10538 => -49,
    10539 => -49,
    10540 => -49,
    10541 => -49,
    10542 => -49,
    10543 => -49,
    10544 => -49,
    10545 => -49,
    10546 => -49,
    10547 => -49,
    10548 => -49,
    10549 => -50,
    10550 => -50,
    10551 => -50,
    10552 => -50,
    10553 => -50,
    10554 => -50,
    10555 => -50,
    10556 => -50,
    10557 => -50,
    10558 => -50,
    10559 => -50,
    10560 => -50,
    10561 => -50,
    10562 => -50,
    10563 => -50,
    10564 => -50,
    10565 => -50,
    10566 => -50,
    10567 => -50,
    10568 => -50,
    10569 => -50,
    10570 => -50,
    10571 => -50,
    10572 => -50,
    10573 => -50,
    10574 => -50,
    10575 => -50,
    10576 => -50,
    10577 => -50,
    10578 => -50,
    10579 => -50,
    10580 => -50,
    10581 => -50,
    10582 => -50,
    10583 => -50,
    10584 => -50,
    10585 => -50,
    10586 => -50,
    10587 => -50,
    10588 => -50,
    10589 => -50,
    10590 => -50,
    10591 => -50,
    10592 => -50,
    10593 => -50,
    10594 => -50,
    10595 => -50,
    10596 => -50,
    10597 => -50,
    10598 => -50,
    10599 => -50,
    10600 => -50,
    10601 => -50,
    10602 => -50,
    10603 => -50,
    10604 => -50,
    10605 => -50,
    10606 => -50,
    10607 => -50,
    10608 => -50,
    10609 => -50,
    10610 => -50,
    10611 => -50,
    10612 => -50,
    10613 => -50,
    10614 => -50,
    10615 => -50,
    10616 => -50,
    10617 => -51,
    10618 => -51,
    10619 => -51,
    10620 => -51,
    10621 => -51,
    10622 => -51,
    10623 => -51,
    10624 => -51,
    10625 => -51,
    10626 => -51,
    10627 => -51,
    10628 => -51,
    10629 => -51,
    10630 => -51,
    10631 => -51,
    10632 => -51,
    10633 => -51,
    10634 => -51,
    10635 => -51,
    10636 => -51,
    10637 => -51,
    10638 => -51,
    10639 => -51,
    10640 => -51,
    10641 => -51,
    10642 => -51,
    10643 => -51,
    10644 => -51,
    10645 => -51,
    10646 => -51,
    10647 => -51,
    10648 => -51,
    10649 => -51,
    10650 => -51,
    10651 => -51,
    10652 => -51,
    10653 => -51,
    10654 => -51,
    10655 => -51,
    10656 => -51,
    10657 => -51,
    10658 => -51,
    10659 => -51,
    10660 => -51,
    10661 => -51,
    10662 => -51,
    10663 => -51,
    10664 => -51,
    10665 => -51,
    10666 => -51,
    10667 => -51,
    10668 => -51,
    10669 => -51,
    10670 => -51,
    10671 => -51,
    10672 => -51,
    10673 => -51,
    10674 => -51,
    10675 => -51,
    10676 => -51,
    10677 => -51,
    10678 => -51,
    10679 => -51,
    10680 => -51,
    10681 => -51,
    10682 => -51,
    10683 => -51,
    10684 => -51,
    10685 => -51,
    10686 => -51,
    10687 => -51,
    10688 => -52,
    10689 => -52,
    10690 => -52,
    10691 => -52,
    10692 => -52,
    10693 => -52,
    10694 => -52,
    10695 => -52,
    10696 => -52,
    10697 => -52,
    10698 => -52,
    10699 => -52,
    10700 => -52,
    10701 => -52,
    10702 => -52,
    10703 => -52,
    10704 => -52,
    10705 => -52,
    10706 => -52,
    10707 => -52,
    10708 => -52,
    10709 => -52,
    10710 => -52,
    10711 => -52,
    10712 => -52,
    10713 => -52,
    10714 => -52,
    10715 => -52,
    10716 => -52,
    10717 => -52,
    10718 => -52,
    10719 => -52,
    10720 => -52,
    10721 => -52,
    10722 => -52,
    10723 => -52,
    10724 => -52,
    10725 => -52,
    10726 => -52,
    10727 => -52,
    10728 => -52,
    10729 => -52,
    10730 => -52,
    10731 => -52,
    10732 => -52,
    10733 => -52,
    10734 => -52,
    10735 => -52,
    10736 => -52,
    10737 => -52,
    10738 => -52,
    10739 => -52,
    10740 => -52,
    10741 => -52,
    10742 => -52,
    10743 => -52,
    10744 => -52,
    10745 => -52,
    10746 => -52,
    10747 => -52,
    10748 => -52,
    10749 => -52,
    10750 => -52,
    10751 => -52,
    10752 => -52,
    10753 => -52,
    10754 => -52,
    10755 => -52,
    10756 => -52,
    10757 => -52,
    10758 => -52,
    10759 => -52,
    10760 => -52,
    10761 => -53,
    10762 => -53,
    10763 => -53,
    10764 => -53,
    10765 => -53,
    10766 => -53,
    10767 => -53,
    10768 => -53,
    10769 => -53,
    10770 => -53,
    10771 => -53,
    10772 => -53,
    10773 => -53,
    10774 => -53,
    10775 => -53,
    10776 => -53,
    10777 => -53,
    10778 => -53,
    10779 => -53,
    10780 => -53,
    10781 => -53,
    10782 => -53,
    10783 => -53,
    10784 => -53,
    10785 => -53,
    10786 => -53,
    10787 => -53,
    10788 => -53,
    10789 => -53,
    10790 => -53,
    10791 => -53,
    10792 => -53,
    10793 => -53,
    10794 => -53,
    10795 => -53,
    10796 => -53,
    10797 => -53,
    10798 => -53,
    10799 => -53,
    10800 => -53,
    10801 => -53,
    10802 => -53,
    10803 => -53,
    10804 => -53,
    10805 => -53,
    10806 => -53,
    10807 => -53,
    10808 => -53,
    10809 => -53,
    10810 => -53,
    10811 => -53,
    10812 => -53,
    10813 => -53,
    10814 => -53,
    10815 => -53,
    10816 => -53,
    10817 => -53,
    10818 => -53,
    10819 => -53,
    10820 => -53,
    10821 => -53,
    10822 => -53,
    10823 => -53,
    10824 => -53,
    10825 => -53,
    10826 => -53,
    10827 => -53,
    10828 => -53,
    10829 => -53,
    10830 => -53,
    10831 => -53,
    10832 => -53,
    10833 => -53,
    10834 => -53,
    10835 => -53,
    10836 => -53,
    10837 => -53,
    10838 => -54,
    10839 => -54,
    10840 => -54,
    10841 => -54,
    10842 => -54,
    10843 => -54,
    10844 => -54,
    10845 => -54,
    10846 => -54,
    10847 => -54,
    10848 => -54,
    10849 => -54,
    10850 => -54,
    10851 => -54,
    10852 => -54,
    10853 => -54,
    10854 => -54,
    10855 => -54,
    10856 => -54,
    10857 => -54,
    10858 => -54,
    10859 => -54,
    10860 => -54,
    10861 => -54,
    10862 => -54,
    10863 => -54,
    10864 => -54,
    10865 => -54,
    10866 => -54,
    10867 => -54,
    10868 => -54,
    10869 => -54,
    10870 => -54,
    10871 => -54,
    10872 => -54,
    10873 => -54,
    10874 => -54,
    10875 => -54,
    10876 => -54,
    10877 => -54,
    10878 => -54,
    10879 => -54,
    10880 => -54,
    10881 => -54,
    10882 => -54,
    10883 => -54,
    10884 => -54,
    10885 => -54,
    10886 => -54,
    10887 => -54,
    10888 => -54,
    10889 => -54,
    10890 => -54,
    10891 => -54,
    10892 => -54,
    10893 => -54,
    10894 => -54,
    10895 => -54,
    10896 => -54,
    10897 => -54,
    10898 => -54,
    10899 => -54,
    10900 => -54,
    10901 => -54,
    10902 => -54,
    10903 => -54,
    10904 => -54,
    10905 => -54,
    10906 => -54,
    10907 => -54,
    10908 => -54,
    10909 => -54,
    10910 => -54,
    10911 => -54,
    10912 => -54,
    10913 => -54,
    10914 => -54,
    10915 => -54,
    10916 => -54,
    10917 => -54,
    10918 => -55,
    10919 => -55,
    10920 => -55,
    10921 => -55,
    10922 => -55,
    10923 => -55,
    10924 => -55,
    10925 => -55,
    10926 => -55,
    10927 => -55,
    10928 => -55,
    10929 => -55,
    10930 => -55,
    10931 => -55,
    10932 => -55,
    10933 => -55,
    10934 => -55,
    10935 => -55,
    10936 => -55,
    10937 => -55,
    10938 => -55,
    10939 => -55,
    10940 => -55,
    10941 => -55,
    10942 => -55,
    10943 => -55,
    10944 => -55,
    10945 => -55,
    10946 => -55,
    10947 => -55,
    10948 => -55,
    10949 => -55,
    10950 => -55,
    10951 => -55,
    10952 => -55,
    10953 => -55,
    10954 => -55,
    10955 => -55,
    10956 => -55,
    10957 => -55,
    10958 => -55,
    10959 => -55,
    10960 => -55,
    10961 => -55,
    10962 => -55,
    10963 => -55,
    10964 => -55,
    10965 => -55,
    10966 => -55,
    10967 => -55,
    10968 => -55,
    10969 => -55,
    10970 => -55,
    10971 => -55,
    10972 => -55,
    10973 => -55,
    10974 => -55,
    10975 => -55,
    10976 => -55,
    10977 => -55,
    10978 => -55,
    10979 => -55,
    10980 => -55,
    10981 => -55,
    10982 => -55,
    10983 => -55,
    10984 => -55,
    10985 => -55,
    10986 => -55,
    10987 => -55,
    10988 => -55,
    10989 => -55,
    10990 => -55,
    10991 => -55,
    10992 => -55,
    10993 => -55,
    10994 => -55,
    10995 => -55,
    10996 => -55,
    10997 => -55,
    10998 => -55,
    10999 => -55,
    11000 => -55,
    11001 => -55,
    11002 => -55,
    11003 => -56,
    11004 => -56,
    11005 => -56,
    11006 => -56,
    11007 => -56,
    11008 => -56,
    11009 => -56,
    11010 => -56,
    11011 => -56,
    11012 => -56,
    11013 => -56,
    11014 => -56,
    11015 => -56,
    11016 => -56,
    11017 => -56,
    11018 => -56,
    11019 => -56,
    11020 => -56,
    11021 => -56,
    11022 => -56,
    11023 => -56,
    11024 => -56,
    11025 => -56,
    11026 => -56,
    11027 => -56,
    11028 => -56,
    11029 => -56,
    11030 => -56,
    11031 => -56,
    11032 => -56,
    11033 => -56,
    11034 => -56,
    11035 => -56,
    11036 => -56,
    11037 => -56,
    11038 => -56,
    11039 => -56,
    11040 => -56,
    11041 => -56,
    11042 => -56,
    11043 => -56,
    11044 => -56,
    11045 => -56,
    11046 => -56,
    11047 => -56,
    11048 => -56,
    11049 => -56,
    11050 => -56,
    11051 => -56,
    11052 => -56,
    11053 => -56,
    11054 => -56,
    11055 => -56,
    11056 => -56,
    11057 => -56,
    11058 => -56,
    11059 => -56,
    11060 => -56,
    11061 => -56,
    11062 => -56,
    11063 => -56,
    11064 => -56,
    11065 => -56,
    11066 => -56,
    11067 => -56,
    11068 => -56,
    11069 => -56,
    11070 => -56,
    11071 => -56,
    11072 => -56,
    11073 => -56,
    11074 => -56,
    11075 => -56,
    11076 => -56,
    11077 => -56,
    11078 => -56,
    11079 => -56,
    11080 => -56,
    11081 => -56,
    11082 => -56,
    11083 => -56,
    11084 => -56,
    11085 => -56,
    11086 => -56,
    11087 => -56,
    11088 => -56,
    11089 => -56,
    11090 => -56,
    11091 => -56,
    11092 => -56,
    11093 => -56,
    11094 => -57,
    11095 => -57,
    11096 => -57,
    11097 => -57,
    11098 => -57,
    11099 => -57,
    11100 => -57,
    11101 => -57,
    11102 => -57,
    11103 => -57,
    11104 => -57,
    11105 => -57,
    11106 => -57,
    11107 => -57,
    11108 => -57,
    11109 => -57,
    11110 => -57,
    11111 => -57,
    11112 => -57,
    11113 => -57,
    11114 => -57,
    11115 => -57,
    11116 => -57,
    11117 => -57,
    11118 => -57,
    11119 => -57,
    11120 => -57,
    11121 => -57,
    11122 => -57,
    11123 => -57,
    11124 => -57,
    11125 => -57,
    11126 => -57,
    11127 => -57,
    11128 => -57,
    11129 => -57,
    11130 => -57,
    11131 => -57,
    11132 => -57,
    11133 => -57,
    11134 => -57,
    11135 => -57,
    11136 => -57,
    11137 => -57,
    11138 => -57,
    11139 => -57,
    11140 => -57,
    11141 => -57,
    11142 => -57,
    11143 => -57,
    11144 => -57,
    11145 => -57,
    11146 => -57,
    11147 => -57,
    11148 => -57,
    11149 => -57,
    11150 => -57,
    11151 => -57,
    11152 => -57,
    11153 => -57,
    11154 => -57,
    11155 => -57,
    11156 => -57,
    11157 => -57,
    11158 => -57,
    11159 => -57,
    11160 => -57,
    11161 => -57,
    11162 => -57,
    11163 => -57,
    11164 => -57,
    11165 => -57,
    11166 => -57,
    11167 => -57,
    11168 => -57,
    11169 => -57,
    11170 => -57,
    11171 => -57,
    11172 => -57,
    11173 => -57,
    11174 => -57,
    11175 => -57,
    11176 => -57,
    11177 => -57,
    11178 => -57,
    11179 => -57,
    11180 => -57,
    11181 => -57,
    11182 => -57,
    11183 => -57,
    11184 => -57,
    11185 => -57,
    11186 => -57,
    11187 => -57,
    11188 => -57,
    11189 => -57,
    11190 => -57,
    11191 => -58,
    11192 => -58,
    11193 => -58,
    11194 => -58,
    11195 => -58,
    11196 => -58,
    11197 => -58,
    11198 => -58,
    11199 => -58,
    11200 => -58,
    11201 => -58,
    11202 => -58,
    11203 => -58,
    11204 => -58,
    11205 => -58,
    11206 => -58,
    11207 => -58,
    11208 => -58,
    11209 => -58,
    11210 => -58,
    11211 => -58,
    11212 => -58,
    11213 => -58,
    11214 => -58,
    11215 => -58,
    11216 => -58,
    11217 => -58,
    11218 => -58,
    11219 => -58,
    11220 => -58,
    11221 => -58,
    11222 => -58,
    11223 => -58,
    11224 => -58,
    11225 => -58,
    11226 => -58,
    11227 => -58,
    11228 => -58,
    11229 => -58,
    11230 => -58,
    11231 => -58,
    11232 => -58,
    11233 => -58,
    11234 => -58,
    11235 => -58,
    11236 => -58,
    11237 => -58,
    11238 => -58,
    11239 => -58,
    11240 => -58,
    11241 => -58,
    11242 => -58,
    11243 => -58,
    11244 => -58,
    11245 => -58,
    11246 => -58,
    11247 => -58,
    11248 => -58,
    11249 => -58,
    11250 => -58,
    11251 => -58,
    11252 => -58,
    11253 => -58,
    11254 => -58,
    11255 => -58,
    11256 => -58,
    11257 => -58,
    11258 => -58,
    11259 => -58,
    11260 => -58,
    11261 => -58,
    11262 => -58,
    11263 => -58,
    11264 => -58,
    11265 => -58,
    11266 => -58,
    11267 => -58,
    11268 => -58,
    11269 => -58,
    11270 => -58,
    11271 => -58,
    11272 => -58,
    11273 => -58,
    11274 => -58,
    11275 => -58,
    11276 => -58,
    11277 => -58,
    11278 => -58,
    11279 => -58,
    11280 => -58,
    11281 => -58,
    11282 => -58,
    11283 => -58,
    11284 => -58,
    11285 => -58,
    11286 => -58,
    11287 => -58,
    11288 => -58,
    11289 => -58,
    11290 => -58,
    11291 => -58,
    11292 => -58,
    11293 => -58,
    11294 => -58,
    11295 => -58,
    11296 => -58,
    11297 => -59,
    11298 => -59,
    11299 => -59,
    11300 => -59,
    11301 => -59,
    11302 => -59,
    11303 => -59,
    11304 => -59,
    11305 => -59,
    11306 => -59,
    11307 => -59,
    11308 => -59,
    11309 => -59,
    11310 => -59,
    11311 => -59,
    11312 => -59,
    11313 => -59,
    11314 => -59,
    11315 => -59,
    11316 => -59,
    11317 => -59,
    11318 => -59,
    11319 => -59,
    11320 => -59,
    11321 => -59,
    11322 => -59,
    11323 => -59,
    11324 => -59,
    11325 => -59,
    11326 => -59,
    11327 => -59,
    11328 => -59,
    11329 => -59,
    11330 => -59,
    11331 => -59,
    11332 => -59,
    11333 => -59,
    11334 => -59,
    11335 => -59,
    11336 => -59,
    11337 => -59,
    11338 => -59,
    11339 => -59,
    11340 => -59,
    11341 => -59,
    11342 => -59,
    11343 => -59,
    11344 => -59,
    11345 => -59,
    11346 => -59,
    11347 => -59,
    11348 => -59,
    11349 => -59,
    11350 => -59,
    11351 => -59,
    11352 => -59,
    11353 => -59,
    11354 => -59,
    11355 => -59,
    11356 => -59,
    11357 => -59,
    11358 => -59,
    11359 => -59,
    11360 => -59,
    11361 => -59,
    11362 => -59,
    11363 => -59,
    11364 => -59,
    11365 => -59,
    11366 => -59,
    11367 => -59,
    11368 => -59,
    11369 => -59,
    11370 => -59,
    11371 => -59,
    11372 => -59,
    11373 => -59,
    11374 => -59,
    11375 => -59,
    11376 => -59,
    11377 => -59,
    11378 => -59,
    11379 => -59,
    11380 => -59,
    11381 => -59,
    11382 => -59,
    11383 => -59,
    11384 => -59,
    11385 => -59,
    11386 => -59,
    11387 => -59,
    11388 => -59,
    11389 => -59,
    11390 => -59,
    11391 => -59,
    11392 => -59,
    11393 => -59,
    11394 => -59,
    11395 => -59,
    11396 => -59,
    11397 => -59,
    11398 => -59,
    11399 => -59,
    11400 => -59,
    11401 => -59,
    11402 => -59,
    11403 => -59,
    11404 => -59,
    11405 => -59,
    11406 => -59,
    11407 => -59,
    11408 => -59,
    11409 => -59,
    11410 => -59,
    11411 => -59,
    11412 => -59,
    11413 => -59,
    11414 => -59,
    11415 => -60,
    11416 => -60,
    11417 => -60,
    11418 => -60,
    11419 => -60,
    11420 => -60,
    11421 => -60,
    11422 => -60,
    11423 => -60,
    11424 => -60,
    11425 => -60,
    11426 => -60,
    11427 => -60,
    11428 => -60,
    11429 => -60,
    11430 => -60,
    11431 => -60,
    11432 => -60,
    11433 => -60,
    11434 => -60,
    11435 => -60,
    11436 => -60,
    11437 => -60,
    11438 => -60,
    11439 => -60,
    11440 => -60,
    11441 => -60,
    11442 => -60,
    11443 => -60,
    11444 => -60,
    11445 => -60,
    11446 => -60,
    11447 => -60,
    11448 => -60,
    11449 => -60,
    11450 => -60,
    11451 => -60,
    11452 => -60,
    11453 => -60,
    11454 => -60,
    11455 => -60,
    11456 => -60,
    11457 => -60,
    11458 => -60,
    11459 => -60,
    11460 => -60,
    11461 => -60,
    11462 => -60,
    11463 => -60,
    11464 => -60,
    11465 => -60,
    11466 => -60,
    11467 => -60,
    11468 => -60,
    11469 => -60,
    11470 => -60,
    11471 => -60,
    11472 => -60,
    11473 => -60,
    11474 => -60,
    11475 => -60,
    11476 => -60,
    11477 => -60,
    11478 => -60,
    11479 => -60,
    11480 => -60,
    11481 => -60,
    11482 => -60,
    11483 => -60,
    11484 => -60,
    11485 => -60,
    11486 => -60,
    11487 => -60,
    11488 => -60,
    11489 => -60,
    11490 => -60,
    11491 => -60,
    11492 => -60,
    11493 => -60,
    11494 => -60,
    11495 => -60,
    11496 => -60,
    11497 => -60,
    11498 => -60,
    11499 => -60,
    11500 => -60,
    11501 => -60,
    11502 => -60,
    11503 => -60,
    11504 => -60,
    11505 => -60,
    11506 => -60,
    11507 => -60,
    11508 => -60,
    11509 => -60,
    11510 => -60,
    11511 => -60,
    11512 => -60,
    11513 => -60,
    11514 => -60,
    11515 => -60,
    11516 => -60,
    11517 => -60,
    11518 => -60,
    11519 => -60,
    11520 => -60,
    11521 => -60,
    11522 => -60,
    11523 => -60,
    11524 => -60,
    11525 => -60,
    11526 => -60,
    11527 => -60,
    11528 => -60,
    11529 => -60,
    11530 => -60,
    11531 => -60,
    11532 => -60,
    11533 => -60,
    11534 => -60,
    11535 => -60,
    11536 => -60,
    11537 => -60,
    11538 => -60,
    11539 => -60,
    11540 => -60,
    11541 => -60,
    11542 => -60,
    11543 => -60,
    11544 => -60,
    11545 => -60,
    11546 => -60,
    11547 => -60,
    11548 => -60,
    11549 => -60,
    11550 => -60,
    11551 => -61,
    11552 => -61,
    11553 => -61,
    11554 => -61,
    11555 => -61,
    11556 => -61,
    11557 => -61,
    11558 => -61,
    11559 => -61,
    11560 => -61,
    11561 => -61,
    11562 => -61,
    11563 => -61,
    11564 => -61,
    11565 => -61,
    11566 => -61,
    11567 => -61,
    11568 => -61,
    11569 => -61,
    11570 => -61,
    11571 => -61,
    11572 => -61,
    11573 => -61,
    11574 => -61,
    11575 => -61,
    11576 => -61,
    11577 => -61,
    11578 => -61,
    11579 => -61,
    11580 => -61,
    11581 => -61,
    11582 => -61,
    11583 => -61,
    11584 => -61,
    11585 => -61,
    11586 => -61,
    11587 => -61,
    11588 => -61,
    11589 => -61,
    11590 => -61,
    11591 => -61,
    11592 => -61,
    11593 => -61,
    11594 => -61,
    11595 => -61,
    11596 => -61,
    11597 => -61,
    11598 => -61,
    11599 => -61,
    11600 => -61,
    11601 => -61,
    11602 => -61,
    11603 => -61,
    11604 => -61,
    11605 => -61,
    11606 => -61,
    11607 => -61,
    11608 => -61,
    11609 => -61,
    11610 => -61,
    11611 => -61,
    11612 => -61,
    11613 => -61,
    11614 => -61,
    11615 => -61,
    11616 => -61,
    11617 => -61,
    11618 => -61,
    11619 => -61,
    11620 => -61,
    11621 => -61,
    11622 => -61,
    11623 => -61,
    11624 => -61,
    11625 => -61,
    11626 => -61,
    11627 => -61,
    11628 => -61,
    11629 => -61,
    11630 => -61,
    11631 => -61,
    11632 => -61,
    11633 => -61,
    11634 => -61,
    11635 => -61,
    11636 => -61,
    11637 => -61,
    11638 => -61,
    11639 => -61,
    11640 => -61,
    11641 => -61,
    11642 => -61,
    11643 => -61,
    11644 => -61,
    11645 => -61,
    11646 => -61,
    11647 => -61,
    11648 => -61,
    11649 => -61,
    11650 => -61,
    11651 => -61,
    11652 => -61,
    11653 => -61,
    11654 => -61,
    11655 => -61,
    11656 => -61,
    11657 => -61,
    11658 => -61,
    11659 => -61,
    11660 => -61,
    11661 => -61,
    11662 => -61,
    11663 => -61,
    11664 => -61,
    11665 => -61,
    11666 => -61,
    11667 => -61,
    11668 => -61,
    11669 => -61,
    11670 => -61,
    11671 => -61,
    11672 => -61,
    11673 => -61,
    11674 => -61,
    11675 => -61,
    11676 => -61,
    11677 => -61,
    11678 => -61,
    11679 => -61,
    11680 => -61,
    11681 => -61,
    11682 => -61,
    11683 => -61,
    11684 => -61,
    11685 => -61,
    11686 => -61,
    11687 => -61,
    11688 => -61,
    11689 => -61,
    11690 => -61,
    11691 => -61,
    11692 => -61,
    11693 => -61,
    11694 => -61,
    11695 => -61,
    11696 => -61,
    11697 => -61,
    11698 => -61,
    11699 => -61,
    11700 => -61,
    11701 => -61,
    11702 => -61,
    11703 => -61,
    11704 => -61,
    11705 => -61,
    11706 => -61,
    11707 => -61,
    11708 => -61,
    11709 => -61,
    11710 => -61,
    11711 => -61,
    11712 => -61,
    11713 => -61,
    11714 => -61,
    11715 => -61,
    11716 => -61,
    11717 => -61,
    11718 => -62,
    11719 => -62,
    11720 => -62,
    11721 => -62,
    11722 => -62,
    11723 => -62,
    11724 => -62,
    11725 => -62,
    11726 => -62,
    11727 => -62,
    11728 => -62,
    11729 => -62,
    11730 => -62,
    11731 => -62,
    11732 => -62,
    11733 => -62,
    11734 => -62,
    11735 => -62,
    11736 => -62,
    11737 => -62,
    11738 => -62,
    11739 => -62,
    11740 => -62,
    11741 => -62,
    11742 => -62,
    11743 => -62,
    11744 => -62,
    11745 => -62,
    11746 => -62,
    11747 => -62,
    11748 => -62,
    11749 => -62,
    11750 => -62,
    11751 => -62,
    11752 => -62,
    11753 => -62,
    11754 => -62,
    11755 => -62,
    11756 => -62,
    11757 => -62,
    11758 => -62,
    11759 => -62,
    11760 => -62,
    11761 => -62,
    11762 => -62,
    11763 => -62,
    11764 => -62,
    11765 => -62,
    11766 => -62,
    11767 => -62,
    11768 => -62,
    11769 => -62,
    11770 => -62,
    11771 => -62,
    11772 => -62,
    11773 => -62,
    11774 => -62,
    11775 => -62,
    11776 => -62,
    11777 => -62,
    11778 => -62,
    11779 => -62,
    11780 => -62,
    11781 => -62,
    11782 => -62,
    11783 => -62,
    11784 => -62,
    11785 => -62,
    11786 => -62,
    11787 => -62,
    11788 => -62,
    11789 => -62,
    11790 => -62,
    11791 => -62,
    11792 => -62,
    11793 => -62,
    11794 => -62,
    11795 => -62,
    11796 => -62,
    11797 => -62,
    11798 => -62,
    11799 => -62,
    11800 => -62,
    11801 => -62,
    11802 => -62,
    11803 => -62,
    11804 => -62,
    11805 => -62,
    11806 => -62,
    11807 => -62,
    11808 => -62,
    11809 => -62,
    11810 => -62,
    11811 => -62,
    11812 => -62,
    11813 => -62,
    11814 => -62,
    11815 => -62,
    11816 => -62,
    11817 => -62,
    11818 => -62,
    11819 => -62,
    11820 => -62,
    11821 => -62,
    11822 => -62,
    11823 => -62,
    11824 => -62,
    11825 => -62,
    11826 => -62,
    11827 => -62,
    11828 => -62,
    11829 => -62,
    11830 => -62,
    11831 => -62,
    11832 => -62,
    11833 => -62,
    11834 => -62,
    11835 => -62,
    11836 => -62,
    11837 => -62,
    11838 => -62,
    11839 => -62,
    11840 => -62,
    11841 => -62,
    11842 => -62,
    11843 => -62,
    11844 => -62,
    11845 => -62,
    11846 => -62,
    11847 => -62,
    11848 => -62,
    11849 => -62,
    11850 => -62,
    11851 => -62,
    11852 => -62,
    11853 => -62,
    11854 => -62,
    11855 => -62,
    11856 => -62,
    11857 => -62,
    11858 => -62,
    11859 => -62,
    11860 => -62,
    11861 => -62,
    11862 => -62,
    11863 => -62,
    11864 => -62,
    11865 => -62,
    11866 => -62,
    11867 => -62,
    11868 => -62,
    11869 => -62,
    11870 => -62,
    11871 => -62,
    11872 => -62,
    11873 => -62,
    11874 => -62,
    11875 => -62,
    11876 => -62,
    11877 => -62,
    11878 => -62,
    11879 => -62,
    11880 => -62,
    11881 => -62,
    11882 => -62,
    11883 => -62,
    11884 => -62,
    11885 => -62,
    11886 => -62,
    11887 => -62,
    11888 => -62,
    11889 => -62,
    11890 => -62,
    11891 => -62,
    11892 => -62,
    11893 => -62,
    11894 => -62,
    11895 => -62,
    11896 => -62,
    11897 => -62,
    11898 => -62,
    11899 => -62,
    11900 => -62,
    11901 => -62,
    11902 => -62,
    11903 => -62,
    11904 => -62,
    11905 => -62,
    11906 => -62,
    11907 => -62,
    11908 => -62,
    11909 => -62,
    11910 => -62,
    11911 => -62,
    11912 => -62,
    11913 => -62,
    11914 => -62,
    11915 => -62,
    11916 => -62,
    11917 => -62,
    11918 => -62,
    11919 => -62,
    11920 => -62,
    11921 => -62,
    11922 => -62,
    11923 => -62,
    11924 => -62,
    11925 => -62,
    11926 => -62,
    11927 => -62,
    11928 => -62,
    11929 => -62,
    11930 => -62,
    11931 => -62,
    11932 => -62,
    11933 => -62,
    11934 => -62,
    11935 => -62,
    11936 => -62,
    11937 => -62,
    11938 => -62,
    11939 => -62,
    11940 => -62,
    11941 => -62,
    11942 => -62,
    11943 => -62,
    11944 => -62,
    11945 => -62,
    11946 => -62,
    11947 => -62,
    11948 => -62,
    11949 => -62,
    11950 => -62,
    11951 => -62,
    11952 => -62,
    11953 => -62,
    11954 => -62,
    11955 => -62,
    11956 => -62,
    11957 => -62,
    11958 => -62,
    11959 => -62,
    11960 => -63,
    11961 => -63,
    11962 => -63,
    11963 => -63,
    11964 => -63,
    11965 => -63,
    11966 => -63,
    11967 => -63,
    11968 => -63,
    11969 => -63,
    11970 => -63,
    11971 => -63,
    11972 => -63,
    11973 => -63,
    11974 => -63,
    11975 => -63,
    11976 => -63,
    11977 => -63,
    11978 => -63,
    11979 => -63,
    11980 => -63,
    11981 => -63,
    11982 => -63,
    11983 => -63,
    11984 => -63,
    11985 => -63,
    11986 => -63,
    11987 => -63,
    11988 => -63,
    11989 => -63,
    11990 => -63,
    11991 => -63,
    11992 => -63,
    11993 => -63,
    11994 => -63,
    11995 => -63,
    11996 => -63,
    11997 => -63,
    11998 => -63,
    11999 => -63,
    12000 => -63,
    12001 => -63,
    12002 => -63,
    12003 => -63,
    12004 => -63,
    12005 => -63,
    12006 => -63,
    12007 => -63,
    12008 => -63,
    12009 => -63,
    12010 => -63,
    12011 => -63,
    12012 => -63,
    12013 => -63,
    12014 => -63,
    12015 => -63,
    12016 => -63,
    12017 => -63,
    12018 => -63,
    12019 => -63,
    12020 => -63,
    12021 => -63,
    12022 => -63,
    12023 => -63,
    12024 => -63,
    12025 => -63,
    12026 => -63,
    12027 => -63,
    12028 => -63,
    12029 => -63,
    12030 => -63,
    12031 => -63,
    12032 => -63,
    12033 => -63,
    12034 => -63,
    12035 => -63,
    12036 => -63,
    12037 => -63,
    12038 => -63,
    12039 => -63,
    12040 => -63,
    12041 => -63,
    12042 => -63,
    12043 => -63,
    12044 => -63,
    12045 => -63,
    12046 => -63,
    12047 => -63,
    12048 => -63,
    12049 => -63,
    12050 => -63,
    12051 => -63,
    12052 => -63,
    12053 => -63,
    12054 => -63,
    12055 => -63,
    12056 => -63,
    12057 => -63,
    12058 => -63,
    12059 => -63,
    12060 => -63,
    12061 => -63,
    12062 => -63,
    12063 => -63,
    12064 => -63,
    12065 => -63,
    12066 => -63,
    12067 => -63,
    12068 => -63,
    12069 => -63,
    12070 => -63,
    12071 => -63,
    12072 => -63,
    12073 => -63,
    12074 => -63,
    12075 => -63,
    12076 => -63,
    12077 => -63,
    12078 => -63,
    12079 => -63,
    12080 => -63,
    12081 => -63,
    12082 => -63,
    12083 => -63,
    12084 => -63,
    12085 => -63,
    12086 => -63,
    12087 => -63,
    12088 => -63,
    12089 => -63,
    12090 => -63,
    12091 => -63,
    12092 => -63,
    12093 => -63,
    12094 => -63,
    12095 => -63,
    12096 => -63,
    12097 => -63,
    12098 => -63,
    12099 => -63,
    12100 => -63,
    12101 => -63,
    12102 => -63,
    12103 => -63,
    12104 => -63,
    12105 => -63,
    12106 => -63,
    12107 => -63,
    12108 => -63,
    12109 => -63,
    12110 => -63,
    12111 => -63,
    12112 => -63,
    12113 => -63,
    12114 => -63,
    12115 => -63,
    12116 => -63,
    12117 => -63,
    12118 => -63,
    12119 => -63,
    12120 => -63,
    12121 => -63,
    12122 => -63,
    12123 => -63,
    12124 => -63,
    12125 => -63,
    12126 => -63,
    12127 => -63,
    12128 => -63,
    12129 => -63,
    12130 => -63,
    12131 => -63,
    12132 => -63,
    12133 => -63,
    12134 => -63,
    12135 => -63,
    12136 => -63,
    12137 => -63,
    12138 => -63,
    12139 => -63,
    12140 => -63,
    12141 => -63,
    12142 => -63,
    12143 => -63,
    12144 => -63,
    12145 => -63,
    12146 => -63,
    12147 => -63,
    12148 => -63,
    12149 => -63,
    12150 => -63,
    12151 => -63,
    12152 => -63,
    12153 => -63,
    12154 => -63,
    12155 => -63,
    12156 => -63,
    12157 => -63,
    12158 => -63,
    12159 => -63,
    12160 => -63,
    12161 => -63,
    12162 => -63,
    12163 => -63,
    12164 => -63,
    12165 => -63,
    12166 => -63,
    12167 => -63,
    12168 => -63,
    12169 => -63,
    12170 => -63,
    12171 => -63,
    12172 => -63,
    12173 => -63,
    12174 => -63,
    12175 => -63,
    12176 => -63,
    12177 => -63,
    12178 => -63,
    12179 => -63,
    12180 => -63,
    12181 => -63,
    12182 => -63,
    12183 => -63,
    12184 => -63,
    12185 => -63,
    12186 => -63,
    12187 => -63,
    12188 => -63,
    12189 => -63,
    12190 => -63,
    12191 => -63,
    12192 => -63,
    12193 => -63,
    12194 => -63,
    12195 => -63,
    12196 => -63,
    12197 => -63,
    12198 => -63,
    12199 => -63,
    12200 => -63,
    12201 => -63,
    12202 => -63,
    12203 => -63,
    12204 => -63,
    12205 => -63,
    12206 => -63,
    12207 => -63,
    12208 => -63,
    12209 => -63,
    12210 => -63,
    12211 => -63,
    12212 => -63,
    12213 => -63,
    12214 => -63,
    12215 => -63,
    12216 => -63,
    12217 => -63,
    12218 => -63,
    12219 => -63,
    12220 => -63,
    12221 => -63,
    12222 => -63,
    12223 => -63,
    12224 => -63,
    12225 => -63,
    12226 => -63,
    12227 => -63,
    12228 => -63,
    12229 => -63,
    12230 => -63,
    12231 => -63,
    12232 => -63,
    12233 => -63,
    12234 => -63,
    12235 => -63,
    12236 => -63,
    12237 => -63,
    12238 => -63,
    12239 => -63,
    12240 => -63,
    12241 => -63,
    12242 => -63,
    12243 => -63,
    12244 => -63,
    12245 => -63,
    12246 => -63,
    12247 => -63,
    12248 => -63,
    12249 => -63,
    12250 => -63,
    12251 => -63,
    12252 => -63,
    12253 => -63,
    12254 => -63,
    12255 => -63,
    12256 => -63,
    12257 => -63,
    12258 => -63,
    12259 => -63,
    12260 => -63,
    12261 => -63,
    12262 => -63,
    12263 => -63,
    12264 => -63,
    12265 => -63,
    12266 => -63,
    12267 => -63,
    12268 => -63,
    12269 => -63,
    12270 => -63,
    12271 => -63,
    12272 => -63,
    12273 => -63,
    12274 => -63,
    12275 => -63,
    12276 => -63,
    12277 => -63,
    12278 => -63,
    12279 => -63,
    12280 => -63,
    12281 => -63,
    12282 => -63,
    12283 => -63,
    12284 => -63,
    12285 => -63,
    12286 => -63,
    12287 => -63,
    12288 => -63,
    12289 => -63,
    12290 => -63,
    12291 => -63,
    12292 => -63,
    12293 => -63,
    12294 => -63,
    12295 => -63,
    12296 => -63,
    12297 => -63,
    12298 => -63,
    12299 => -63,
    12300 => -63,
    12301 => -63,
    12302 => -63,
    12303 => -63,
    12304 => -63,
    12305 => -63,
    12306 => -63,
    12307 => -63,
    12308 => -63,
    12309 => -63,
    12310 => -63,
    12311 => -63,
    12312 => -63,
    12313 => -63,
    12314 => -63,
    12315 => -63,
    12316 => -63,
    12317 => -63,
    12318 => -63,
    12319 => -63,
    12320 => -63,
    12321 => -63,
    12322 => -63,
    12323 => -63,
    12324 => -63,
    12325 => -63,
    12326 => -63,
    12327 => -63,
    12328 => -63,
    12329 => -63,
    12330 => -63,
    12331 => -63,
    12332 => -63,
    12333 => -63,
    12334 => -63,
    12335 => -63,
    12336 => -63,
    12337 => -63,
    12338 => -63,
    12339 => -63,
    12340 => -63,
    12341 => -63,
    12342 => -63,
    12343 => -63,
    12344 => -63,
    12345 => -63,
    12346 => -63,
    12347 => -63,
    12348 => -63,
    12349 => -63,
    12350 => -63,
    12351 => -63,
    12352 => -63,
    12353 => -63,
    12354 => -63,
    12355 => -63,
    12356 => -63,
    12357 => -63,
    12358 => -63,
    12359 => -63,
    12360 => -63,
    12361 => -63,
    12362 => -63,
    12363 => -63,
    12364 => -63,
    12365 => -63,
    12366 => -63,
    12367 => -63,
    12368 => -63,
    12369 => -63,
    12370 => -63,
    12371 => -63,
    12372 => -63,
    12373 => -63,
    12374 => -63,
    12375 => -63,
    12376 => -63,
    12377 => -63,
    12378 => -63,
    12379 => -63,
    12380 => -63,
    12381 => -63,
    12382 => -63,
    12383 => -63,
    12384 => -63,
    12385 => -63,
    12386 => -63,
    12387 => -63,
    12388 => -63,
    12389 => -63,
    12390 => -63,
    12391 => -63,
    12392 => -63,
    12393 => -63,
    12394 => -63,
    12395 => -63,
    12396 => -63,
    12397 => -63,
    12398 => -63,
    12399 => -63,
    12400 => -63,
    12401 => -63,
    12402 => -63,
    12403 => -63,
    12404 => -63,
    12405 => -63,
    12406 => -63,
    12407 => -63,
    12408 => -63,
    12409 => -63,
    12410 => -63,
    12411 => -63,
    12412 => -63,
    12413 => -63,
    12414 => -63,
    12415 => -63,
    12416 => -63,
    12417 => -63,
    12418 => -63,
    12419 => -63,
    12420 => -63,
    12421 => -63,
    12422 => -63,
    12423 => -63,
    12424 => -63,
    12425 => -63,
    12426 => -63,
    12427 => -63,
    12428 => -63,
    12429 => -63,
    12430 => -63,
    12431 => -63,
    12432 => -63,
    12433 => -63,
    12434 => -63,
    12435 => -63,
    12436 => -63,
    12437 => -63,
    12438 => -63,
    12439 => -63,
    12440 => -63,
    12441 => -63,
    12442 => -63,
    12443 => -63,
    12444 => -63,
    12445 => -63,
    12446 => -63,
    12447 => -63,
    12448 => -63,
    12449 => -63,
    12450 => -63,
    12451 => -63,
    12452 => -63,
    12453 => -63,
    12454 => -63,
    12455 => -63,
    12456 => -63,
    12457 => -63,
    12458 => -63,
    12459 => -63,
    12460 => -63,
    12461 => -63,
    12462 => -63,
    12463 => -63,
    12464 => -63,
    12465 => -63,
    12466 => -63,
    12467 => -63,
    12468 => -63,
    12469 => -63,
    12470 => -63,
    12471 => -63,
    12472 => -63,
    12473 => -63,
    12474 => -63,
    12475 => -63,
    12476 => -63,
    12477 => -63,
    12478 => -63,
    12479 => -63,
    12480 => -63,
    12481 => -63,
    12482 => -63,
    12483 => -63,
    12484 => -63,
    12485 => -63,
    12486 => -63,
    12487 => -63,
    12488 => -63,
    12489 => -63,
    12490 => -63,
    12491 => -63,
    12492 => -63,
    12493 => -63,
    12494 => -63,
    12495 => -63,
    12496 => -63,
    12497 => -63,
    12498 => -63,
    12499 => -63,
    12500 => -63,
    12501 => -63,
    12502 => -63,
    12503 => -63,
    12504 => -63,
    12505 => -63,
    12506 => -63,
    12507 => -63,
    12508 => -63,
    12509 => -63,
    12510 => -63,
    12511 => -63,
    12512 => -63,
    12513 => -63,
    12514 => -63,
    12515 => -63,
    12516 => -63,
    12517 => -63,
    12518 => -63,
    12519 => -63,
    12520 => -63,
    12521 => -63,
    12522 => -63,
    12523 => -63,
    12524 => -63,
    12525 => -63,
    12526 => -63,
    12527 => -63,
    12528 => -63,
    12529 => -63,
    12530 => -63,
    12531 => -63,
    12532 => -63,
    12533 => -63,
    12534 => -63,
    12535 => -63,
    12536 => -63,
    12537 => -63,
    12538 => -63,
    12539 => -63,
    12540 => -63,
    12541 => -63,
    12542 => -63,
    12543 => -63,
    12544 => -63,
    12545 => -63,
    12546 => -63,
    12547 => -63,
    12548 => -63,
    12549 => -63,
    12550 => -63,
    12551 => -63,
    12552 => -63,
    12553 => -63,
    12554 => -63,
    12555 => -63,
    12556 => -63,
    12557 => -63,
    12558 => -63,
    12559 => -63,
    12560 => -63,
    12561 => -63,
    12562 => -63,
    12563 => -63,
    12564 => -63,
    12565 => -63,
    12566 => -63,
    12567 => -63,
    12568 => -63,
    12569 => -63,
    12570 => -63,
    12571 => -63,
    12572 => -63,
    12573 => -63,
    12574 => -63,
    12575 => -63,
    12576 => -63,
    12577 => -63,
    12578 => -63,
    12579 => -63,
    12580 => -63,
    12581 => -63,
    12582 => -63,
    12583 => -63,
    12584 => -63,
    12585 => -63,
    12586 => -63,
    12587 => -63,
    12588 => -63,
    12589 => -63,
    12590 => -63,
    12591 => -63,
    12592 => -63,
    12593 => -63,
    12594 => -63,
    12595 => -63,
    12596 => -63,
    12597 => -63,
    12598 => -63,
    12599 => -63,
    12600 => -63,
    12601 => -63,
    12602 => -63,
    12603 => -63,
    12604 => -63,
    12605 => -63,
    12606 => -63,
    12607 => -63,
    12608 => -63,
    12609 => -63,
    12610 => -63,
    12611 => -63,
    12612 => -63,
    12613 => -63,
    12614 => -63,
    12615 => -63,
    12616 => -63,
    12617 => -62,
    12618 => -62,
    12619 => -62,
    12620 => -62,
    12621 => -62,
    12622 => -62,
    12623 => -62,
    12624 => -62,
    12625 => -62,
    12626 => -62,
    12627 => -62,
    12628 => -62,
    12629 => -62,
    12630 => -62,
    12631 => -62,
    12632 => -62,
    12633 => -62,
    12634 => -62,
    12635 => -62,
    12636 => -62,
    12637 => -62,
    12638 => -62,
    12639 => -62,
    12640 => -62,
    12641 => -62,
    12642 => -62,
    12643 => -62,
    12644 => -62,
    12645 => -62,
    12646 => -62,
    12647 => -62,
    12648 => -62,
    12649 => -62,
    12650 => -62,
    12651 => -62,
    12652 => -62,
    12653 => -62,
    12654 => -62,
    12655 => -62,
    12656 => -62,
    12657 => -62,
    12658 => -62,
    12659 => -62,
    12660 => -62,
    12661 => -62,
    12662 => -62,
    12663 => -62,
    12664 => -62,
    12665 => -62,
    12666 => -62,
    12667 => -62,
    12668 => -62,
    12669 => -62,
    12670 => -62,
    12671 => -62,
    12672 => -62,
    12673 => -62,
    12674 => -62,
    12675 => -62,
    12676 => -62,
    12677 => -62,
    12678 => -62,
    12679 => -62,
    12680 => -62,
    12681 => -62,
    12682 => -62,
    12683 => -62,
    12684 => -62,
    12685 => -62,
    12686 => -62,
    12687 => -62,
    12688 => -62,
    12689 => -62,
    12690 => -62,
    12691 => -62,
    12692 => -62,
    12693 => -62,
    12694 => -62,
    12695 => -62,
    12696 => -62,
    12697 => -62,
    12698 => -62,
    12699 => -62,
    12700 => -62,
    12701 => -62,
    12702 => -62,
    12703 => -62,
    12704 => -62,
    12705 => -62,
    12706 => -62,
    12707 => -62,
    12708 => -62,
    12709 => -62,
    12710 => -62,
    12711 => -62,
    12712 => -62,
    12713 => -62,
    12714 => -62,
    12715 => -62,
    12716 => -62,
    12717 => -62,
    12718 => -62,
    12719 => -62,
    12720 => -62,
    12721 => -62,
    12722 => -62,
    12723 => -62,
    12724 => -62,
    12725 => -62,
    12726 => -62,
    12727 => -62,
    12728 => -62,
    12729 => -62,
    12730 => -62,
    12731 => -62,
    12732 => -62,
    12733 => -62,
    12734 => -62,
    12735 => -62,
    12736 => -62,
    12737 => -62,
    12738 => -62,
    12739 => -62,
    12740 => -62,
    12741 => -62,
    12742 => -62,
    12743 => -62,
    12744 => -62,
    12745 => -62,
    12746 => -62,
    12747 => -62,
    12748 => -62,
    12749 => -62,
    12750 => -62,
    12751 => -62,
    12752 => -62,
    12753 => -62,
    12754 => -62,
    12755 => -62,
    12756 => -62,
    12757 => -62,
    12758 => -62,
    12759 => -62,
    12760 => -62,
    12761 => -62,
    12762 => -62,
    12763 => -62,
    12764 => -62,
    12765 => -62,
    12766 => -62,
    12767 => -62,
    12768 => -62,
    12769 => -62,
    12770 => -62,
    12771 => -62,
    12772 => -62,
    12773 => -62,
    12774 => -62,
    12775 => -62,
    12776 => -62,
    12777 => -62,
    12778 => -62,
    12779 => -62,
    12780 => -62,
    12781 => -62,
    12782 => -62,
    12783 => -62,
    12784 => -62,
    12785 => -62,
    12786 => -62,
    12787 => -62,
    12788 => -62,
    12789 => -62,
    12790 => -62,
    12791 => -62,
    12792 => -62,
    12793 => -62,
    12794 => -62,
    12795 => -62,
    12796 => -62,
    12797 => -62,
    12798 => -62,
    12799 => -62,
    12800 => -62,
    12801 => -62,
    12802 => -62,
    12803 => -62,
    12804 => -62,
    12805 => -62,
    12806 => -62,
    12807 => -62,
    12808 => -62,
    12809 => -62,
    12810 => -62,
    12811 => -62,
    12812 => -62,
    12813 => -62,
    12814 => -62,
    12815 => -62,
    12816 => -62,
    12817 => -62,
    12818 => -62,
    12819 => -62,
    12820 => -62,
    12821 => -62,
    12822 => -62,
    12823 => -62,
    12824 => -62,
    12825 => -62,
    12826 => -62,
    12827 => -62,
    12828 => -62,
    12829 => -62,
    12830 => -62,
    12831 => -62,
    12832 => -62,
    12833 => -62,
    12834 => -62,
    12835 => -62,
    12836 => -62,
    12837 => -62,
    12838 => -62,
    12839 => -62,
    12840 => -62,
    12841 => -62,
    12842 => -62,
    12843 => -62,
    12844 => -62,
    12845 => -62,
    12846 => -62,
    12847 => -62,
    12848 => -62,
    12849 => -62,
    12850 => -62,
    12851 => -62,
    12852 => -62,
    12853 => -62,
    12854 => -62,
    12855 => -62,
    12856 => -62,
    12857 => -62,
    12858 => -62,
    12859 => -61,
    12860 => -61,
    12861 => -61,
    12862 => -61,
    12863 => -61,
    12864 => -61,
    12865 => -61,
    12866 => -61,
    12867 => -61,
    12868 => -61,
    12869 => -61,
    12870 => -61,
    12871 => -61,
    12872 => -61,
    12873 => -61,
    12874 => -61,
    12875 => -61,
    12876 => -61,
    12877 => -61,
    12878 => -61,
    12879 => -61,
    12880 => -61,
    12881 => -61,
    12882 => -61,
    12883 => -61,
    12884 => -61,
    12885 => -61,
    12886 => -61,
    12887 => -61,
    12888 => -61,
    12889 => -61,
    12890 => -61,
    12891 => -61,
    12892 => -61,
    12893 => -61,
    12894 => -61,
    12895 => -61,
    12896 => -61,
    12897 => -61,
    12898 => -61,
    12899 => -61,
    12900 => -61,
    12901 => -61,
    12902 => -61,
    12903 => -61,
    12904 => -61,
    12905 => -61,
    12906 => -61,
    12907 => -61,
    12908 => -61,
    12909 => -61,
    12910 => -61,
    12911 => -61,
    12912 => -61,
    12913 => -61,
    12914 => -61,
    12915 => -61,
    12916 => -61,
    12917 => -61,
    12918 => -61,
    12919 => -61,
    12920 => -61,
    12921 => -61,
    12922 => -61,
    12923 => -61,
    12924 => -61,
    12925 => -61,
    12926 => -61,
    12927 => -61,
    12928 => -61,
    12929 => -61,
    12930 => -61,
    12931 => -61,
    12932 => -61,
    12933 => -61,
    12934 => -61,
    12935 => -61,
    12936 => -61,
    12937 => -61,
    12938 => -61,
    12939 => -61,
    12940 => -61,
    12941 => -61,
    12942 => -61,
    12943 => -61,
    12944 => -61,
    12945 => -61,
    12946 => -61,
    12947 => -61,
    12948 => -61,
    12949 => -61,
    12950 => -61,
    12951 => -61,
    12952 => -61,
    12953 => -61,
    12954 => -61,
    12955 => -61,
    12956 => -61,
    12957 => -61,
    12958 => -61,
    12959 => -61,
    12960 => -61,
    12961 => -61,
    12962 => -61,
    12963 => -61,
    12964 => -61,
    12965 => -61,
    12966 => -61,
    12967 => -61,
    12968 => -61,
    12969 => -61,
    12970 => -61,
    12971 => -61,
    12972 => -61,
    12973 => -61,
    12974 => -61,
    12975 => -61,
    12976 => -61,
    12977 => -61,
    12978 => -61,
    12979 => -61,
    12980 => -61,
    12981 => -61,
    12982 => -61,
    12983 => -61,
    12984 => -61,
    12985 => -61,
    12986 => -61,
    12987 => -61,
    12988 => -61,
    12989 => -61,
    12990 => -61,
    12991 => -61,
    12992 => -61,
    12993 => -61,
    12994 => -61,
    12995 => -61,
    12996 => -61,
    12997 => -61,
    12998 => -61,
    12999 => -61,
    13000 => -61,
    13001 => -61,
    13002 => -61,
    13003 => -61,
    13004 => -61,
    13005 => -61,
    13006 => -61,
    13007 => -61,
    13008 => -61,
    13009 => -61,
    13010 => -61,
    13011 => -61,
    13012 => -61,
    13013 => -61,
    13014 => -61,
    13015 => -61,
    13016 => -61,
    13017 => -61,
    13018 => -61,
    13019 => -61,
    13020 => -61,
    13021 => -61,
    13022 => -61,
    13023 => -61,
    13024 => -61,
    13025 => -61,
    13026 => -60,
    13027 => -60,
    13028 => -60,
    13029 => -60,
    13030 => -60,
    13031 => -60,
    13032 => -60,
    13033 => -60,
    13034 => -60,
    13035 => -60,
    13036 => -60,
    13037 => -60,
    13038 => -60,
    13039 => -60,
    13040 => -60,
    13041 => -60,
    13042 => -60,
    13043 => -60,
    13044 => -60,
    13045 => -60,
    13046 => -60,
    13047 => -60,
    13048 => -60,
    13049 => -60,
    13050 => -60,
    13051 => -60,
    13052 => -60,
    13053 => -60,
    13054 => -60,
    13055 => -60,
    13056 => -60,
    13057 => -60,
    13058 => -60,
    13059 => -60,
    13060 => -60,
    13061 => -60,
    13062 => -60,
    13063 => -60,
    13064 => -60,
    13065 => -60,
    13066 => -60,
    13067 => -60,
    13068 => -60,
    13069 => -60,
    13070 => -60,
    13071 => -60,
    13072 => -60,
    13073 => -60,
    13074 => -60,
    13075 => -60,
    13076 => -60,
    13077 => -60,
    13078 => -60,
    13079 => -60,
    13080 => -60,
    13081 => -60,
    13082 => -60,
    13083 => -60,
    13084 => -60,
    13085 => -60,
    13086 => -60,
    13087 => -60,
    13088 => -60,
    13089 => -60,
    13090 => -60,
    13091 => -60,
    13092 => -60,
    13093 => -60,
    13094 => -60,
    13095 => -60,
    13096 => -60,
    13097 => -60,
    13098 => -60,
    13099 => -60,
    13100 => -60,
    13101 => -60,
    13102 => -60,
    13103 => -60,
    13104 => -60,
    13105 => -60,
    13106 => -60,
    13107 => -60,
    13108 => -60,
    13109 => -60,
    13110 => -60,
    13111 => -60,
    13112 => -60,
    13113 => -60,
    13114 => -60,
    13115 => -60,
    13116 => -60,
    13117 => -60,
    13118 => -60,
    13119 => -60,
    13120 => -60,
    13121 => -60,
    13122 => -60,
    13123 => -60,
    13124 => -60,
    13125 => -60,
    13126 => -60,
    13127 => -60,
    13128 => -60,
    13129 => -60,
    13130 => -60,
    13131 => -60,
    13132 => -60,
    13133 => -60,
    13134 => -60,
    13135 => -60,
    13136 => -60,
    13137 => -60,
    13138 => -60,
    13139 => -60,
    13140 => -60,
    13141 => -60,
    13142 => -60,
    13143 => -60,
    13144 => -60,
    13145 => -60,
    13146 => -60,
    13147 => -60,
    13148 => -60,
    13149 => -60,
    13150 => -60,
    13151 => -60,
    13152 => -60,
    13153 => -60,
    13154 => -60,
    13155 => -60,
    13156 => -60,
    13157 => -60,
    13158 => -60,
    13159 => -60,
    13160 => -60,
    13161 => -60,
    13162 => -59,
    13163 => -59,
    13164 => -59,
    13165 => -59,
    13166 => -59,
    13167 => -59,
    13168 => -59,
    13169 => -59,
    13170 => -59,
    13171 => -59,
    13172 => -59,
    13173 => -59,
    13174 => -59,
    13175 => -59,
    13176 => -59,
    13177 => -59,
    13178 => -59,
    13179 => -59,
    13180 => -59,
    13181 => -59,
    13182 => -59,
    13183 => -59,
    13184 => -59,
    13185 => -59,
    13186 => -59,
    13187 => -59,
    13188 => -59,
    13189 => -59,
    13190 => -59,
    13191 => -59,
    13192 => -59,
    13193 => -59,
    13194 => -59,
    13195 => -59,
    13196 => -59,
    13197 => -59,
    13198 => -59,
    13199 => -59,
    13200 => -59,
    13201 => -59,
    13202 => -59,
    13203 => -59,
    13204 => -59,
    13205 => -59,
    13206 => -59,
    13207 => -59,
    13208 => -59,
    13209 => -59,
    13210 => -59,
    13211 => -59,
    13212 => -59,
    13213 => -59,
    13214 => -59,
    13215 => -59,
    13216 => -59,
    13217 => -59,
    13218 => -59,
    13219 => -59,
    13220 => -59,
    13221 => -59,
    13222 => -59,
    13223 => -59,
    13224 => -59,
    13225 => -59,
    13226 => -59,
    13227 => -59,
    13228 => -59,
    13229 => -59,
    13230 => -59,
    13231 => -59,
    13232 => -59,
    13233 => -59,
    13234 => -59,
    13235 => -59,
    13236 => -59,
    13237 => -59,
    13238 => -59,
    13239 => -59,
    13240 => -59,
    13241 => -59,
    13242 => -59,
    13243 => -59,
    13244 => -59,
    13245 => -59,
    13246 => -59,
    13247 => -59,
    13248 => -59,
    13249 => -59,
    13250 => -59,
    13251 => -59,
    13252 => -59,
    13253 => -59,
    13254 => -59,
    13255 => -59,
    13256 => -59,
    13257 => -59,
    13258 => -59,
    13259 => -59,
    13260 => -59,
    13261 => -59,
    13262 => -59,
    13263 => -59,
    13264 => -59,
    13265 => -59,
    13266 => -59,
    13267 => -59,
    13268 => -59,
    13269 => -59,
    13270 => -59,
    13271 => -59,
    13272 => -59,
    13273 => -59,
    13274 => -59,
    13275 => -59,
    13276 => -59,
    13277 => -59,
    13278 => -59,
    13279 => -59,
    13280 => -58,
    13281 => -58,
    13282 => -58,
    13283 => -58,
    13284 => -58,
    13285 => -58,
    13286 => -58,
    13287 => -58,
    13288 => -58,
    13289 => -58,
    13290 => -58,
    13291 => -58,
    13292 => -58,
    13293 => -58,
    13294 => -58,
    13295 => -58,
    13296 => -58,
    13297 => -58,
    13298 => -58,
    13299 => -58,
    13300 => -58,
    13301 => -58,
    13302 => -58,
    13303 => -58,
    13304 => -58,
    13305 => -58,
    13306 => -58,
    13307 => -58,
    13308 => -58,
    13309 => -58,
    13310 => -58,
    13311 => -58,
    13312 => -58,
    13313 => -58,
    13314 => -58,
    13315 => -58,
    13316 => -58,
    13317 => -58,
    13318 => -58,
    13319 => -58,
    13320 => -58,
    13321 => -58,
    13322 => -58,
    13323 => -58,
    13324 => -58,
    13325 => -58,
    13326 => -58,
    13327 => -58,
    13328 => -58,
    13329 => -58,
    13330 => -58,
    13331 => -58,
    13332 => -58,
    13333 => -58,
    13334 => -58,
    13335 => -58,
    13336 => -58,
    13337 => -58,
    13338 => -58,
    13339 => -58,
    13340 => -58,
    13341 => -58,
    13342 => -58,
    13343 => -58,
    13344 => -58,
    13345 => -58,
    13346 => -58,
    13347 => -58,
    13348 => -58,
    13349 => -58,
    13350 => -58,
    13351 => -58,
    13352 => -58,
    13353 => -58,
    13354 => -58,
    13355 => -58,
    13356 => -58,
    13357 => -58,
    13358 => -58,
    13359 => -58,
    13360 => -58,
    13361 => -58,
    13362 => -58,
    13363 => -58,
    13364 => -58,
    13365 => -58,
    13366 => -58,
    13367 => -58,
    13368 => -58,
    13369 => -58,
    13370 => -58,
    13371 => -58,
    13372 => -58,
    13373 => -58,
    13374 => -58,
    13375 => -58,
    13376 => -58,
    13377 => -58,
    13378 => -58,
    13379 => -58,
    13380 => -58,
    13381 => -58,
    13382 => -58,
    13383 => -58,
    13384 => -58,
    13385 => -58,
    13386 => -57,
    13387 => -57,
    13388 => -57,
    13389 => -57,
    13390 => -57,
    13391 => -57,
    13392 => -57,
    13393 => -57,
    13394 => -57,
    13395 => -57,
    13396 => -57,
    13397 => -57,
    13398 => -57,
    13399 => -57,
    13400 => -57,
    13401 => -57,
    13402 => -57,
    13403 => -57,
    13404 => -57,
    13405 => -57,
    13406 => -57,
    13407 => -57,
    13408 => -57,
    13409 => -57,
    13410 => -57,
    13411 => -57,
    13412 => -57,
    13413 => -57,
    13414 => -57,
    13415 => -57,
    13416 => -57,
    13417 => -57,
    13418 => -57,
    13419 => -57,
    13420 => -57,
    13421 => -57,
    13422 => -57,
    13423 => -57,
    13424 => -57,
    13425 => -57,
    13426 => -57,
    13427 => -57,
    13428 => -57,
    13429 => -57,
    13430 => -57,
    13431 => -57,
    13432 => -57,
    13433 => -57,
    13434 => -57,
    13435 => -57,
    13436 => -57,
    13437 => -57,
    13438 => -57,
    13439 => -57,
    13440 => -57,
    13441 => -57,
    13442 => -57,
    13443 => -57,
    13444 => -57,
    13445 => -57,
    13446 => -57,
    13447 => -57,
    13448 => -57,
    13449 => -57,
    13450 => -57,
    13451 => -57,
    13452 => -57,
    13453 => -57,
    13454 => -57,
    13455 => -57,
    13456 => -57,
    13457 => -57,
    13458 => -57,
    13459 => -57,
    13460 => -57,
    13461 => -57,
    13462 => -57,
    13463 => -57,
    13464 => -57,
    13465 => -57,
    13466 => -57,
    13467 => -57,
    13468 => -57,
    13469 => -57,
    13470 => -57,
    13471 => -57,
    13472 => -57,
    13473 => -57,
    13474 => -57,
    13475 => -57,
    13476 => -57,
    13477 => -57,
    13478 => -57,
    13479 => -57,
    13480 => -57,
    13481 => -57,
    13482 => -57,
    13483 => -56,
    13484 => -56,
    13485 => -56,
    13486 => -56,
    13487 => -56,
    13488 => -56,
    13489 => -56,
    13490 => -56,
    13491 => -56,
    13492 => -56,
    13493 => -56,
    13494 => -56,
    13495 => -56,
    13496 => -56,
    13497 => -56,
    13498 => -56,
    13499 => -56,
    13500 => -56,
    13501 => -56,
    13502 => -56,
    13503 => -56,
    13504 => -56,
    13505 => -56,
    13506 => -56,
    13507 => -56,
    13508 => -56,
    13509 => -56,
    13510 => -56,
    13511 => -56,
    13512 => -56,
    13513 => -56,
    13514 => -56,
    13515 => -56,
    13516 => -56,
    13517 => -56,
    13518 => -56,
    13519 => -56,
    13520 => -56,
    13521 => -56,
    13522 => -56,
    13523 => -56,
    13524 => -56,
    13525 => -56,
    13526 => -56,
    13527 => -56,
    13528 => -56,
    13529 => -56,
    13530 => -56,
    13531 => -56,
    13532 => -56,
    13533 => -56,
    13534 => -56,
    13535 => -56,
    13536 => -56,
    13537 => -56,
    13538 => -56,
    13539 => -56,
    13540 => -56,
    13541 => -56,
    13542 => -56,
    13543 => -56,
    13544 => -56,
    13545 => -56,
    13546 => -56,
    13547 => -56,
    13548 => -56,
    13549 => -56,
    13550 => -56,
    13551 => -56,
    13552 => -56,
    13553 => -56,
    13554 => -56,
    13555 => -56,
    13556 => -56,
    13557 => -56,
    13558 => -56,
    13559 => -56,
    13560 => -56,
    13561 => -56,
    13562 => -56,
    13563 => -56,
    13564 => -56,
    13565 => -56,
    13566 => -56,
    13567 => -56,
    13568 => -56,
    13569 => -56,
    13570 => -56,
    13571 => -56,
    13572 => -56,
    13573 => -56,
    13574 => -55,
    13575 => -55,
    13576 => -55,
    13577 => -55,
    13578 => -55,
    13579 => -55,
    13580 => -55,
    13581 => -55,
    13582 => -55,
    13583 => -55,
    13584 => -55,
    13585 => -55,
    13586 => -55,
    13587 => -55,
    13588 => -55,
    13589 => -55,
    13590 => -55,
    13591 => -55,
    13592 => -55,
    13593 => -55,
    13594 => -55,
    13595 => -55,
    13596 => -55,
    13597 => -55,
    13598 => -55,
    13599 => -55,
    13600 => -55,
    13601 => -55,
    13602 => -55,
    13603 => -55,
    13604 => -55,
    13605 => -55,
    13606 => -55,
    13607 => -55,
    13608 => -55,
    13609 => -55,
    13610 => -55,
    13611 => -55,
    13612 => -55,
    13613 => -55,
    13614 => -55,
    13615 => -55,
    13616 => -55,
    13617 => -55,
    13618 => -55,
    13619 => -55,
    13620 => -55,
    13621 => -55,
    13622 => -55,
    13623 => -55,
    13624 => -55,
    13625 => -55,
    13626 => -55,
    13627 => -55,
    13628 => -55,
    13629 => -55,
    13630 => -55,
    13631 => -55,
    13632 => -55,
    13633 => -55,
    13634 => -55,
    13635 => -55,
    13636 => -55,
    13637 => -55,
    13638 => -55,
    13639 => -55,
    13640 => -55,
    13641 => -55,
    13642 => -55,
    13643 => -55,
    13644 => -55,
    13645 => -55,
    13646 => -55,
    13647 => -55,
    13648 => -55,
    13649 => -55,
    13650 => -55,
    13651 => -55,
    13652 => -55,
    13653 => -55,
    13654 => -55,
    13655 => -55,
    13656 => -55,
    13657 => -55,
    13658 => -55,
    13659 => -54,
    13660 => -54,
    13661 => -54,
    13662 => -54,
    13663 => -54,
    13664 => -54,
    13665 => -54,
    13666 => -54,
    13667 => -54,
    13668 => -54,
    13669 => -54,
    13670 => -54,
    13671 => -54,
    13672 => -54,
    13673 => -54,
    13674 => -54,
    13675 => -54,
    13676 => -54,
    13677 => -54,
    13678 => -54,
    13679 => -54,
    13680 => -54,
    13681 => -54,
    13682 => -54,
    13683 => -54,
    13684 => -54,
    13685 => -54,
    13686 => -54,
    13687 => -54,
    13688 => -54,
    13689 => -54,
    13690 => -54,
    13691 => -54,
    13692 => -54,
    13693 => -54,
    13694 => -54,
    13695 => -54,
    13696 => -54,
    13697 => -54,
    13698 => -54,
    13699 => -54,
    13700 => -54,
    13701 => -54,
    13702 => -54,
    13703 => -54,
    13704 => -54,
    13705 => -54,
    13706 => -54,
    13707 => -54,
    13708 => -54,
    13709 => -54,
    13710 => -54,
    13711 => -54,
    13712 => -54,
    13713 => -54,
    13714 => -54,
    13715 => -54,
    13716 => -54,
    13717 => -54,
    13718 => -54,
    13719 => -54,
    13720 => -54,
    13721 => -54,
    13722 => -54,
    13723 => -54,
    13724 => -54,
    13725 => -54,
    13726 => -54,
    13727 => -54,
    13728 => -54,
    13729 => -54,
    13730 => -54,
    13731 => -54,
    13732 => -54,
    13733 => -54,
    13734 => -54,
    13735 => -54,
    13736 => -54,
    13737 => -54,
    13738 => -54,
    13739 => -53,
    13740 => -53,
    13741 => -53,
    13742 => -53,
    13743 => -53,
    13744 => -53,
    13745 => -53,
    13746 => -53,
    13747 => -53,
    13748 => -53,
    13749 => -53,
    13750 => -53,
    13751 => -53,
    13752 => -53,
    13753 => -53,
    13754 => -53,
    13755 => -53,
    13756 => -53,
    13757 => -53,
    13758 => -53,
    13759 => -53,
    13760 => -53,
    13761 => -53,
    13762 => -53,
    13763 => -53,
    13764 => -53,
    13765 => -53,
    13766 => -53,
    13767 => -53,
    13768 => -53,
    13769 => -53,
    13770 => -53,
    13771 => -53,
    13772 => -53,
    13773 => -53,
    13774 => -53,
    13775 => -53,
    13776 => -53,
    13777 => -53,
    13778 => -53,
    13779 => -53,
    13780 => -53,
    13781 => -53,
    13782 => -53,
    13783 => -53,
    13784 => -53,
    13785 => -53,
    13786 => -53,
    13787 => -53,
    13788 => -53,
    13789 => -53,
    13790 => -53,
    13791 => -53,
    13792 => -53,
    13793 => -53,
    13794 => -53,
    13795 => -53,
    13796 => -53,
    13797 => -53,
    13798 => -53,
    13799 => -53,
    13800 => -53,
    13801 => -53,
    13802 => -53,
    13803 => -53,
    13804 => -53,
    13805 => -53,
    13806 => -53,
    13807 => -53,
    13808 => -53,
    13809 => -53,
    13810 => -53,
    13811 => -53,
    13812 => -53,
    13813 => -53,
    13814 => -53,
    13815 => -53,
    13816 => -52,
    13817 => -52,
    13818 => -52,
    13819 => -52,
    13820 => -52,
    13821 => -52,
    13822 => -52,
    13823 => -52,
    13824 => -52,
    13825 => -52,
    13826 => -52,
    13827 => -52,
    13828 => -52,
    13829 => -52,
    13830 => -52,
    13831 => -52,
    13832 => -52,
    13833 => -52,
    13834 => -52,
    13835 => -52,
    13836 => -52,
    13837 => -52,
    13838 => -52,
    13839 => -52,
    13840 => -52,
    13841 => -52,
    13842 => -52,
    13843 => -52,
    13844 => -52,
    13845 => -52,
    13846 => -52,
    13847 => -52,
    13848 => -52,
    13849 => -52,
    13850 => -52,
    13851 => -52,
    13852 => -52,
    13853 => -52,
    13854 => -52,
    13855 => -52,
    13856 => -52,
    13857 => -52,
    13858 => -52,
    13859 => -52,
    13860 => -52,
    13861 => -52,
    13862 => -52,
    13863 => -52,
    13864 => -52,
    13865 => -52,
    13866 => -52,
    13867 => -52,
    13868 => -52,
    13869 => -52,
    13870 => -52,
    13871 => -52,
    13872 => -52,
    13873 => -52,
    13874 => -52,
    13875 => -52,
    13876 => -52,
    13877 => -52,
    13878 => -52,
    13879 => -52,
    13880 => -52,
    13881 => -52,
    13882 => -52,
    13883 => -52,
    13884 => -52,
    13885 => -52,
    13886 => -52,
    13887 => -52,
    13888 => -52,
    13889 => -51,
    13890 => -51,
    13891 => -51,
    13892 => -51,
    13893 => -51,
    13894 => -51,
    13895 => -51,
    13896 => -51,
    13897 => -51,
    13898 => -51,
    13899 => -51,
    13900 => -51,
    13901 => -51,
    13902 => -51,
    13903 => -51,
    13904 => -51,
    13905 => -51,
    13906 => -51,
    13907 => -51,
    13908 => -51,
    13909 => -51,
    13910 => -51,
    13911 => -51,
    13912 => -51,
    13913 => -51,
    13914 => -51,
    13915 => -51,
    13916 => -51,
    13917 => -51,
    13918 => -51,
    13919 => -51,
    13920 => -51,
    13921 => -51,
    13922 => -51,
    13923 => -51,
    13924 => -51,
    13925 => -51,
    13926 => -51,
    13927 => -51,
    13928 => -51,
    13929 => -51,
    13930 => -51,
    13931 => -51,
    13932 => -51,
    13933 => -51,
    13934 => -51,
    13935 => -51,
    13936 => -51,
    13937 => -51,
    13938 => -51,
    13939 => -51,
    13940 => -51,
    13941 => -51,
    13942 => -51,
    13943 => -51,
    13944 => -51,
    13945 => -51,
    13946 => -51,
    13947 => -51,
    13948 => -51,
    13949 => -51,
    13950 => -51,
    13951 => -51,
    13952 => -51,
    13953 => -51,
    13954 => -51,
    13955 => -51,
    13956 => -51,
    13957 => -51,
    13958 => -51,
    13959 => -51,
    13960 => -50,
    13961 => -50,
    13962 => -50,
    13963 => -50,
    13964 => -50,
    13965 => -50,
    13966 => -50,
    13967 => -50,
    13968 => -50,
    13969 => -50,
    13970 => -50,
    13971 => -50,
    13972 => -50,
    13973 => -50,
    13974 => -50,
    13975 => -50,
    13976 => -50,
    13977 => -50,
    13978 => -50,
    13979 => -50,
    13980 => -50,
    13981 => -50,
    13982 => -50,
    13983 => -50,
    13984 => -50,
    13985 => -50,
    13986 => -50,
    13987 => -50,
    13988 => -50,
    13989 => -50,
    13990 => -50,
    13991 => -50,
    13992 => -50,
    13993 => -50,
    13994 => -50,
    13995 => -50,
    13996 => -50,
    13997 => -50,
    13998 => -50,
    13999 => -50,
    14000 => -50,
    14001 => -50,
    14002 => -50,
    14003 => -50,
    14004 => -50,
    14005 => -50,
    14006 => -50,
    14007 => -50,
    14008 => -50,
    14009 => -50,
    14010 => -50,
    14011 => -50,
    14012 => -50,
    14013 => -50,
    14014 => -50,
    14015 => -50,
    14016 => -50,
    14017 => -50,
    14018 => -50,
    14019 => -50,
    14020 => -50,
    14021 => -50,
    14022 => -50,
    14023 => -50,
    14024 => -50,
    14025 => -50,
    14026 => -50,
    14027 => -50,
    14028 => -49,
    14029 => -49,
    14030 => -49,
    14031 => -49,
    14032 => -49,
    14033 => -49,
    14034 => -49,
    14035 => -49,
    14036 => -49,
    14037 => -49,
    14038 => -49,
    14039 => -49,
    14040 => -49,
    14041 => -49,
    14042 => -49,
    14043 => -49,
    14044 => -49,
    14045 => -49,
    14046 => -49,
    14047 => -49,
    14048 => -49,
    14049 => -49,
    14050 => -49,
    14051 => -49,
    14052 => -49,
    14053 => -49,
    14054 => -49,
    14055 => -49,
    14056 => -49,
    14057 => -49,
    14058 => -49,
    14059 => -49,
    14060 => -49,
    14061 => -49,
    14062 => -49,
    14063 => -49,
    14064 => -49,
    14065 => -49,
    14066 => -49,
    14067 => -49,
    14068 => -49,
    14069 => -49,
    14070 => -49,
    14071 => -49,
    14072 => -49,
    14073 => -49,
    14074 => -49,
    14075 => -49,
    14076 => -49,
    14077 => -49,
    14078 => -49,
    14079 => -49,
    14080 => -49,
    14081 => -49,
    14082 => -49,
    14083 => -49,
    14084 => -49,
    14085 => -49,
    14086 => -49,
    14087 => -49,
    14088 => -49,
    14089 => -49,
    14090 => -49,
    14091 => -49,
    14092 => -49,
    14093 => -48,
    14094 => -48,
    14095 => -48,
    14096 => -48,
    14097 => -48,
    14098 => -48,
    14099 => -48,
    14100 => -48,
    14101 => -48,
    14102 => -48,
    14103 => -48,
    14104 => -48,
    14105 => -48,
    14106 => -48,
    14107 => -48,
    14108 => -48,
    14109 => -48,
    14110 => -48,
    14111 => -48,
    14112 => -48,
    14113 => -48,
    14114 => -48,
    14115 => -48,
    14116 => -48,
    14117 => -48,
    14118 => -48,
    14119 => -48,
    14120 => -48,
    14121 => -48,
    14122 => -48,
    14123 => -48,
    14124 => -48,
    14125 => -48,
    14126 => -48,
    14127 => -48,
    14128 => -48,
    14129 => -48,
    14130 => -48,
    14131 => -48,
    14132 => -48,
    14133 => -48,
    14134 => -48,
    14135 => -48,
    14136 => -48,
    14137 => -48,
    14138 => -48,
    14139 => -48,
    14140 => -48,
    14141 => -48,
    14142 => -48,
    14143 => -48,
    14144 => -48,
    14145 => -48,
    14146 => -48,
    14147 => -48,
    14148 => -48,
    14149 => -48,
    14150 => -48,
    14151 => -48,
    14152 => -48,
    14153 => -48,
    14154 => -48,
    14155 => -48,
    14156 => -48,
    14157 => -47,
    14158 => -47,
    14159 => -47,
    14160 => -47,
    14161 => -47,
    14162 => -47,
    14163 => -47,
    14164 => -47,
    14165 => -47,
    14166 => -47,
    14167 => -47,
    14168 => -47,
    14169 => -47,
    14170 => -47,
    14171 => -47,
    14172 => -47,
    14173 => -47,
    14174 => -47,
    14175 => -47,
    14176 => -47,
    14177 => -47,
    14178 => -47,
    14179 => -47,
    14180 => -47,
    14181 => -47,
    14182 => -47,
    14183 => -47,
    14184 => -47,
    14185 => -47,
    14186 => -47,
    14187 => -47,
    14188 => -47,
    14189 => -47,
    14190 => -47,
    14191 => -47,
    14192 => -47,
    14193 => -47,
    14194 => -47,
    14195 => -47,
    14196 => -47,
    14197 => -47,
    14198 => -47,
    14199 => -47,
    14200 => -47,
    14201 => -47,
    14202 => -47,
    14203 => -47,
    14204 => -47,
    14205 => -47,
    14206 => -47,
    14207 => -47,
    14208 => -47,
    14209 => -47,
    14210 => -47,
    14211 => -47,
    14212 => -47,
    14213 => -47,
    14214 => -47,
    14215 => -47,
    14216 => -47,
    14217 => -47,
    14218 => -47,
    14219 => -47,
    14220 => -46,
    14221 => -46,
    14222 => -46,
    14223 => -46,
    14224 => -46,
    14225 => -46,
    14226 => -46,
    14227 => -46,
    14228 => -46,
    14229 => -46,
    14230 => -46,
    14231 => -46,
    14232 => -46,
    14233 => -46,
    14234 => -46,
    14235 => -46,
    14236 => -46,
    14237 => -46,
    14238 => -46,
    14239 => -46,
    14240 => -46,
    14241 => -46,
    14242 => -46,
    14243 => -46,
    14244 => -46,
    14245 => -46,
    14246 => -46,
    14247 => -46,
    14248 => -46,
    14249 => -46,
    14250 => -46,
    14251 => -46,
    14252 => -46,
    14253 => -46,
    14254 => -46,
    14255 => -46,
    14256 => -46,
    14257 => -46,
    14258 => -46,
    14259 => -46,
    14260 => -46,
    14261 => -46,
    14262 => -46,
    14263 => -46,
    14264 => -46,
    14265 => -46,
    14266 => -46,
    14267 => -46,
    14268 => -46,
    14269 => -46,
    14270 => -46,
    14271 => -46,
    14272 => -46,
    14273 => -46,
    14274 => -46,
    14275 => -46,
    14276 => -46,
    14277 => -46,
    14278 => -46,
    14279 => -46,
    14280 => -45,
    14281 => -45,
    14282 => -45,
    14283 => -45,
    14284 => -45,
    14285 => -45,
    14286 => -45,
    14287 => -45,
    14288 => -45,
    14289 => -45,
    14290 => -45,
    14291 => -45,
    14292 => -45,
    14293 => -45,
    14294 => -45,
    14295 => -45,
    14296 => -45,
    14297 => -45,
    14298 => -45,
    14299 => -45,
    14300 => -45,
    14301 => -45,
    14302 => -45,
    14303 => -45,
    14304 => -45,
    14305 => -45,
    14306 => -45,
    14307 => -45,
    14308 => -45,
    14309 => -45,
    14310 => -45,
    14311 => -45,
    14312 => -45,
    14313 => -45,
    14314 => -45,
    14315 => -45,
    14316 => -45,
    14317 => -45,
    14318 => -45,
    14319 => -45,
    14320 => -45,
    14321 => -45,
    14322 => -45,
    14323 => -45,
    14324 => -45,
    14325 => -45,
    14326 => -45,
    14327 => -45,
    14328 => -45,
    14329 => -45,
    14330 => -45,
    14331 => -45,
    14332 => -45,
    14333 => -45,
    14334 => -45,
    14335 => -45,
    14336 => -45,
    14337 => -45,
    14338 => -45,
    14339 => -44,
    14340 => -44,
    14341 => -44,
    14342 => -44,
    14343 => -44,
    14344 => -44,
    14345 => -44,
    14346 => -44,
    14347 => -44,
    14348 => -44,
    14349 => -44,
    14350 => -44,
    14351 => -44,
    14352 => -44,
    14353 => -44,
    14354 => -44,
    14355 => -44,
    14356 => -44,
    14357 => -44,
    14358 => -44,
    14359 => -44,
    14360 => -44,
    14361 => -44,
    14362 => -44,
    14363 => -44,
    14364 => -44,
    14365 => -44,
    14366 => -44,
    14367 => -44,
    14368 => -44,
    14369 => -44,
    14370 => -44,
    14371 => -44,
    14372 => -44,
    14373 => -44,
    14374 => -44,
    14375 => -44,
    14376 => -44,
    14377 => -44,
    14378 => -44,
    14379 => -44,
    14380 => -44,
    14381 => -44,
    14382 => -44,
    14383 => -44,
    14384 => -44,
    14385 => -44,
    14386 => -44,
    14387 => -44,
    14388 => -44,
    14389 => -44,
    14390 => -44,
    14391 => -44,
    14392 => -44,
    14393 => -44,
    14394 => -44,
    14395 => -44,
    14396 => -44,
    14397 => -43,
    14398 => -43,
    14399 => -43,
    14400 => -43,
    14401 => -43,
    14402 => -43,
    14403 => -43,
    14404 => -43,
    14405 => -43,
    14406 => -43,
    14407 => -43,
    14408 => -43,
    14409 => -43,
    14410 => -43,
    14411 => -43,
    14412 => -43,
    14413 => -43,
    14414 => -43,
    14415 => -43,
    14416 => -43,
    14417 => -43,
    14418 => -43,
    14419 => -43,
    14420 => -43,
    14421 => -43,
    14422 => -43,
    14423 => -43,
    14424 => -43,
    14425 => -43,
    14426 => -43,
    14427 => -43,
    14428 => -43,
    14429 => -43,
    14430 => -43,
    14431 => -43,
    14432 => -43,
    14433 => -43,
    14434 => -43,
    14435 => -43,
    14436 => -43,
    14437 => -43,
    14438 => -43,
    14439 => -43,
    14440 => -43,
    14441 => -43,
    14442 => -43,
    14443 => -43,
    14444 => -43,
    14445 => -43,
    14446 => -43,
    14447 => -43,
    14448 => -43,
    14449 => -43,
    14450 => -43,
    14451 => -43,
    14452 => -43,
    14453 => -43,
    14454 => -42,
    14455 => -42,
    14456 => -42,
    14457 => -42,
    14458 => -42,
    14459 => -42,
    14460 => -42,
    14461 => -42,
    14462 => -42,
    14463 => -42,
    14464 => -42,
    14465 => -42,
    14466 => -42,
    14467 => -42,
    14468 => -42,
    14469 => -42,
    14470 => -42,
    14471 => -42,
    14472 => -42,
    14473 => -42,
    14474 => -42,
    14475 => -42,
    14476 => -42,
    14477 => -42,
    14478 => -42,
    14479 => -42,
    14480 => -42,
    14481 => -42,
    14482 => -42,
    14483 => -42,
    14484 => -42,
    14485 => -42,
    14486 => -42,
    14487 => -42,
    14488 => -42,
    14489 => -42,
    14490 => -42,
    14491 => -42,
    14492 => -42,
    14493 => -42,
    14494 => -42,
    14495 => -42,
    14496 => -42,
    14497 => -42,
    14498 => -42,
    14499 => -42,
    14500 => -42,
    14501 => -42,
    14502 => -42,
    14503 => -42,
    14504 => -42,
    14505 => -42,
    14506 => -42,
    14507 => -42,
    14508 => -42,
    14509 => -41,
    14510 => -41,
    14511 => -41,
    14512 => -41,
    14513 => -41,
    14514 => -41,
    14515 => -41,
    14516 => -41,
    14517 => -41,
    14518 => -41,
    14519 => -41,
    14520 => -41,
    14521 => -41,
    14522 => -41,
    14523 => -41,
    14524 => -41,
    14525 => -41,
    14526 => -41,
    14527 => -41,
    14528 => -41,
    14529 => -41,
    14530 => -41,
    14531 => -41,
    14532 => -41,
    14533 => -41,
    14534 => -41,
    14535 => -41,
    14536 => -41,
    14537 => -41,
    14538 => -41,
    14539 => -41,
    14540 => -41,
    14541 => -41,
    14542 => -41,
    14543 => -41,
    14544 => -41,
    14545 => -41,
    14546 => -41,
    14547 => -41,
    14548 => -41,
    14549 => -41,
    14550 => -41,
    14551 => -41,
    14552 => -41,
    14553 => -41,
    14554 => -41,
    14555 => -41,
    14556 => -41,
    14557 => -41,
    14558 => -41,
    14559 => -41,
    14560 => -41,
    14561 => -41,
    14562 => -41,
    14563 => -41,
    14564 => -40,
    14565 => -40,
    14566 => -40,
    14567 => -40,
    14568 => -40,
    14569 => -40,
    14570 => -40,
    14571 => -40,
    14572 => -40,
    14573 => -40,
    14574 => -40,
    14575 => -40,
    14576 => -40,
    14577 => -40,
    14578 => -40,
    14579 => -40,
    14580 => -40,
    14581 => -40,
    14582 => -40,
    14583 => -40,
    14584 => -40,
    14585 => -40,
    14586 => -40,
    14587 => -40,
    14588 => -40,
    14589 => -40,
    14590 => -40,
    14591 => -40,
    14592 => -40,
    14593 => -40,
    14594 => -40,
    14595 => -40,
    14596 => -40,
    14597 => -40,
    14598 => -40,
    14599 => -40,
    14600 => -40,
    14601 => -40,
    14602 => -40,
    14603 => -40,
    14604 => -40,
    14605 => -40,
    14606 => -40,
    14607 => -40,
    14608 => -40,
    14609 => -40,
    14610 => -40,
    14611 => -40,
    14612 => -40,
    14613 => -40,
    14614 => -40,
    14615 => -40,
    14616 => -40,
    14617 => -39,
    14618 => -39,
    14619 => -39,
    14620 => -39,
    14621 => -39,
    14622 => -39,
    14623 => -39,
    14624 => -39,
    14625 => -39,
    14626 => -39,
    14627 => -39,
    14628 => -39,
    14629 => -39,
    14630 => -39,
    14631 => -39,
    14632 => -39,
    14633 => -39,
    14634 => -39,
    14635 => -39,
    14636 => -39,
    14637 => -39,
    14638 => -39,
    14639 => -39,
    14640 => -39,
    14641 => -39,
    14642 => -39,
    14643 => -39,
    14644 => -39,
    14645 => -39,
    14646 => -39,
    14647 => -39,
    14648 => -39,
    14649 => -39,
    14650 => -39,
    14651 => -39,
    14652 => -39,
    14653 => -39,
    14654 => -39,
    14655 => -39,
    14656 => -39,
    14657 => -39,
    14658 => -39,
    14659 => -39,
    14660 => -39,
    14661 => -39,
    14662 => -39,
    14663 => -39,
    14664 => -39,
    14665 => -39,
    14666 => -39,
    14667 => -39,
    14668 => -39,
    14669 => -39,
    14670 => -38,
    14671 => -38,
    14672 => -38,
    14673 => -38,
    14674 => -38,
    14675 => -38,
    14676 => -38,
    14677 => -38,
    14678 => -38,
    14679 => -38,
    14680 => -38,
    14681 => -38,
    14682 => -38,
    14683 => -38,
    14684 => -38,
    14685 => -38,
    14686 => -38,
    14687 => -38,
    14688 => -38,
    14689 => -38,
    14690 => -38,
    14691 => -38,
    14692 => -38,
    14693 => -38,
    14694 => -38,
    14695 => -38,
    14696 => -38,
    14697 => -38,
    14698 => -38,
    14699 => -38,
    14700 => -38,
    14701 => -38,
    14702 => -38,
    14703 => -38,
    14704 => -38,
    14705 => -38,
    14706 => -38,
    14707 => -38,
    14708 => -38,
    14709 => -38,
    14710 => -38,
    14711 => -38,
    14712 => -38,
    14713 => -38,
    14714 => -38,
    14715 => -38,
    14716 => -38,
    14717 => -38,
    14718 => -38,
    14719 => -38,
    14720 => -38,
    14721 => -38,
    14722 => -37,
    14723 => -37,
    14724 => -37,
    14725 => -37,
    14726 => -37,
    14727 => -37,
    14728 => -37,
    14729 => -37,
    14730 => -37,
    14731 => -37,
    14732 => -37,
    14733 => -37,
    14734 => -37,
    14735 => -37,
    14736 => -37,
    14737 => -37,
    14738 => -37,
    14739 => -37,
    14740 => -37,
    14741 => -37,
    14742 => -37,
    14743 => -37,
    14744 => -37,
    14745 => -37,
    14746 => -37,
    14747 => -37,
    14748 => -37,
    14749 => -37,
    14750 => -37,
    14751 => -37,
    14752 => -37,
    14753 => -37,
    14754 => -37,
    14755 => -37,
    14756 => -37,
    14757 => -37,
    14758 => -37,
    14759 => -37,
    14760 => -37,
    14761 => -37,
    14762 => -37,
    14763 => -37,
    14764 => -37,
    14765 => -37,
    14766 => -37,
    14767 => -37,
    14768 => -37,
    14769 => -37,
    14770 => -37,
    14771 => -37,
    14772 => -37,
    14773 => -36,
    14774 => -36,
    14775 => -36,
    14776 => -36,
    14777 => -36,
    14778 => -36,
    14779 => -36,
    14780 => -36,
    14781 => -36,
    14782 => -36,
    14783 => -36,
    14784 => -36,
    14785 => -36,
    14786 => -36,
    14787 => -36,
    14788 => -36,
    14789 => -36,
    14790 => -36,
    14791 => -36,
    14792 => -36,
    14793 => -36,
    14794 => -36,
    14795 => -36,
    14796 => -36,
    14797 => -36,
    14798 => -36,
    14799 => -36,
    14800 => -36,
    14801 => -36,
    14802 => -36,
    14803 => -36,
    14804 => -36,
    14805 => -36,
    14806 => -36,
    14807 => -36,
    14808 => -36,
    14809 => -36,
    14810 => -36,
    14811 => -36,
    14812 => -36,
    14813 => -36,
    14814 => -36,
    14815 => -36,
    14816 => -36,
    14817 => -36,
    14818 => -36,
    14819 => -36,
    14820 => -36,
    14821 => -36,
    14822 => -36,
    14823 => -36,
    14824 => -35,
    14825 => -35,
    14826 => -35,
    14827 => -35,
    14828 => -35,
    14829 => -35,
    14830 => -35,
    14831 => -35,
    14832 => -35,
    14833 => -35,
    14834 => -35,
    14835 => -35,
    14836 => -35,
    14837 => -35,
    14838 => -35,
    14839 => -35,
    14840 => -35,
    14841 => -35,
    14842 => -35,
    14843 => -35,
    14844 => -35,
    14845 => -35,
    14846 => -35,
    14847 => -35,
    14848 => -35,
    14849 => -35,
    14850 => -35,
    14851 => -35,
    14852 => -35,
    14853 => -35,
    14854 => -35,
    14855 => -35,
    14856 => -35,
    14857 => -35,
    14858 => -35,
    14859 => -35,
    14860 => -35,
    14861 => -35,
    14862 => -35,
    14863 => -35,
    14864 => -35,
    14865 => -35,
    14866 => -35,
    14867 => -35,
    14868 => -35,
    14869 => -35,
    14870 => -35,
    14871 => -35,
    14872 => -35,
    14873 => -34,
    14874 => -34,
    14875 => -34,
    14876 => -34,
    14877 => -34,
    14878 => -34,
    14879 => -34,
    14880 => -34,
    14881 => -34,
    14882 => -34,
    14883 => -34,
    14884 => -34,
    14885 => -34,
    14886 => -34,
    14887 => -34,
    14888 => -34,
    14889 => -34,
    14890 => -34,
    14891 => -34,
    14892 => -34,
    14893 => -34,
    14894 => -34,
    14895 => -34,
    14896 => -34,
    14897 => -34,
    14898 => -34,
    14899 => -34,
    14900 => -34,
    14901 => -34,
    14902 => -34,
    14903 => -34,
    14904 => -34,
    14905 => -34,
    14906 => -34,
    14907 => -34,
    14908 => -34,
    14909 => -34,
    14910 => -34,
    14911 => -34,
    14912 => -34,
    14913 => -34,
    14914 => -34,
    14915 => -34,
    14916 => -34,
    14917 => -34,
    14918 => -34,
    14919 => -34,
    14920 => -34,
    14921 => -34,
    14922 => -34,
    14923 => -33,
    14924 => -33,
    14925 => -33,
    14926 => -33,
    14927 => -33,
    14928 => -33,
    14929 => -33,
    14930 => -33,
    14931 => -33,
    14932 => -33,
    14933 => -33,
    14934 => -33,
    14935 => -33,
    14936 => -33,
    14937 => -33,
    14938 => -33,
    14939 => -33,
    14940 => -33,
    14941 => -33,
    14942 => -33,
    14943 => -33,
    14944 => -33,
    14945 => -33,
    14946 => -33,
    14947 => -33,
    14948 => -33,
    14949 => -33,
    14950 => -33,
    14951 => -33,
    14952 => -33,
    14953 => -33,
    14954 => -33,
    14955 => -33,
    14956 => -33,
    14957 => -33,
    14958 => -33,
    14959 => -33,
    14960 => -33,
    14961 => -33,
    14962 => -33,
    14963 => -33,
    14964 => -33,
    14965 => -33,
    14966 => -33,
    14967 => -33,
    14968 => -33,
    14969 => -33,
    14970 => -33,
    14971 => -32,
    14972 => -32,
    14973 => -32,
    14974 => -32,
    14975 => -32,
    14976 => -32,
    14977 => -32,
    14978 => -32,
    14979 => -32,
    14980 => -32,
    14981 => -32,
    14982 => -32,
    14983 => -32,
    14984 => -32,
    14985 => -32,
    14986 => -32,
    14987 => -32,
    14988 => -32,
    14989 => -32,
    14990 => -32,
    14991 => -32,
    14992 => -32,
    14993 => -32,
    14994 => -32,
    14995 => -32,
    14996 => -32,
    14997 => -32,
    14998 => -32,
    14999 => -32,
    15000 => -32,
    15001 => -32,
    15002 => -32,
    15003 => -32,
    15004 => -32,
    15005 => -32,
    15006 => -32,
    15007 => -32,
    15008 => -32,
    15009 => -32,
    15010 => -32,
    15011 => -32,
    15012 => -32,
    15013 => -32,
    15014 => -32,
    15015 => -32,
    15016 => -32,
    15017 => -32,
    15018 => -32,
    15019 => -31,
    15020 => -31,
    15021 => -31,
    15022 => -31,
    15023 => -31,
    15024 => -31,
    15025 => -31,
    15026 => -31,
    15027 => -31,
    15028 => -31,
    15029 => -31,
    15030 => -31,
    15031 => -31,
    15032 => -31,
    15033 => -31,
    15034 => -31,
    15035 => -31,
    15036 => -31,
    15037 => -31,
    15038 => -31,
    15039 => -31,
    15040 => -31,
    15041 => -31,
    15042 => -31,
    15043 => -31,
    15044 => -31,
    15045 => -31,
    15046 => -31,
    15047 => -31,
    15048 => -31,
    15049 => -31,
    15050 => -31,
    15051 => -31,
    15052 => -31,
    15053 => -31,
    15054 => -31,
    15055 => -31,
    15056 => -31,
    15057 => -31,
    15058 => -31,
    15059 => -31,
    15060 => -31,
    15061 => -31,
    15062 => -31,
    15063 => -31,
    15064 => -31,
    15065 => -31,
    15066 => -31,
    15067 => -30,
    15068 => -30,
    15069 => -30,
    15070 => -30,
    15071 => -30,
    15072 => -30,
    15073 => -30,
    15074 => -30,
    15075 => -30,
    15076 => -30,
    15077 => -30,
    15078 => -30,
    15079 => -30,
    15080 => -30,
    15081 => -30,
    15082 => -30,
    15083 => -30,
    15084 => -30,
    15085 => -30,
    15086 => -30,
    15087 => -30,
    15088 => -30,
    15089 => -30,
    15090 => -30,
    15091 => -30,
    15092 => -30,
    15093 => -30,
    15094 => -30,
    15095 => -30,
    15096 => -30,
    15097 => -30,
    15098 => -30,
    15099 => -30,
    15100 => -30,
    15101 => -30,
    15102 => -30,
    15103 => -30,
    15104 => -30,
    15105 => -30,
    15106 => -30,
    15107 => -30,
    15108 => -30,
    15109 => -30,
    15110 => -30,
    15111 => -30,
    15112 => -30,
    15113 => -30,
    15114 => -29,
    15115 => -29,
    15116 => -29,
    15117 => -29,
    15118 => -29,
    15119 => -29,
    15120 => -29,
    15121 => -29,
    15122 => -29,
    15123 => -29,
    15124 => -29,
    15125 => -29,
    15126 => -29,
    15127 => -29,
    15128 => -29,
    15129 => -29,
    15130 => -29,
    15131 => -29,
    15132 => -29,
    15133 => -29,
    15134 => -29,
    15135 => -29,
    15136 => -29,
    15137 => -29,
    15138 => -29,
    15139 => -29,
    15140 => -29,
    15141 => -29,
    15142 => -29,
    15143 => -29,
    15144 => -29,
    15145 => -29,
    15146 => -29,
    15147 => -29,
    15148 => -29,
    15149 => -29,
    15150 => -29,
    15151 => -29,
    15152 => -29,
    15153 => -29,
    15154 => -29,
    15155 => -29,
    15156 => -29,
    15157 => -29,
    15158 => -29,
    15159 => -29,
    15160 => -28,
    15161 => -28,
    15162 => -28,
    15163 => -28,
    15164 => -28,
    15165 => -28,
    15166 => -28,
    15167 => -28,
    15168 => -28,
    15169 => -28,
    15170 => -28,
    15171 => -28,
    15172 => -28,
    15173 => -28,
    15174 => -28,
    15175 => -28,
    15176 => -28,
    15177 => -28,
    15178 => -28,
    15179 => -28,
    15180 => -28,
    15181 => -28,
    15182 => -28,
    15183 => -28,
    15184 => -28,
    15185 => -28,
    15186 => -28,
    15187 => -28,
    15188 => -28,
    15189 => -28,
    15190 => -28,
    15191 => -28,
    15192 => -28,
    15193 => -28,
    15194 => -28,
    15195 => -28,
    15196 => -28,
    15197 => -28,
    15198 => -28,
    15199 => -28,
    15200 => -28,
    15201 => -28,
    15202 => -28,
    15203 => -28,
    15204 => -28,
    15205 => -28,
    15206 => -28,
    15207 => -27,
    15208 => -27,
    15209 => -27,
    15210 => -27,
    15211 => -27,
    15212 => -27,
    15213 => -27,
    15214 => -27,
    15215 => -27,
    15216 => -27,
    15217 => -27,
    15218 => -27,
    15219 => -27,
    15220 => -27,
    15221 => -27,
    15222 => -27,
    15223 => -27,
    15224 => -27,
    15225 => -27,
    15226 => -27,
    15227 => -27,
    15228 => -27,
    15229 => -27,
    15230 => -27,
    15231 => -27,
    15232 => -27,
    15233 => -27,
    15234 => -27,
    15235 => -27,
    15236 => -27,
    15237 => -27,
    15238 => -27,
    15239 => -27,
    15240 => -27,
    15241 => -27,
    15242 => -27,
    15243 => -27,
    15244 => -27,
    15245 => -27,
    15246 => -27,
    15247 => -27,
    15248 => -27,
    15249 => -27,
    15250 => -27,
    15251 => -27,
    15252 => -26,
    15253 => -26,
    15254 => -26,
    15255 => -26,
    15256 => -26,
    15257 => -26,
    15258 => -26,
    15259 => -26,
    15260 => -26,
    15261 => -26,
    15262 => -26,
    15263 => -26,
    15264 => -26,
    15265 => -26,
    15266 => -26,
    15267 => -26,
    15268 => -26,
    15269 => -26,
    15270 => -26,
    15271 => -26,
    15272 => -26,
    15273 => -26,
    15274 => -26,
    15275 => -26,
    15276 => -26,
    15277 => -26,
    15278 => -26,
    15279 => -26,
    15280 => -26,
    15281 => -26,
    15282 => -26,
    15283 => -26,
    15284 => -26,
    15285 => -26,
    15286 => -26,
    15287 => -26,
    15288 => -26,
    15289 => -26,
    15290 => -26,
    15291 => -26,
    15292 => -26,
    15293 => -26,
    15294 => -26,
    15295 => -26,
    15296 => -26,
    15297 => -26,
    15298 => -25,
    15299 => -25,
    15300 => -25,
    15301 => -25,
    15302 => -25,
    15303 => -25,
    15304 => -25,
    15305 => -25,
    15306 => -25,
    15307 => -25,
    15308 => -25,
    15309 => -25,
    15310 => -25,
    15311 => -25,
    15312 => -25,
    15313 => -25,
    15314 => -25,
    15315 => -25,
    15316 => -25,
    15317 => -25,
    15318 => -25,
    15319 => -25,
    15320 => -25,
    15321 => -25,
    15322 => -25,
    15323 => -25,
    15324 => -25,
    15325 => -25,
    15326 => -25,
    15327 => -25,
    15328 => -25,
    15329 => -25,
    15330 => -25,
    15331 => -25,
    15332 => -25,
    15333 => -25,
    15334 => -25,
    15335 => -25,
    15336 => -25,
    15337 => -25,
    15338 => -25,
    15339 => -25,
    15340 => -25,
    15341 => -25,
    15342 => -25,
    15343 => -24,
    15344 => -24,
    15345 => -24,
    15346 => -24,
    15347 => -24,
    15348 => -24,
    15349 => -24,
    15350 => -24,
    15351 => -24,
    15352 => -24,
    15353 => -24,
    15354 => -24,
    15355 => -24,
    15356 => -24,
    15357 => -24,
    15358 => -24,
    15359 => -24,
    15360 => -24,
    15361 => -24,
    15362 => -24,
    15363 => -24,
    15364 => -24,
    15365 => -24,
    15366 => -24,
    15367 => -24,
    15368 => -24,
    15369 => -24,
    15370 => -24,
    15371 => -24,
    15372 => -24,
    15373 => -24,
    15374 => -24,
    15375 => -24,
    15376 => -24,
    15377 => -24,
    15378 => -24,
    15379 => -24,
    15380 => -24,
    15381 => -24,
    15382 => -24,
    15383 => -24,
    15384 => -24,
    15385 => -24,
    15386 => -24,
    15387 => -24,
    15388 => -23,
    15389 => -23,
    15390 => -23,
    15391 => -23,
    15392 => -23,
    15393 => -23,
    15394 => -23,
    15395 => -23,
    15396 => -23,
    15397 => -23,
    15398 => -23,
    15399 => -23,
    15400 => -23,
    15401 => -23,
    15402 => -23,
    15403 => -23,
    15404 => -23,
    15405 => -23,
    15406 => -23,
    15407 => -23,
    15408 => -23,
    15409 => -23,
    15410 => -23,
    15411 => -23,
    15412 => -23,
    15413 => -23,
    15414 => -23,
    15415 => -23,
    15416 => -23,
    15417 => -23,
    15418 => -23,
    15419 => -23,
    15420 => -23,
    15421 => -23,
    15422 => -23,
    15423 => -23,
    15424 => -23,
    15425 => -23,
    15426 => -23,
    15427 => -23,
    15428 => -23,
    15429 => -23,
    15430 => -23,
    15431 => -23,
    15432 => -22,
    15433 => -22,
    15434 => -22,
    15435 => -22,
    15436 => -22,
    15437 => -22,
    15438 => -22,
    15439 => -22,
    15440 => -22,
    15441 => -22,
    15442 => -22,
    15443 => -22,
    15444 => -22,
    15445 => -22,
    15446 => -22,
    15447 => -22,
    15448 => -22,
    15449 => -22,
    15450 => -22,
    15451 => -22,
    15452 => -22,
    15453 => -22,
    15454 => -22,
    15455 => -22,
    15456 => -22,
    15457 => -22,
    15458 => -22,
    15459 => -22,
    15460 => -22,
    15461 => -22,
    15462 => -22,
    15463 => -22,
    15464 => -22,
    15465 => -22,
    15466 => -22,
    15467 => -22,
    15468 => -22,
    15469 => -22,
    15470 => -22,
    15471 => -22,
    15472 => -22,
    15473 => -22,
    15474 => -22,
    15475 => -22,
    15476 => -21,
    15477 => -21,
    15478 => -21,
    15479 => -21,
    15480 => -21,
    15481 => -21,
    15482 => -21,
    15483 => -21,
    15484 => -21,
    15485 => -21,
    15486 => -21,
    15487 => -21,
    15488 => -21,
    15489 => -21,
    15490 => -21,
    15491 => -21,
    15492 => -21,
    15493 => -21,
    15494 => -21,
    15495 => -21,
    15496 => -21,
    15497 => -21,
    15498 => -21,
    15499 => -21,
    15500 => -21,
    15501 => -21,
    15502 => -21,
    15503 => -21,
    15504 => -21,
    15505 => -21,
    15506 => -21,
    15507 => -21,
    15508 => -21,
    15509 => -21,
    15510 => -21,
    15511 => -21,
    15512 => -21,
    15513 => -21,
    15514 => -21,
    15515 => -21,
    15516 => -21,
    15517 => -21,
    15518 => -21,
    15519 => -21,
    15520 => -20,
    15521 => -20,
    15522 => -20,
    15523 => -20,
    15524 => -20,
    15525 => -20,
    15526 => -20,
    15527 => -20,
    15528 => -20,
    15529 => -20,
    15530 => -20,
    15531 => -20,
    15532 => -20,
    15533 => -20,
    15534 => -20,
    15535 => -20,
    15536 => -20,
    15537 => -20,
    15538 => -20,
    15539 => -20,
    15540 => -20,
    15541 => -20,
    15542 => -20,
    15543 => -20,
    15544 => -20,
    15545 => -20,
    15546 => -20,
    15547 => -20,
    15548 => -20,
    15549 => -20,
    15550 => -20,
    15551 => -20,
    15552 => -20,
    15553 => -20,
    15554 => -20,
    15555 => -20,
    15556 => -20,
    15557 => -20,
    15558 => -20,
    15559 => -20,
    15560 => -20,
    15561 => -20,
    15562 => -20,
    15563 => -20,
    15564 => -19,
    15565 => -19,
    15566 => -19,
    15567 => -19,
    15568 => -19,
    15569 => -19,
    15570 => -19,
    15571 => -19,
    15572 => -19,
    15573 => -19,
    15574 => -19,
    15575 => -19,
    15576 => -19,
    15577 => -19,
    15578 => -19,
    15579 => -19,
    15580 => -19,
    15581 => -19,
    15582 => -19,
    15583 => -19,
    15584 => -19,
    15585 => -19,
    15586 => -19,
    15587 => -19,
    15588 => -19,
    15589 => -19,
    15590 => -19,
    15591 => -19,
    15592 => -19,
    15593 => -19,
    15594 => -19,
    15595 => -19,
    15596 => -19,
    15597 => -19,
    15598 => -19,
    15599 => -19,
    15600 => -19,
    15601 => -19,
    15602 => -19,
    15603 => -19,
    15604 => -19,
    15605 => -19,
    15606 => -19,
    15607 => -18,
    15608 => -18,
    15609 => -18,
    15610 => -18,
    15611 => -18,
    15612 => -18,
    15613 => -18,
    15614 => -18,
    15615 => -18,
    15616 => -18,
    15617 => -18,
    15618 => -18,
    15619 => -18,
    15620 => -18,
    15621 => -18,
    15622 => -18,
    15623 => -18,
    15624 => -18,
    15625 => -18,
    15626 => -18,
    15627 => -18,
    15628 => -18,
    15629 => -18,
    15630 => -18,
    15631 => -18,
    15632 => -18,
    15633 => -18,
    15634 => -18,
    15635 => -18,
    15636 => -18,
    15637 => -18,
    15638 => -18,
    15639 => -18,
    15640 => -18,
    15641 => -18,
    15642 => -18,
    15643 => -18,
    15644 => -18,
    15645 => -18,
    15646 => -18,
    15647 => -18,
    15648 => -18,
    15649 => -18,
    15650 => -18,
    15651 => -17,
    15652 => -17,
    15653 => -17,
    15654 => -17,
    15655 => -17,
    15656 => -17,
    15657 => -17,
    15658 => -17,
    15659 => -17,
    15660 => -17,
    15661 => -17,
    15662 => -17,
    15663 => -17,
    15664 => -17,
    15665 => -17,
    15666 => -17,
    15667 => -17,
    15668 => -17,
    15669 => -17,
    15670 => -17,
    15671 => -17,
    15672 => -17,
    15673 => -17,
    15674 => -17,
    15675 => -17,
    15676 => -17,
    15677 => -17,
    15678 => -17,
    15679 => -17,
    15680 => -17,
    15681 => -17,
    15682 => -17,
    15683 => -17,
    15684 => -17,
    15685 => -17,
    15686 => -17,
    15687 => -17,
    15688 => -17,
    15689 => -17,
    15690 => -17,
    15691 => -17,
    15692 => -17,
    15693 => -16,
    15694 => -16,
    15695 => -16,
    15696 => -16,
    15697 => -16,
    15698 => -16,
    15699 => -16,
    15700 => -16,
    15701 => -16,
    15702 => -16,
    15703 => -16,
    15704 => -16,
    15705 => -16,
    15706 => -16,
    15707 => -16,
    15708 => -16,
    15709 => -16,
    15710 => -16,
    15711 => -16,
    15712 => -16,
    15713 => -16,
    15714 => -16,
    15715 => -16,
    15716 => -16,
    15717 => -16,
    15718 => -16,
    15719 => -16,
    15720 => -16,
    15721 => -16,
    15722 => -16,
    15723 => -16,
    15724 => -16,
    15725 => -16,
    15726 => -16,
    15727 => -16,
    15728 => -16,
    15729 => -16,
    15730 => -16,
    15731 => -16,
    15732 => -16,
    15733 => -16,
    15734 => -16,
    15735 => -16,
    15736 => -15,
    15737 => -15,
    15738 => -15,
    15739 => -15,
    15740 => -15,
    15741 => -15,
    15742 => -15,
    15743 => -15,
    15744 => -15,
    15745 => -15,
    15746 => -15,
    15747 => -15,
    15748 => -15,
    15749 => -15,
    15750 => -15,
    15751 => -15,
    15752 => -15,
    15753 => -15,
    15754 => -15,
    15755 => -15,
    15756 => -15,
    15757 => -15,
    15758 => -15,
    15759 => -15,
    15760 => -15,
    15761 => -15,
    15762 => -15,
    15763 => -15,
    15764 => -15,
    15765 => -15,
    15766 => -15,
    15767 => -15,
    15768 => -15,
    15769 => -15,
    15770 => -15,
    15771 => -15,
    15772 => -15,
    15773 => -15,
    15774 => -15,
    15775 => -15,
    15776 => -15,
    15777 => -15,
    15778 => -15,
    15779 => -14,
    15780 => -14,
    15781 => -14,
    15782 => -14,
    15783 => -14,
    15784 => -14,
    15785 => -14,
    15786 => -14,
    15787 => -14,
    15788 => -14,
    15789 => -14,
    15790 => -14,
    15791 => -14,
    15792 => -14,
    15793 => -14,
    15794 => -14,
    15795 => -14,
    15796 => -14,
    15797 => -14,
    15798 => -14,
    15799 => -14,
    15800 => -14,
    15801 => -14,
    15802 => -14,
    15803 => -14,
    15804 => -14,
    15805 => -14,
    15806 => -14,
    15807 => -14,
    15808 => -14,
    15809 => -14,
    15810 => -14,
    15811 => -14,
    15812 => -14,
    15813 => -14,
    15814 => -14,
    15815 => -14,
    15816 => -14,
    15817 => -14,
    15818 => -14,
    15819 => -14,
    15820 => -14,
    15821 => -13,
    15822 => -13,
    15823 => -13,
    15824 => -13,
    15825 => -13,
    15826 => -13,
    15827 => -13,
    15828 => -13,
    15829 => -13,
    15830 => -13,
    15831 => -13,
    15832 => -13,
    15833 => -13,
    15834 => -13,
    15835 => -13,
    15836 => -13,
    15837 => -13,
    15838 => -13,
    15839 => -13,
    15840 => -13,
    15841 => -13,
    15842 => -13,
    15843 => -13,
    15844 => -13,
    15845 => -13,
    15846 => -13,
    15847 => -13,
    15848 => -13,
    15849 => -13,
    15850 => -13,
    15851 => -13,
    15852 => -13,
    15853 => -13,
    15854 => -13,
    15855 => -13,
    15856 => -13,
    15857 => -13,
    15858 => -13,
    15859 => -13,
    15860 => -13,
    15861 => -13,
    15862 => -13,
    15863 => -13,
    15864 => -12,
    15865 => -12,
    15866 => -12,
    15867 => -12,
    15868 => -12,
    15869 => -12,
    15870 => -12,
    15871 => -12,
    15872 => -12,
    15873 => -12,
    15874 => -12,
    15875 => -12,
    15876 => -12,
    15877 => -12,
    15878 => -12,
    15879 => -12,
    15880 => -12,
    15881 => -12,
    15882 => -12,
    15883 => -12,
    15884 => -12,
    15885 => -12,
    15886 => -12,
    15887 => -12,
    15888 => -12,
    15889 => -12,
    15890 => -12,
    15891 => -12,
    15892 => -12,
    15893 => -12,
    15894 => -12,
    15895 => -12,
    15896 => -12,
    15897 => -12,
    15898 => -12,
    15899 => -12,
    15900 => -12,
    15901 => -12,
    15902 => -12,
    15903 => -12,
    15904 => -12,
    15905 => -12,
    15906 => -11,
    15907 => -11,
    15908 => -11,
    15909 => -11,
    15910 => -11,
    15911 => -11,
    15912 => -11,
    15913 => -11,
    15914 => -11,
    15915 => -11,
    15916 => -11,
    15917 => -11,
    15918 => -11,
    15919 => -11,
    15920 => -11,
    15921 => -11,
    15922 => -11,
    15923 => -11,
    15924 => -11,
    15925 => -11,
    15926 => -11,
    15927 => -11,
    15928 => -11,
    15929 => -11,
    15930 => -11,
    15931 => -11,
    15932 => -11,
    15933 => -11,
    15934 => -11,
    15935 => -11,
    15936 => -11,
    15937 => -11,
    15938 => -11,
    15939 => -11,
    15940 => -11,
    15941 => -11,
    15942 => -11,
    15943 => -11,
    15944 => -11,
    15945 => -11,
    15946 => -11,
    15947 => -11,
    15948 => -10,
    15949 => -10,
    15950 => -10,
    15951 => -10,
    15952 => -10,
    15953 => -10,
    15954 => -10,
    15955 => -10,
    15956 => -10,
    15957 => -10,
    15958 => -10,
    15959 => -10,
    15960 => -10,
    15961 => -10,
    15962 => -10,
    15963 => -10,
    15964 => -10,
    15965 => -10,
    15966 => -10,
    15967 => -10,
    15968 => -10,
    15969 => -10,
    15970 => -10,
    15971 => -10,
    15972 => -10,
    15973 => -10,
    15974 => -10,
    15975 => -10,
    15976 => -10,
    15977 => -10,
    15978 => -10,
    15979 => -10,
    15980 => -10,
    15981 => -10,
    15982 => -10,
    15983 => -10,
    15984 => -10,
    15985 => -10,
    15986 => -10,
    15987 => -10,
    15988 => -10,
    15989 => -10,
    15990 => -9,
    15991 => -9,
    15992 => -9,
    15993 => -9,
    15994 => -9,
    15995 => -9,
    15996 => -9,
    15997 => -9,
    15998 => -9,
    15999 => -9,
    16000 => -9,
    16001 => -9,
    16002 => -9,
    16003 => -9,
    16004 => -9,
    16005 => -9,
    16006 => -9,
    16007 => -9,
    16008 => -9,
    16009 => -9,
    16010 => -9,
    16011 => -9,
    16012 => -9,
    16013 => -9,
    16014 => -9,
    16015 => -9,
    16016 => -9,
    16017 => -9,
    16018 => -9,
    16019 => -9,
    16020 => -9,
    16021 => -9,
    16022 => -9,
    16023 => -9,
    16024 => -9,
    16025 => -9,
    16026 => -9,
    16027 => -9,
    16028 => -9,
    16029 => -9,
    16030 => -9,
    16031 => -9,
    16032 => -8,
    16033 => -8,
    16034 => -8,
    16035 => -8,
    16036 => -8,
    16037 => -8,
    16038 => -8,
    16039 => -8,
    16040 => -8,
    16041 => -8,
    16042 => -8,
    16043 => -8,
    16044 => -8,
    16045 => -8,
    16046 => -8,
    16047 => -8,
    16048 => -8,
    16049 => -8,
    16050 => -8,
    16051 => -8,
    16052 => -8,
    16053 => -8,
    16054 => -8,
    16055 => -8,
    16056 => -8,
    16057 => -8,
    16058 => -8,
    16059 => -8,
    16060 => -8,
    16061 => -8,
    16062 => -8,
    16063 => -8,
    16064 => -8,
    16065 => -8,
    16066 => -8,
    16067 => -8,
    16068 => -8,
    16069 => -8,
    16070 => -8,
    16071 => -8,
    16072 => -8,
    16073 => -7,
    16074 => -7,
    16075 => -7,
    16076 => -7,
    16077 => -7,
    16078 => -7,
    16079 => -7,
    16080 => -7,
    16081 => -7,
    16082 => -7,
    16083 => -7,
    16084 => -7,
    16085 => -7,
    16086 => -7,
    16087 => -7,
    16088 => -7,
    16089 => -7,
    16090 => -7,
    16091 => -7,
    16092 => -7,
    16093 => -7,
    16094 => -7,
    16095 => -7,
    16096 => -7,
    16097 => -7,
    16098 => -7,
    16099 => -7,
    16100 => -7,
    16101 => -7,
    16102 => -7,
    16103 => -7,
    16104 => -7,
    16105 => -7,
    16106 => -7,
    16107 => -7,
    16108 => -7,
    16109 => -7,
    16110 => -7,
    16111 => -7,
    16112 => -7,
    16113 => -7,
    16114 => -7,
    16115 => -6,
    16116 => -6,
    16117 => -6,
    16118 => -6,
    16119 => -6,
    16120 => -6,
    16121 => -6,
    16122 => -6,
    16123 => -6,
    16124 => -6,
    16125 => -6,
    16126 => -6,
    16127 => -6,
    16128 => -6,
    16129 => -6,
    16130 => -6,
    16131 => -6,
    16132 => -6,
    16133 => -6,
    16134 => -6,
    16135 => -6,
    16136 => -6,
    16137 => -6,
    16138 => -6,
    16139 => -6,
    16140 => -6,
    16141 => -6,
    16142 => -6,
    16143 => -6,
    16144 => -6,
    16145 => -6,
    16146 => -6,
    16147 => -6,
    16148 => -6,
    16149 => -6,
    16150 => -6,
    16151 => -6,
    16152 => -6,
    16153 => -6,
    16154 => -6,
    16155 => -6,
    16156 => -6,
    16157 => -5,
    16158 => -5,
    16159 => -5,
    16160 => -5,
    16161 => -5,
    16162 => -5,
    16163 => -5,
    16164 => -5,
    16165 => -5,
    16166 => -5,
    16167 => -5,
    16168 => -5,
    16169 => -5,
    16170 => -5,
    16171 => -5,
    16172 => -5,
    16173 => -5,
    16174 => -5,
    16175 => -5,
    16176 => -5,
    16177 => -5,
    16178 => -5,
    16179 => -5,
    16180 => -5,
    16181 => -5,
    16182 => -5,
    16183 => -5,
    16184 => -5,
    16185 => -5,
    16186 => -5,
    16187 => -5,
    16188 => -5,
    16189 => -5,
    16190 => -5,
    16191 => -5,
    16192 => -5,
    16193 => -5,
    16194 => -5,
    16195 => -5,
    16196 => -5,
    16197 => -5,
    16198 => -4,
    16199 => -4,
    16200 => -4,
    16201 => -4,
    16202 => -4,
    16203 => -4,
    16204 => -4,
    16205 => -4,
    16206 => -4,
    16207 => -4,
    16208 => -4,
    16209 => -4,
    16210 => -4,
    16211 => -4,
    16212 => -4,
    16213 => -4,
    16214 => -4,
    16215 => -4,
    16216 => -4,
    16217 => -4,
    16218 => -4,
    16219 => -4,
    16220 => -4,
    16221 => -4,
    16222 => -4,
    16223 => -4,
    16224 => -4,
    16225 => -4,
    16226 => -4,
    16227 => -4,
    16228 => -4,
    16229 => -4,
    16230 => -4,
    16231 => -4,
    16232 => -4,
    16233 => -4,
    16234 => -4,
    16235 => -4,
    16236 => -4,
    16237 => -4,
    16238 => -4,
    16239 => -4,
    16240 => -3,
    16241 => -3,
    16242 => -3,
    16243 => -3,
    16244 => -3,
    16245 => -3,
    16246 => -3,
    16247 => -3,
    16248 => -3,
    16249 => -3,
    16250 => -3,
    16251 => -3,
    16252 => -3,
    16253 => -3,
    16254 => -3,
    16255 => -3,
    16256 => -3,
    16257 => -3,
    16258 => -3,
    16259 => -3,
    16260 => -3,
    16261 => -3,
    16262 => -3,
    16263 => -3,
    16264 => -3,
    16265 => -3,
    16266 => -3,
    16267 => -3,
    16268 => -3,
    16269 => -3,
    16270 => -3,
    16271 => -3,
    16272 => -3,
    16273 => -3,
    16274 => -3,
    16275 => -3,
    16276 => -3,
    16277 => -3,
    16278 => -3,
    16279 => -3,
    16280 => -3,
    16281 => -2,
    16282 => -2,
    16283 => -2,
    16284 => -2,
    16285 => -2,
    16286 => -2,
    16287 => -2,
    16288 => -2,
    16289 => -2,
    16290 => -2,
    16291 => -2,
    16292 => -2,
    16293 => -2,
    16294 => -2,
    16295 => -2,
    16296 => -2,
    16297 => -2,
    16298 => -2,
    16299 => -2,
    16300 => -2,
    16301 => -2,
    16302 => -2,
    16303 => -2,
    16304 => -2,
    16305 => -2,
    16306 => -2,
    16307 => -2,
    16308 => -2,
    16309 => -2,
    16310 => -2,
    16311 => -2,
    16312 => -2,
    16313 => -2,
    16314 => -2,
    16315 => -2,
    16316 => -2,
    16317 => -2,
    16318 => -2,
    16319 => -2,
    16320 => -2,
    16321 => -2,
    16322 => -1,
    16323 => -1,
    16324 => -1,
    16325 => -1,
    16326 => -1,
    16327 => -1,
    16328 => -1,
    16329 => -1,
    16330 => -1,
    16331 => -1,
    16332 => -1,
    16333 => -1,
    16334 => -1,
    16335 => -1,
    16336 => -1,
    16337 => -1,
    16338 => -1,
    16339 => -1,
    16340 => -1,
    16341 => -1,
    16342 => -1,
    16343 => -1,
    16344 => -1,
    16345 => -1,
    16346 => -1,
    16347 => -1,
    16348 => -1,
    16349 => -1,
    16350 => -1,
    16351 => -1,
    16352 => -1,
    16353 => -1,
    16354 => -1,
    16355 => -1,
    16356 => -1,
    16357 => -1,
    16358 => -1,
    16359 => -1,
    16360 => -1,
    16361 => -1,
    16362 => -1,
    16363 => -1,
    16364 => 0,
    16365 => 0,
    16366 => 0,
    16367 => 0,
    16368 => 0,
    16369 => 0,
    16370 => 0,
    16371 => 0,
    16372 => 0,
    16373 => 0,
    16374 => 0,
    16375 => 0,
    16376 => 0,
    16377 => 0,
    16378 => 0,
    16379 => 0,
    16380 => 0,
    16381 => 0,
    16382 => 0,
    16383 => 0
  );

begin
  lut_out <= std_logic_vector(to_signed(LUT(to_integer(unsigned(address))),P));
end architecture;
